//Benchmark atmr_misex3_1774_0.0313

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1288_, ori_ori_n1289_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1509_, mai_mai_n1510_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1539_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  INV        o0001(.A(d), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(g), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(g), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  NO2        o0010(.A(ori_ori_n38_), .B(n), .Y(ori_ori_n39_));
  INV        o0011(.A(h), .Y(ori_ori_n40_));
  NAi21      o0012(.An(j), .B(l), .Y(ori_ori_n41_));
  NAi32      o0013(.An(n), .Bn(g), .C(m), .Y(ori_ori_n42_));
  NO3        o0014(.A(ori_ori_n42_), .B(ori_ori_n41_), .C(ori_ori_n40_), .Y(ori_ori_n43_));
  NAi31      o0015(.An(n), .B(m), .C(l), .Y(ori_ori_n44_));
  INV        o0016(.A(i), .Y(ori_ori_n45_));
  AN2        o0017(.A(h), .B(g), .Y(ori_ori_n46_));
  NA2        o0018(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o0019(.A(ori_ori_n47_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NAi21      o0020(.An(n), .B(m), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(l), .Y(ori_ori_n50_));
  NOi32      o0022(.An(k), .Bn(h), .C(g), .Y(ori_ori_n51_));
  INV        o0023(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NO2        o0024(.A(ori_ori_n52_), .B(ori_ori_n49_), .Y(ori_ori_n53_));
  NO3        o0025(.A(ori_ori_n53_), .B(ori_ori_n48_), .C(ori_ori_n43_), .Y(ori_ori_n54_));
  AOI210     o0026(.A0(ori_ori_n54_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n55_));
  INV        o0027(.A(c), .Y(ori_ori_n56_));
  NA2        o0028(.A(e), .B(b), .Y(ori_ori_n57_));
  NO2        o0029(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0030(.A(d), .Y(ori_ori_n59_));
  NAi21      o0031(.An(i), .B(h), .Y(ori_ori_n60_));
  NAi41      o0032(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n61_));
  NA2        o0033(.A(g), .B(f), .Y(ori_ori_n62_));
  NO2        o0034(.A(ori_ori_n62_), .B(ori_ori_n61_), .Y(ori_ori_n63_));
  NAi21      o0035(.An(i), .B(j), .Y(ori_ori_n64_));
  NAi32      o0036(.An(n), .Bn(k), .C(m), .Y(ori_ori_n65_));
  NAi31      o0037(.An(l), .B(m), .C(k), .Y(ori_ori_n66_));
  NAi21      o0038(.An(e), .B(h), .Y(ori_ori_n67_));
  NAi41      o0039(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n68_));
  INV        o0040(.A(m), .Y(ori_ori_n69_));
  NOi21      o0041(.An(k), .B(l), .Y(ori_ori_n70_));
  NA2        o0042(.A(ori_ori_n70_), .B(ori_ori_n69_), .Y(ori_ori_n71_));
  AN4        o0043(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n72_));
  NOi31      o0044(.An(h), .B(g), .C(f), .Y(ori_ori_n73_));
  NA2        o0045(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  NAi32      o0046(.An(m), .Bn(k), .C(j), .Y(ori_ori_n75_));
  NOi32      o0047(.An(h), .Bn(g), .C(f), .Y(ori_ori_n76_));
  NA2        o0048(.A(ori_ori_n76_), .B(ori_ori_n72_), .Y(ori_ori_n77_));
  OA220      o0049(.A0(ori_ori_n77_), .A1(ori_ori_n75_), .B0(ori_ori_n74_), .B1(ori_ori_n71_), .Y(ori_ori_n78_));
  INV        o0050(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  INV        o0051(.A(n), .Y(ori_ori_n80_));
  NOi32      o0052(.An(e), .Bn(b), .C(d), .Y(ori_ori_n81_));
  NA2        o0053(.A(ori_ori_n81_), .B(ori_ori_n80_), .Y(ori_ori_n82_));
  INV        o0054(.A(j), .Y(ori_ori_n83_));
  AN3        o0055(.A(m), .B(k), .C(i), .Y(ori_ori_n84_));
  NA3        o0056(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(g), .Y(ori_ori_n85_));
  NO2        o0057(.A(ori_ori_n85_), .B(f), .Y(ori_ori_n86_));
  NAi32      o0058(.An(g), .Bn(f), .C(h), .Y(ori_ori_n87_));
  NAi31      o0059(.An(j), .B(m), .C(l), .Y(ori_ori_n88_));
  NO2        o0060(.A(ori_ori_n88_), .B(ori_ori_n87_), .Y(ori_ori_n89_));
  NA2        o0061(.A(m), .B(l), .Y(ori_ori_n90_));
  NAi31      o0062(.An(k), .B(j), .C(g), .Y(ori_ori_n91_));
  NO3        o0063(.A(ori_ori_n91_), .B(ori_ori_n90_), .C(f), .Y(ori_ori_n92_));
  AN2        o0064(.A(j), .B(g), .Y(ori_ori_n93_));
  NOi32      o0065(.An(m), .Bn(l), .C(i), .Y(ori_ori_n94_));
  NOi21      o0066(.An(g), .B(i), .Y(ori_ori_n95_));
  NOi32      o0067(.An(m), .Bn(j), .C(k), .Y(ori_ori_n96_));
  AOI220     o0068(.A0(ori_ori_n96_), .A1(ori_ori_n95_), .B0(ori_ori_n94_), .B1(ori_ori_n93_), .Y(ori_ori_n97_));
  NO2        o0069(.A(ori_ori_n97_), .B(f), .Y(ori_ori_n98_));
  NO4        o0070(.A(ori_ori_n98_), .B(ori_ori_n92_), .C(ori_ori_n89_), .D(ori_ori_n86_), .Y(ori_ori_n99_));
  NAi41      o0071(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n100_));
  AN2        o0072(.A(e), .B(b), .Y(ori_ori_n101_));
  NOi31      o0073(.An(c), .B(h), .C(f), .Y(ori_ori_n102_));
  NA2        o0074(.A(ori_ori_n102_), .B(ori_ori_n101_), .Y(ori_ori_n103_));
  NO2        o0075(.A(ori_ori_n103_), .B(ori_ori_n100_), .Y(ori_ori_n104_));
  NOi21      o0076(.An(i), .B(h), .Y(ori_ori_n105_));
  INV        o0077(.A(a), .Y(ori_ori_n106_));
  NA2        o0078(.A(ori_ori_n101_), .B(ori_ori_n106_), .Y(ori_ori_n107_));
  INV        o0079(.A(l), .Y(ori_ori_n108_));
  NOi21      o0080(.An(m), .B(n), .Y(ori_ori_n109_));
  AN2        o0081(.A(k), .B(h), .Y(ori_ori_n110_));
  INV        o0082(.A(b), .Y(ori_ori_n111_));
  NA2        o0083(.A(l), .B(j), .Y(ori_ori_n112_));
  AN2        o0084(.A(k), .B(i), .Y(ori_ori_n113_));
  NA2        o0085(.A(ori_ori_n113_), .B(ori_ori_n112_), .Y(ori_ori_n114_));
  NA2        o0086(.A(g), .B(e), .Y(ori_ori_n115_));
  NOi32      o0087(.An(c), .Bn(a), .C(d), .Y(ori_ori_n116_));
  NA2        o0088(.A(ori_ori_n116_), .B(ori_ori_n109_), .Y(ori_ori_n117_));
  INV        o0089(.A(ori_ori_n104_), .Y(ori_ori_n118_));
  OAI210     o0090(.A0(ori_ori_n99_), .A1(ori_ori_n82_), .B0(ori_ori_n118_), .Y(ori_ori_n119_));
  NOi31      o0091(.An(k), .B(m), .C(j), .Y(ori_ori_n120_));
  NA3        o0092(.A(ori_ori_n120_), .B(ori_ori_n73_), .C(ori_ori_n72_), .Y(ori_ori_n121_));
  NOi31      o0093(.An(k), .B(m), .C(i), .Y(ori_ori_n122_));
  NA3        o0094(.A(ori_ori_n122_), .B(ori_ori_n76_), .C(ori_ori_n72_), .Y(ori_ori_n123_));
  NA2        o0095(.A(ori_ori_n123_), .B(ori_ori_n121_), .Y(ori_ori_n124_));
  NOi32      o0096(.An(f), .Bn(b), .C(e), .Y(ori_ori_n125_));
  NAi21      o0097(.An(g), .B(h), .Y(ori_ori_n126_));
  NAi21      o0098(.An(m), .B(n), .Y(ori_ori_n127_));
  NAi41      o0099(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n128_));
  NAi31      o0100(.An(j), .B(k), .C(h), .Y(ori_ori_n129_));
  NO3        o0101(.A(ori_ori_n129_), .B(ori_ori_n128_), .C(ori_ori_n127_), .Y(ori_ori_n130_));
  INV        o0102(.A(ori_ori_n130_), .Y(ori_ori_n131_));
  NO2        o0103(.A(k), .B(j), .Y(ori_ori_n132_));
  NO2        o0104(.A(ori_ori_n132_), .B(ori_ori_n127_), .Y(ori_ori_n133_));
  AN2        o0105(.A(k), .B(j), .Y(ori_ori_n134_));
  NAi21      o0106(.An(c), .B(b), .Y(ori_ori_n135_));
  NA2        o0107(.A(f), .B(d), .Y(ori_ori_n136_));
  NO4        o0108(.A(ori_ori_n136_), .B(ori_ori_n135_), .C(ori_ori_n134_), .D(ori_ori_n126_), .Y(ori_ori_n137_));
  NA2        o0109(.A(h), .B(c), .Y(ori_ori_n138_));
  NAi31      o0110(.An(f), .B(e), .C(b), .Y(ori_ori_n139_));
  NA2        o0111(.A(ori_ori_n137_), .B(ori_ori_n133_), .Y(ori_ori_n140_));
  NA2        o0112(.A(d), .B(b), .Y(ori_ori_n141_));
  NAi21      o0113(.An(e), .B(f), .Y(ori_ori_n142_));
  NO2        o0114(.A(ori_ori_n142_), .B(ori_ori_n141_), .Y(ori_ori_n143_));
  NA2        o0115(.A(b), .B(a), .Y(ori_ori_n144_));
  NAi21      o0116(.An(e), .B(g), .Y(ori_ori_n145_));
  NAi21      o0117(.An(c), .B(d), .Y(ori_ori_n146_));
  NAi31      o0118(.An(l), .B(k), .C(h), .Y(ori_ori_n147_));
  NO2        o0119(.A(ori_ori_n127_), .B(ori_ori_n147_), .Y(ori_ori_n148_));
  NA2        o0120(.A(ori_ori_n148_), .B(ori_ori_n143_), .Y(ori_ori_n149_));
  NAi41      o0121(.An(ori_ori_n124_), .B(ori_ori_n149_), .C(ori_ori_n140_), .D(ori_ori_n131_), .Y(ori_ori_n150_));
  NAi31      o0122(.An(e), .B(f), .C(b), .Y(ori_ori_n151_));
  NOi21      o0123(.An(g), .B(d), .Y(ori_ori_n152_));
  NO2        o0124(.A(ori_ori_n152_), .B(ori_ori_n151_), .Y(ori_ori_n153_));
  NOi21      o0125(.An(h), .B(i), .Y(ori_ori_n154_));
  NOi21      o0126(.An(k), .B(m), .Y(ori_ori_n155_));
  NA3        o0127(.A(ori_ori_n155_), .B(ori_ori_n154_), .C(n), .Y(ori_ori_n156_));
  NOi21      o0128(.An(ori_ori_n153_), .B(ori_ori_n156_), .Y(ori_ori_n157_));
  NOi21      o0129(.An(h), .B(g), .Y(ori_ori_n158_));
  NO2        o0130(.A(ori_ori_n136_), .B(ori_ori_n135_), .Y(ori_ori_n159_));
  NAi31      o0131(.An(l), .B(j), .C(h), .Y(ori_ori_n160_));
  NO2        o0132(.A(ori_ori_n160_), .B(ori_ori_n49_), .Y(ori_ori_n161_));
  NA2        o0133(.A(ori_ori_n161_), .B(ori_ori_n63_), .Y(ori_ori_n162_));
  NOi32      o0134(.An(n), .Bn(k), .C(m), .Y(ori_ori_n163_));
  INV        o0135(.A(ori_ori_n162_), .Y(ori_ori_n164_));
  NAi31      o0136(.An(d), .B(f), .C(c), .Y(ori_ori_n165_));
  NAi31      o0137(.An(e), .B(f), .C(c), .Y(ori_ori_n166_));
  NA2        o0138(.A(ori_ori_n166_), .B(ori_ori_n165_), .Y(ori_ori_n167_));
  NA2        o0139(.A(j), .B(h), .Y(ori_ori_n168_));
  OR3        o0140(.A(n), .B(m), .C(k), .Y(ori_ori_n169_));
  NO2        o0141(.A(ori_ori_n169_), .B(ori_ori_n168_), .Y(ori_ori_n170_));
  NAi32      o0142(.An(m), .Bn(k), .C(n), .Y(ori_ori_n171_));
  NO2        o0143(.A(ori_ori_n171_), .B(ori_ori_n168_), .Y(ori_ori_n172_));
  AOI220     o0144(.A0(ori_ori_n172_), .A1(ori_ori_n153_), .B0(ori_ori_n170_), .B1(ori_ori_n167_), .Y(ori_ori_n173_));
  NO2        o0145(.A(n), .B(m), .Y(ori_ori_n174_));
  NA2        o0146(.A(ori_ori_n174_), .B(ori_ori_n50_), .Y(ori_ori_n175_));
  NAi21      o0147(.An(f), .B(e), .Y(ori_ori_n176_));
  NA2        o0148(.A(d), .B(c), .Y(ori_ori_n177_));
  NO2        o0149(.A(ori_ori_n177_), .B(ori_ori_n176_), .Y(ori_ori_n178_));
  NOi21      o0150(.An(ori_ori_n178_), .B(ori_ori_n175_), .Y(ori_ori_n179_));
  NAi31      o0151(.An(m), .B(n), .C(b), .Y(ori_ori_n180_));
  NA2        o0152(.A(k), .B(i), .Y(ori_ori_n181_));
  NAi21      o0153(.An(h), .B(f), .Y(ori_ori_n182_));
  NO2        o0154(.A(ori_ori_n182_), .B(ori_ori_n181_), .Y(ori_ori_n183_));
  NO2        o0155(.A(ori_ori_n180_), .B(ori_ori_n146_), .Y(ori_ori_n184_));
  NA2        o0156(.A(ori_ori_n184_), .B(ori_ori_n183_), .Y(ori_ori_n185_));
  NOi32      o0157(.An(f), .Bn(c), .C(d), .Y(ori_ori_n186_));
  NOi32      o0158(.An(f), .Bn(c), .C(e), .Y(ori_ori_n187_));
  NO2        o0159(.A(ori_ori_n187_), .B(ori_ori_n186_), .Y(ori_ori_n188_));
  NO3        o0160(.A(n), .B(m), .C(j), .Y(ori_ori_n189_));
  NA2        o0161(.A(ori_ori_n189_), .B(ori_ori_n110_), .Y(ori_ori_n190_));
  AO210      o0162(.A0(ori_ori_n190_), .A1(ori_ori_n175_), .B0(ori_ori_n188_), .Y(ori_ori_n191_));
  NAi41      o0163(.An(ori_ori_n179_), .B(ori_ori_n191_), .C(ori_ori_n185_), .D(ori_ori_n173_), .Y(ori_ori_n192_));
  OR4        o0164(.A(ori_ori_n192_), .B(ori_ori_n164_), .C(ori_ori_n157_), .D(ori_ori_n150_), .Y(ori_ori_n193_));
  NO4        o0165(.A(ori_ori_n193_), .B(ori_ori_n119_), .C(ori_ori_n79_), .D(ori_ori_n55_), .Y(ori_ori_n194_));
  NA3        o0166(.A(m), .B(ori_ori_n108_), .C(j), .Y(ori_ori_n195_));
  NAi31      o0167(.An(n), .B(h), .C(g), .Y(ori_ori_n196_));
  NO2        o0168(.A(ori_ori_n196_), .B(ori_ori_n195_), .Y(ori_ori_n197_));
  NOi32      o0169(.An(m), .Bn(k), .C(l), .Y(ori_ori_n198_));
  NA3        o0170(.A(ori_ori_n198_), .B(ori_ori_n83_), .C(g), .Y(ori_ori_n199_));
  NO2        o0171(.A(ori_ori_n199_), .B(n), .Y(ori_ori_n200_));
  NOi21      o0172(.An(k), .B(j), .Y(ori_ori_n201_));
  NA4        o0173(.A(ori_ori_n201_), .B(ori_ori_n109_), .C(i), .D(g), .Y(ori_ori_n202_));
  AN2        o0174(.A(i), .B(g), .Y(ori_ori_n203_));
  INV        o0175(.A(ori_ori_n202_), .Y(ori_ori_n204_));
  NO3        o0176(.A(ori_ori_n204_), .B(ori_ori_n200_), .C(ori_ori_n197_), .Y(ori_ori_n205_));
  NAi41      o0177(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n206_));
  INV        o0178(.A(ori_ori_n206_), .Y(ori_ori_n207_));
  INV        o0179(.A(f), .Y(ori_ori_n208_));
  INV        o0180(.A(g), .Y(ori_ori_n209_));
  NOi31      o0181(.An(i), .B(j), .C(h), .Y(ori_ori_n210_));
  NOi21      o0182(.An(l), .B(m), .Y(ori_ori_n211_));
  NA2        o0183(.A(ori_ori_n211_), .B(ori_ori_n210_), .Y(ori_ori_n212_));
  NO3        o0184(.A(ori_ori_n212_), .B(ori_ori_n209_), .C(ori_ori_n208_), .Y(ori_ori_n213_));
  NA2        o0185(.A(ori_ori_n213_), .B(ori_ori_n207_), .Y(ori_ori_n214_));
  OAI210     o0186(.A0(ori_ori_n205_), .A1(ori_ori_n32_), .B0(ori_ori_n214_), .Y(ori_ori_n215_));
  NOi21      o0187(.An(n), .B(m), .Y(ori_ori_n216_));
  NOi32      o0188(.An(l), .Bn(i), .C(j), .Y(ori_ori_n217_));
  NA2        o0189(.A(ori_ori_n217_), .B(ori_ori_n216_), .Y(ori_ori_n218_));
  OR2        o0190(.A(ori_ori_n75_), .B(ori_ori_n74_), .Y(ori_ori_n219_));
  NAi21      o0191(.An(j), .B(h), .Y(ori_ori_n220_));
  XN2        o0192(.A(i), .B(h), .Y(ori_ori_n221_));
  NA2        o0193(.A(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  NOi31      o0194(.An(k), .B(n), .C(m), .Y(ori_ori_n223_));
  NOi31      o0195(.An(ori_ori_n223_), .B(ori_ori_n177_), .C(ori_ori_n176_), .Y(ori_ori_n224_));
  NA2        o0196(.A(ori_ori_n224_), .B(ori_ori_n222_), .Y(ori_ori_n225_));
  NAi31      o0197(.An(f), .B(e), .C(c), .Y(ori_ori_n226_));
  NO4        o0198(.A(ori_ori_n226_), .B(ori_ori_n169_), .C(ori_ori_n168_), .D(ori_ori_n59_), .Y(ori_ori_n227_));
  NA3        o0199(.A(e), .B(c), .C(b), .Y(ori_ori_n228_));
  NAi32      o0200(.An(m), .Bn(i), .C(k), .Y(ori_ori_n229_));
  INV        o0201(.A(k), .Y(ori_ori_n230_));
  INV        o0202(.A(ori_ori_n227_), .Y(ori_ori_n231_));
  NAi21      o0203(.An(n), .B(a), .Y(ori_ori_n232_));
  NO2        o0204(.A(ori_ori_n232_), .B(ori_ori_n141_), .Y(ori_ori_n233_));
  NAi41      o0205(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n234_));
  NO2        o0206(.A(ori_ori_n234_), .B(e), .Y(ori_ori_n235_));
  NA2        o0207(.A(ori_ori_n235_), .B(ori_ori_n233_), .Y(ori_ori_n236_));
  AN4        o0208(.A(ori_ori_n236_), .B(ori_ori_n231_), .C(ori_ori_n225_), .D(ori_ori_n219_), .Y(ori_ori_n237_));
  OR2        o0209(.A(h), .B(g), .Y(ori_ori_n238_));
  NO2        o0210(.A(ori_ori_n238_), .B(ori_ori_n100_), .Y(ori_ori_n239_));
  NA2        o0211(.A(ori_ori_n239_), .B(ori_ori_n125_), .Y(ori_ori_n240_));
  NAi41      o0212(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n241_));
  NO2        o0213(.A(ori_ori_n241_), .B(ori_ori_n208_), .Y(ori_ori_n242_));
  NA2        o0214(.A(ori_ori_n155_), .B(ori_ori_n105_), .Y(ori_ori_n243_));
  NAi21      o0215(.An(ori_ori_n243_), .B(ori_ori_n242_), .Y(ori_ori_n244_));
  NO2        o0216(.A(n), .B(a), .Y(ori_ori_n245_));
  NAi31      o0217(.An(ori_ori_n234_), .B(ori_ori_n245_), .C(ori_ori_n101_), .Y(ori_ori_n246_));
  AN2        o0218(.A(ori_ori_n246_), .B(ori_ori_n244_), .Y(ori_ori_n247_));
  NAi21      o0219(.An(h), .B(i), .Y(ori_ori_n248_));
  NA2        o0220(.A(ori_ori_n174_), .B(k), .Y(ori_ori_n249_));
  NO2        o0221(.A(ori_ori_n249_), .B(ori_ori_n248_), .Y(ori_ori_n250_));
  NA2        o0222(.A(ori_ori_n250_), .B(ori_ori_n186_), .Y(ori_ori_n251_));
  NA3        o0223(.A(ori_ori_n251_), .B(ori_ori_n247_), .C(ori_ori_n240_), .Y(ori_ori_n252_));
  NOi21      o0224(.An(g), .B(e), .Y(ori_ori_n253_));
  NO2        o0225(.A(ori_ori_n68_), .B(ori_ori_n69_), .Y(ori_ori_n254_));
  NA2        o0226(.A(ori_ori_n254_), .B(ori_ori_n253_), .Y(ori_ori_n255_));
  NOi32      o0227(.An(l), .Bn(j), .C(i), .Y(ori_ori_n256_));
  AOI210     o0228(.A0(ori_ori_n70_), .A1(ori_ori_n83_), .B0(ori_ori_n256_), .Y(ori_ori_n257_));
  NO2        o0229(.A(ori_ori_n248_), .B(ori_ori_n44_), .Y(ori_ori_n258_));
  NAi21      o0230(.An(f), .B(g), .Y(ori_ori_n259_));
  NO2        o0231(.A(ori_ori_n259_), .B(ori_ori_n61_), .Y(ori_ori_n260_));
  NO2        o0232(.A(ori_ori_n65_), .B(ori_ori_n112_), .Y(ori_ori_n261_));
  AOI220     o0233(.A0(ori_ori_n261_), .A1(ori_ori_n260_), .B0(ori_ori_n258_), .B1(ori_ori_n63_), .Y(ori_ori_n262_));
  OAI210     o0234(.A0(ori_ori_n257_), .A1(ori_ori_n255_), .B0(ori_ori_n262_), .Y(ori_ori_n263_));
  NOi41      o0235(.An(ori_ori_n237_), .B(ori_ori_n263_), .C(ori_ori_n252_), .D(ori_ori_n215_), .Y(ori_ori_n264_));
  NO4        o0236(.A(ori_ori_n197_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n265_));
  NO2        o0237(.A(ori_ori_n265_), .B(ori_ori_n107_), .Y(ori_ori_n266_));
  NA3        o0238(.A(ori_ori_n59_), .B(c), .C(b), .Y(ori_ori_n267_));
  NAi21      o0239(.An(h), .B(g), .Y(ori_ori_n268_));
  OR4        o0240(.A(ori_ori_n268_), .B(ori_ori_n267_), .C(ori_ori_n218_), .D(e), .Y(ori_ori_n269_));
  NO2        o0241(.A(ori_ori_n243_), .B(ori_ori_n259_), .Y(ori_ori_n270_));
  NAi31      o0242(.An(g), .B(k), .C(h), .Y(ori_ori_n271_));
  NO3        o0243(.A(ori_ori_n127_), .B(ori_ori_n271_), .C(l), .Y(ori_ori_n272_));
  NAi31      o0244(.An(e), .B(d), .C(a), .Y(ori_ori_n273_));
  NA2        o0245(.A(ori_ori_n272_), .B(ori_ori_n125_), .Y(ori_ori_n274_));
  NA2        o0246(.A(ori_ori_n274_), .B(ori_ori_n269_), .Y(ori_ori_n275_));
  NA4        o0247(.A(ori_ori_n155_), .B(ori_ori_n76_), .C(ori_ori_n72_), .D(ori_ori_n112_), .Y(ori_ori_n276_));
  NA3        o0248(.A(ori_ori_n155_), .B(ori_ori_n154_), .C(ori_ori_n80_), .Y(ori_ori_n277_));
  NO2        o0249(.A(ori_ori_n277_), .B(ori_ori_n188_), .Y(ori_ori_n278_));
  NOi21      o0250(.An(ori_ori_n276_), .B(ori_ori_n278_), .Y(ori_ori_n279_));
  NA3        o0251(.A(e), .B(c), .C(b), .Y(ori_ori_n280_));
  NAi32      o0252(.An(k), .Bn(i), .C(j), .Y(ori_ori_n281_));
  NAi31      o0253(.An(h), .B(l), .C(i), .Y(ori_ori_n282_));
  NA3        o0254(.A(ori_ori_n282_), .B(ori_ori_n281_), .C(ori_ori_n160_), .Y(ori_ori_n283_));
  NOi21      o0255(.An(ori_ori_n283_), .B(ori_ori_n49_), .Y(ori_ori_n284_));
  NA2        o0256(.A(ori_ori_n260_), .B(ori_ori_n284_), .Y(ori_ori_n285_));
  NAi21      o0257(.An(l), .B(k), .Y(ori_ori_n286_));
  NO2        o0258(.A(ori_ori_n286_), .B(ori_ori_n49_), .Y(ori_ori_n287_));
  NOi21      o0259(.An(l), .B(j), .Y(ori_ori_n288_));
  NA2        o0260(.A(ori_ori_n158_), .B(ori_ori_n288_), .Y(ori_ori_n289_));
  NAi32      o0261(.An(j), .Bn(h), .C(i), .Y(ori_ori_n290_));
  NAi21      o0262(.An(m), .B(l), .Y(ori_ori_n291_));
  NO3        o0263(.A(ori_ori_n291_), .B(ori_ori_n290_), .C(ori_ori_n80_), .Y(ori_ori_n292_));
  NA2        o0264(.A(h), .B(g), .Y(ori_ori_n293_));
  NA2        o0265(.A(ori_ori_n163_), .B(ori_ori_n45_), .Y(ori_ori_n294_));
  NO2        o0266(.A(ori_ori_n294_), .B(ori_ori_n293_), .Y(ori_ori_n295_));
  OAI210     o0267(.A0(ori_ori_n295_), .A1(ori_ori_n292_), .B0(ori_ori_n159_), .Y(ori_ori_n296_));
  NA3        o0268(.A(ori_ori_n296_), .B(ori_ori_n285_), .C(ori_ori_n279_), .Y(ori_ori_n297_));
  NO2        o0269(.A(ori_ori_n139_), .B(d), .Y(ori_ori_n298_));
  NA2        o0270(.A(ori_ori_n298_), .B(ori_ori_n53_), .Y(ori_ori_n299_));
  NO2        o0271(.A(ori_ori_n103_), .B(ori_ori_n100_), .Y(ori_ori_n300_));
  NAi32      o0272(.An(n), .Bn(m), .C(l), .Y(ori_ori_n301_));
  NO2        o0273(.A(ori_ori_n301_), .B(ori_ori_n290_), .Y(ori_ori_n302_));
  NA2        o0274(.A(ori_ori_n302_), .B(ori_ori_n178_), .Y(ori_ori_n303_));
  NAi31      o0275(.An(k), .B(l), .C(j), .Y(ori_ori_n304_));
  OAI210     o0276(.A0(ori_ori_n286_), .A1(j), .B0(ori_ori_n304_), .Y(ori_ori_n305_));
  NOi21      o0277(.An(ori_ori_n305_), .B(ori_ori_n115_), .Y(ori_ori_n306_));
  NA2        o0278(.A(ori_ori_n303_), .B(ori_ori_n299_), .Y(ori_ori_n307_));
  NO4        o0279(.A(ori_ori_n307_), .B(ori_ori_n297_), .C(ori_ori_n275_), .D(ori_ori_n266_), .Y(ori_ori_n308_));
  NA2        o0280(.A(ori_ori_n250_), .B(ori_ori_n187_), .Y(ori_ori_n309_));
  NAi21      o0281(.An(m), .B(k), .Y(ori_ori_n310_));
  NO2        o0282(.A(ori_ori_n221_), .B(ori_ori_n310_), .Y(ori_ori_n311_));
  NAi41      o0283(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n312_));
  NO2        o0284(.A(ori_ori_n312_), .B(ori_ori_n145_), .Y(ori_ori_n313_));
  NA2        o0285(.A(ori_ori_n313_), .B(ori_ori_n311_), .Y(ori_ori_n314_));
  NAi31      o0286(.An(i), .B(l), .C(h), .Y(ori_ori_n315_));
  NO4        o0287(.A(ori_ori_n315_), .B(ori_ori_n145_), .C(ori_ori_n68_), .D(ori_ori_n69_), .Y(ori_ori_n316_));
  NA2        o0288(.A(e), .B(c), .Y(ori_ori_n317_));
  NO3        o0289(.A(ori_ori_n317_), .B(n), .C(d), .Y(ori_ori_n318_));
  NOi21      o0290(.An(f), .B(h), .Y(ori_ori_n319_));
  NAi31      o0291(.An(d), .B(e), .C(b), .Y(ori_ori_n320_));
  NAi31      o0292(.An(ori_ori_n316_), .B(ori_ori_n314_), .C(ori_ori_n309_), .Y(ori_ori_n321_));
  NO4        o0293(.A(ori_ori_n312_), .B(ori_ori_n75_), .C(ori_ori_n67_), .D(ori_ori_n209_), .Y(ori_ori_n322_));
  NA2        o0294(.A(ori_ori_n245_), .B(ori_ori_n101_), .Y(ori_ori_n323_));
  OR2        o0295(.A(ori_ori_n323_), .B(ori_ori_n199_), .Y(ori_ori_n324_));
  NOi31      o0296(.An(l), .B(n), .C(m), .Y(ori_ori_n325_));
  NA2        o0297(.A(ori_ori_n325_), .B(ori_ori_n210_), .Y(ori_ori_n326_));
  NO2        o0298(.A(ori_ori_n326_), .B(ori_ori_n188_), .Y(ori_ori_n327_));
  NAi32      o0299(.An(ori_ori_n327_), .Bn(ori_ori_n322_), .C(ori_ori_n324_), .Y(ori_ori_n328_));
  NAi32      o0300(.An(m), .Bn(j), .C(k), .Y(ori_ori_n329_));
  NAi41      o0301(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n330_));
  OAI210     o0302(.A0(ori_ori_n206_), .A1(ori_ori_n329_), .B0(ori_ori_n330_), .Y(ori_ori_n331_));
  NOi31      o0303(.An(j), .B(m), .C(k), .Y(ori_ori_n332_));
  NO2        o0304(.A(ori_ori_n120_), .B(ori_ori_n332_), .Y(ori_ori_n333_));
  AN3        o0305(.A(h), .B(g), .C(f), .Y(ori_ori_n334_));
  NAi31      o0306(.An(ori_ori_n333_), .B(ori_ori_n334_), .C(ori_ori_n331_), .Y(ori_ori_n335_));
  NOi32      o0307(.An(m), .Bn(j), .C(l), .Y(ori_ori_n336_));
  NO2        o0308(.A(ori_ori_n336_), .B(ori_ori_n94_), .Y(ori_ori_n337_));
  NAi32      o0309(.An(ori_ori_n337_), .Bn(ori_ori_n196_), .C(ori_ori_n298_), .Y(ori_ori_n338_));
  NO2        o0310(.A(ori_ori_n291_), .B(ori_ori_n290_), .Y(ori_ori_n339_));
  NO2        o0311(.A(ori_ori_n212_), .B(g), .Y(ori_ori_n340_));
  NO2        o0312(.A(ori_ori_n151_), .B(ori_ori_n80_), .Y(ori_ori_n341_));
  AOI220     o0313(.A0(ori_ori_n341_), .A1(ori_ori_n340_), .B0(ori_ori_n242_), .B1(ori_ori_n339_), .Y(ori_ori_n342_));
  NA2        o0314(.A(ori_ori_n229_), .B(ori_ori_n75_), .Y(ori_ori_n343_));
  NA3        o0315(.A(ori_ori_n343_), .B(ori_ori_n334_), .C(ori_ori_n207_), .Y(ori_ori_n344_));
  NA4        o0316(.A(ori_ori_n344_), .B(ori_ori_n342_), .C(ori_ori_n338_), .D(ori_ori_n335_), .Y(ori_ori_n345_));
  NA3        o0317(.A(h), .B(g), .C(f), .Y(ori_ori_n346_));
  NO2        o0318(.A(ori_ori_n346_), .B(ori_ori_n71_), .Y(ori_ori_n347_));
  NA2        o0319(.A(ori_ori_n158_), .B(e), .Y(ori_ori_n348_));
  NO2        o0320(.A(ori_ori_n348_), .B(ori_ori_n41_), .Y(ori_ori_n349_));
  NOi32      o0321(.An(j), .Bn(g), .C(i), .Y(ori_ori_n350_));
  NA3        o0322(.A(ori_ori_n350_), .B(ori_ori_n286_), .C(ori_ori_n109_), .Y(ori_ori_n351_));
  AO210      o0323(.A0(ori_ori_n107_), .A1(ori_ori_n32_), .B0(ori_ori_n351_), .Y(ori_ori_n352_));
  NOi32      o0324(.An(e), .Bn(b), .C(a), .Y(ori_ori_n353_));
  AN2        o0325(.A(l), .B(j), .Y(ori_ori_n354_));
  NO2        o0326(.A(ori_ori_n310_), .B(ori_ori_n354_), .Y(ori_ori_n355_));
  NO3        o0327(.A(ori_ori_n312_), .B(ori_ori_n67_), .C(ori_ori_n209_), .Y(ori_ori_n356_));
  NA2        o0328(.A(ori_ori_n202_), .B(ori_ori_n35_), .Y(ori_ori_n357_));
  AOI220     o0329(.A0(ori_ori_n357_), .A1(ori_ori_n353_), .B0(ori_ori_n356_), .B1(ori_ori_n355_), .Y(ori_ori_n358_));
  NO2        o0330(.A(ori_ori_n320_), .B(n), .Y(ori_ori_n359_));
  NA2        o0331(.A(ori_ori_n203_), .B(k), .Y(ori_ori_n360_));
  NA3        o0332(.A(m), .B(ori_ori_n108_), .C(ori_ori_n208_), .Y(ori_ori_n361_));
  NA4        o0333(.A(ori_ori_n198_), .B(ori_ori_n83_), .C(g), .D(ori_ori_n208_), .Y(ori_ori_n362_));
  OAI210     o0334(.A0(ori_ori_n361_), .A1(ori_ori_n360_), .B0(ori_ori_n362_), .Y(ori_ori_n363_));
  NAi41      o0335(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n364_));
  NA2        o0336(.A(ori_ori_n51_), .B(ori_ori_n109_), .Y(ori_ori_n365_));
  NO2        o0337(.A(ori_ori_n365_), .B(ori_ori_n364_), .Y(ori_ori_n366_));
  NA2        o0338(.A(ori_ori_n363_), .B(ori_ori_n359_), .Y(ori_ori_n367_));
  NA3        o0339(.A(ori_ori_n367_), .B(ori_ori_n358_), .C(ori_ori_n352_), .Y(ori_ori_n368_));
  NO4        o0340(.A(ori_ori_n368_), .B(ori_ori_n345_), .C(ori_ori_n328_), .D(ori_ori_n321_), .Y(ori_ori_n369_));
  NA4        o0341(.A(ori_ori_n369_), .B(ori_ori_n308_), .C(ori_ori_n264_), .D(ori_ori_n194_), .Y(ori10));
  NA3        o0342(.A(m), .B(k), .C(i), .Y(ori_ori_n371_));
  NOi21      o0343(.An(e), .B(f), .Y(ori_ori_n372_));
  NAi31      o0344(.An(b), .B(f), .C(c), .Y(ori_ori_n373_));
  INV        o0345(.A(ori_ori_n373_), .Y(ori_ori_n374_));
  NOi32      o0346(.An(k), .Bn(h), .C(j), .Y(ori_ori_n375_));
  NA2        o0347(.A(ori_ori_n375_), .B(ori_ori_n216_), .Y(ori_ori_n376_));
  NA2        o0348(.A(ori_ori_n156_), .B(ori_ori_n376_), .Y(ori_ori_n377_));
  NA2        o0349(.A(ori_ori_n377_), .B(ori_ori_n374_), .Y(ori_ori_n378_));
  AN2        o0350(.A(j), .B(h), .Y(ori_ori_n379_));
  NO3        o0351(.A(n), .B(m), .C(k), .Y(ori_ori_n380_));
  NA2        o0352(.A(ori_ori_n380_), .B(ori_ori_n379_), .Y(ori_ori_n381_));
  NO3        o0353(.A(ori_ori_n381_), .B(ori_ori_n146_), .C(ori_ori_n208_), .Y(ori_ori_n382_));
  OR2        o0354(.A(m), .B(k), .Y(ori_ori_n383_));
  NO2        o0355(.A(ori_ori_n168_), .B(ori_ori_n383_), .Y(ori_ori_n384_));
  NA4        o0356(.A(n), .B(f), .C(c), .D(ori_ori_n111_), .Y(ori_ori_n385_));
  NOi21      o0357(.An(ori_ori_n384_), .B(ori_ori_n385_), .Y(ori_ori_n386_));
  NOi32      o0358(.An(d), .Bn(a), .C(c), .Y(ori_ori_n387_));
  NA2        o0359(.A(ori_ori_n387_), .B(ori_ori_n176_), .Y(ori_ori_n388_));
  NAi21      o0360(.An(i), .B(g), .Y(ori_ori_n389_));
  NAi31      o0361(.An(k), .B(m), .C(j), .Y(ori_ori_n390_));
  NO3        o0362(.A(ori_ori_n390_), .B(ori_ori_n389_), .C(n), .Y(ori_ori_n391_));
  NOi21      o0363(.An(ori_ori_n391_), .B(ori_ori_n388_), .Y(ori_ori_n392_));
  NO3        o0364(.A(ori_ori_n392_), .B(ori_ori_n386_), .C(ori_ori_n382_), .Y(ori_ori_n393_));
  NO2        o0365(.A(ori_ori_n385_), .B(ori_ori_n291_), .Y(ori_ori_n394_));
  NOi32      o0366(.An(f), .Bn(d), .C(c), .Y(ori_ori_n395_));
  AOI220     o0367(.A0(ori_ori_n395_), .A1(ori_ori_n302_), .B0(ori_ori_n394_), .B1(ori_ori_n210_), .Y(ori_ori_n396_));
  NA3        o0368(.A(ori_ori_n396_), .B(ori_ori_n393_), .C(ori_ori_n378_), .Y(ori_ori_n397_));
  NO2        o0369(.A(ori_ori_n59_), .B(ori_ori_n111_), .Y(ori_ori_n398_));
  NA2        o0370(.A(ori_ori_n245_), .B(ori_ori_n398_), .Y(ori_ori_n399_));
  INV        o0371(.A(e), .Y(ori_ori_n400_));
  NA2        o0372(.A(ori_ori_n46_), .B(e), .Y(ori_ori_n401_));
  OAI220     o0373(.A0(ori_ori_n401_), .A1(ori_ori_n195_), .B0(ori_ori_n199_), .B1(ori_ori_n400_), .Y(ori_ori_n402_));
  NO2        o0374(.A(ori_ori_n85_), .B(ori_ori_n400_), .Y(ori_ori_n403_));
  NO2        o0375(.A(ori_ori_n97_), .B(ori_ori_n400_), .Y(ori_ori_n404_));
  NO3        o0376(.A(ori_ori_n404_), .B(ori_ori_n403_), .C(ori_ori_n402_), .Y(ori_ori_n405_));
  NOi32      o0377(.An(h), .Bn(e), .C(g), .Y(ori_ori_n406_));
  NA3        o0378(.A(ori_ori_n406_), .B(ori_ori_n288_), .C(m), .Y(ori_ori_n407_));
  NOi21      o0379(.An(g), .B(h), .Y(ori_ori_n408_));
  AN3        o0380(.A(m), .B(l), .C(i), .Y(ori_ori_n409_));
  NA3        o0381(.A(ori_ori_n409_), .B(ori_ori_n408_), .C(e), .Y(ori_ori_n410_));
  AN3        o0382(.A(h), .B(g), .C(e), .Y(ori_ori_n411_));
  NA2        o0383(.A(ori_ori_n411_), .B(ori_ori_n94_), .Y(ori_ori_n412_));
  AN3        o0384(.A(ori_ori_n412_), .B(ori_ori_n410_), .C(ori_ori_n407_), .Y(ori_ori_n413_));
  AOI210     o0385(.A0(ori_ori_n413_), .A1(ori_ori_n405_), .B0(ori_ori_n399_), .Y(ori_ori_n414_));
  NA3        o0386(.A(ori_ori_n387_), .B(ori_ori_n176_), .C(ori_ori_n80_), .Y(ori_ori_n415_));
  NAi31      o0387(.An(b), .B(c), .C(a), .Y(ori_ori_n416_));
  NO2        o0388(.A(ori_ori_n416_), .B(n), .Y(ori_ori_n417_));
  NA2        o0389(.A(ori_ori_n51_), .B(m), .Y(ori_ori_n418_));
  NO2        o0390(.A(ori_ori_n418_), .B(ori_ori_n142_), .Y(ori_ori_n419_));
  NO2        o0391(.A(ori_ori_n414_), .B(ori_ori_n397_), .Y(ori_ori_n420_));
  NA2        o0392(.A(i), .B(g), .Y(ori_ori_n421_));
  NOi21      o0393(.An(a), .B(n), .Y(ori_ori_n422_));
  NOi21      o0394(.An(d), .B(c), .Y(ori_ori_n423_));
  NA2        o0395(.A(ori_ori_n423_), .B(ori_ori_n422_), .Y(ori_ori_n424_));
  NA3        o0396(.A(i), .B(g), .C(f), .Y(ori_ori_n425_));
  OR2        o0397(.A(n), .B(m), .Y(ori_ori_n426_));
  NO2        o0398(.A(ori_ori_n426_), .B(ori_ori_n147_), .Y(ori_ori_n427_));
  NO2        o0399(.A(ori_ori_n177_), .B(ori_ori_n142_), .Y(ori_ori_n428_));
  OAI210     o0400(.A0(ori_ori_n427_), .A1(ori_ori_n170_), .B0(ori_ori_n428_), .Y(ori_ori_n429_));
  INV        o0401(.A(ori_ori_n365_), .Y(ori_ori_n430_));
  NA3        o0402(.A(ori_ori_n430_), .B(ori_ori_n353_), .C(d), .Y(ori_ori_n431_));
  NO2        o0403(.A(ori_ori_n416_), .B(ori_ori_n49_), .Y(ori_ori_n432_));
  NAi21      o0404(.An(k), .B(j), .Y(ori_ori_n433_));
  NAi21      o0405(.An(e), .B(d), .Y(ori_ori_n434_));
  INV        o0406(.A(ori_ori_n434_), .Y(ori_ori_n435_));
  NO2        o0407(.A(ori_ori_n249_), .B(ori_ori_n208_), .Y(ori_ori_n436_));
  NA3        o0408(.A(ori_ori_n436_), .B(ori_ori_n435_), .C(ori_ori_n222_), .Y(ori_ori_n437_));
  NA3        o0409(.A(ori_ori_n437_), .B(ori_ori_n431_), .C(ori_ori_n429_), .Y(ori_ori_n438_));
  NO2        o0410(.A(ori_ori_n326_), .B(ori_ori_n208_), .Y(ori_ori_n439_));
  NA2        o0411(.A(ori_ori_n439_), .B(ori_ori_n435_), .Y(ori_ori_n440_));
  NOi31      o0412(.An(n), .B(m), .C(k), .Y(ori_ori_n441_));
  AOI220     o0413(.A0(ori_ori_n441_), .A1(ori_ori_n379_), .B0(ori_ori_n216_), .B1(ori_ori_n50_), .Y(ori_ori_n442_));
  NAi31      o0414(.An(g), .B(f), .C(c), .Y(ori_ori_n443_));
  OR3        o0415(.A(ori_ori_n443_), .B(ori_ori_n442_), .C(e), .Y(ori_ori_n444_));
  NA3        o0416(.A(ori_ori_n444_), .B(ori_ori_n440_), .C(ori_ori_n303_), .Y(ori_ori_n445_));
  NO3        o0417(.A(ori_ori_n445_), .B(ori_ori_n438_), .C(ori_ori_n263_), .Y(ori_ori_n446_));
  NOi32      o0418(.An(c), .Bn(a), .C(b), .Y(ori_ori_n447_));
  NA2        o0419(.A(ori_ori_n447_), .B(ori_ori_n109_), .Y(ori_ori_n448_));
  INV        o0420(.A(ori_ori_n271_), .Y(ori_ori_n449_));
  AN2        o0421(.A(e), .B(d), .Y(ori_ori_n450_));
  INV        o0422(.A(ori_ori_n142_), .Y(ori_ori_n451_));
  NO2        o0423(.A(ori_ori_n126_), .B(ori_ori_n41_), .Y(ori_ori_n452_));
  NO2        o0424(.A(ori_ori_n62_), .B(e), .Y(ori_ori_n453_));
  NOi31      o0425(.An(j), .B(k), .C(i), .Y(ori_ori_n454_));
  NOi21      o0426(.An(ori_ori_n160_), .B(ori_ori_n454_), .Y(ori_ori_n455_));
  NA3        o0427(.A(ori_ori_n455_), .B(ori_ori_n257_), .C(ori_ori_n114_), .Y(ori_ori_n456_));
  AOI220     o0428(.A0(ori_ori_n456_), .A1(ori_ori_n453_), .B0(ori_ori_n452_), .B1(ori_ori_n451_), .Y(ori_ori_n457_));
  NO2        o0429(.A(ori_ori_n457_), .B(ori_ori_n448_), .Y(ori_ori_n458_));
  NO2        o0430(.A(ori_ori_n204_), .B(ori_ori_n200_), .Y(ori_ori_n459_));
  NOi21      o0431(.An(a), .B(b), .Y(ori_ori_n460_));
  NA3        o0432(.A(e), .B(d), .C(c), .Y(ori_ori_n461_));
  NAi21      o0433(.An(ori_ori_n461_), .B(ori_ori_n460_), .Y(ori_ori_n462_));
  NO2        o0434(.A(ori_ori_n415_), .B(ori_ori_n199_), .Y(ori_ori_n463_));
  NOi21      o0435(.An(ori_ori_n462_), .B(ori_ori_n463_), .Y(ori_ori_n464_));
  AOI210     o0436(.A0(ori_ori_n265_), .A1(ori_ori_n459_), .B0(ori_ori_n464_), .Y(ori_ori_n465_));
  NO4        o0437(.A(ori_ori_n182_), .B(ori_ori_n100_), .C(ori_ori_n56_), .D(b), .Y(ori_ori_n466_));
  NA2        o0438(.A(ori_ori_n374_), .B(ori_ori_n148_), .Y(ori_ori_n467_));
  OR2        o0439(.A(k), .B(j), .Y(ori_ori_n468_));
  NA2        o0440(.A(l), .B(k), .Y(ori_ori_n469_));
  NA3        o0441(.A(ori_ori_n469_), .B(ori_ori_n468_), .C(ori_ori_n216_), .Y(ori_ori_n470_));
  AOI210     o0442(.A0(ori_ori_n229_), .A1(ori_ori_n329_), .B0(ori_ori_n80_), .Y(ori_ori_n471_));
  NOi21      o0443(.An(ori_ori_n470_), .B(ori_ori_n471_), .Y(ori_ori_n472_));
  OR3        o0444(.A(ori_ori_n472_), .B(ori_ori_n138_), .C(ori_ori_n128_), .Y(ori_ori_n473_));
  NA3        o0445(.A(ori_ori_n276_), .B(ori_ori_n123_), .C(ori_ori_n121_), .Y(ori_ori_n474_));
  NO3        o0446(.A(ori_ori_n415_), .B(ori_ori_n88_), .C(ori_ori_n126_), .Y(ori_ori_n475_));
  NO3        o0447(.A(ori_ori_n475_), .B(ori_ori_n474_), .C(ori_ori_n316_), .Y(ori_ori_n476_));
  NA3        o0448(.A(ori_ori_n476_), .B(ori_ori_n473_), .C(ori_ori_n467_), .Y(ori_ori_n477_));
  NO4        o0449(.A(ori_ori_n477_), .B(ori_ori_n466_), .C(ori_ori_n465_), .D(ori_ori_n458_), .Y(ori_ori_n478_));
  INV        o0450(.A(e), .Y(ori_ori_n479_));
  NO2        o0451(.A(ori_ori_n182_), .B(ori_ori_n56_), .Y(ori_ori_n480_));
  NAi31      o0452(.An(j), .B(l), .C(i), .Y(ori_ori_n481_));
  OAI210     o0453(.A0(ori_ori_n481_), .A1(ori_ori_n127_), .B0(ori_ori_n100_), .Y(ori_ori_n482_));
  NA3        o0454(.A(ori_ori_n482_), .B(ori_ori_n480_), .C(ori_ori_n479_), .Y(ori_ori_n483_));
  NO3        o0455(.A(ori_ori_n388_), .B(ori_ori_n337_), .C(ori_ori_n196_), .Y(ori_ori_n484_));
  NO2        o0456(.A(ori_ori_n388_), .B(ori_ori_n365_), .Y(ori_ori_n485_));
  NO4        o0457(.A(ori_ori_n485_), .B(ori_ori_n484_), .C(ori_ori_n179_), .D(ori_ori_n300_), .Y(ori_ori_n486_));
  NA3        o0458(.A(ori_ori_n486_), .B(ori_ori_n483_), .C(ori_ori_n237_), .Y(ori_ori_n487_));
  OAI210     o0459(.A0(ori_ori_n122_), .A1(ori_ori_n120_), .B0(n), .Y(ori_ori_n488_));
  NO2        o0460(.A(ori_ori_n488_), .B(ori_ori_n126_), .Y(ori_ori_n489_));
  XO2        o0461(.A(i), .B(h), .Y(ori_ori_n490_));
  NA3        o0462(.A(ori_ori_n490_), .B(ori_ori_n155_), .C(n), .Y(ori_ori_n491_));
  NAi41      o0463(.An(ori_ori_n292_), .B(ori_ori_n491_), .C(ori_ori_n442_), .D(ori_ori_n376_), .Y(ori_ori_n492_));
  NOi32      o0464(.An(ori_ori_n492_), .Bn(ori_ori_n453_), .C(ori_ori_n267_), .Y(ori_ori_n493_));
  NAi31      o0465(.An(c), .B(f), .C(d), .Y(ori_ori_n494_));
  AOI210     o0466(.A0(ori_ori_n277_), .A1(ori_ori_n190_), .B0(ori_ori_n494_), .Y(ori_ori_n495_));
  NOi21      o0467(.An(ori_ori_n78_), .B(ori_ori_n495_), .Y(ori_ori_n496_));
  NA2        o0468(.A(ori_ori_n223_), .B(ori_ori_n105_), .Y(ori_ori_n497_));
  AOI210     o0469(.A0(ori_ori_n497_), .A1(ori_ori_n175_), .B0(ori_ori_n494_), .Y(ori_ori_n498_));
  INV        o0470(.A(ori_ori_n498_), .Y(ori_ori_n499_));
  AO220      o0471(.A0(ori_ori_n284_), .A1(ori_ori_n260_), .B0(ori_ori_n161_), .B1(ori_ori_n63_), .Y(ori_ori_n500_));
  NA3        o0472(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(f), .Y(ori_ori_n501_));
  NO2        o0473(.A(ori_ori_n501_), .B(ori_ori_n424_), .Y(ori_ori_n502_));
  INV        o0474(.A(ori_ori_n502_), .Y(ori_ori_n503_));
  NAi41      o0475(.An(ori_ori_n500_), .B(ori_ori_n503_), .C(ori_ori_n499_), .D(ori_ori_n496_), .Y(ori_ori_n504_));
  NO3        o0476(.A(ori_ori_n504_), .B(ori_ori_n493_), .C(ori_ori_n487_), .Y(ori_ori_n505_));
  NA4        o0477(.A(ori_ori_n505_), .B(ori_ori_n478_), .C(ori_ori_n446_), .D(ori_ori_n420_), .Y(ori11));
  NO2        o0478(.A(ori_ori_n68_), .B(f), .Y(ori_ori_n507_));
  NA2        o0479(.A(j), .B(g), .Y(ori_ori_n508_));
  NAi31      o0480(.An(i), .B(m), .C(l), .Y(ori_ori_n509_));
  NA3        o0481(.A(m), .B(k), .C(j), .Y(ori_ori_n510_));
  OAI220     o0482(.A0(ori_ori_n510_), .A1(ori_ori_n126_), .B0(ori_ori_n509_), .B1(ori_ori_n508_), .Y(ori_ori_n511_));
  NA2        o0483(.A(ori_ori_n511_), .B(ori_ori_n507_), .Y(ori_ori_n512_));
  NOi32      o0484(.An(e), .Bn(b), .C(f), .Y(ori_ori_n513_));
  NA2        o0485(.A(ori_ori_n46_), .B(j), .Y(ori_ori_n514_));
  NO2        o0486(.A(ori_ori_n514_), .B(ori_ori_n294_), .Y(ori_ori_n515_));
  NAi31      o0487(.An(d), .B(e), .C(a), .Y(ori_ori_n516_));
  NO2        o0488(.A(ori_ori_n516_), .B(n), .Y(ori_ori_n517_));
  AOI220     o0489(.A0(ori_ori_n517_), .A1(ori_ori_n98_), .B0(ori_ori_n515_), .B1(ori_ori_n513_), .Y(ori_ori_n518_));
  NAi41      o0490(.An(f), .B(e), .C(c), .D(a), .Y(ori_ori_n519_));
  AN2        o0491(.A(ori_ori_n519_), .B(ori_ori_n364_), .Y(ori_ori_n520_));
  NA2        o0492(.A(j), .B(i), .Y(ori_ori_n521_));
  NAi31      o0493(.An(n), .B(m), .C(k), .Y(ori_ori_n522_));
  NO3        o0494(.A(ori_ori_n522_), .B(ori_ori_n521_), .C(ori_ori_n108_), .Y(ori_ori_n523_));
  NO4        o0495(.A(n), .B(d), .C(ori_ori_n111_), .D(a), .Y(ori_ori_n524_));
  OR2        o0496(.A(n), .B(c), .Y(ori_ori_n525_));
  NO2        o0497(.A(ori_ori_n525_), .B(ori_ori_n144_), .Y(ori_ori_n526_));
  NO2        o0498(.A(ori_ori_n526_), .B(ori_ori_n524_), .Y(ori_ori_n527_));
  NOi32      o0499(.An(g), .Bn(f), .C(i), .Y(ori_ori_n528_));
  AOI220     o0500(.A0(ori_ori_n528_), .A1(ori_ori_n96_), .B0(ori_ori_n511_), .B1(f), .Y(ori_ori_n529_));
  NO2        o0501(.A(ori_ori_n271_), .B(ori_ori_n49_), .Y(ori_ori_n530_));
  NO2        o0502(.A(ori_ori_n529_), .B(ori_ori_n527_), .Y(ori_ori_n531_));
  INV        o0503(.A(ori_ori_n531_), .Y(ori_ori_n532_));
  NA2        o0504(.A(ori_ori_n134_), .B(ori_ori_n34_), .Y(ori_ori_n533_));
  OAI220     o0505(.A0(ori_ori_n533_), .A1(m), .B0(ori_ori_n514_), .B1(ori_ori_n229_), .Y(ori_ori_n534_));
  NOi41      o0506(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n535_));
  NAi32      o0507(.An(e), .Bn(b), .C(c), .Y(ori_ori_n536_));
  OR2        o0508(.A(ori_ori_n536_), .B(ori_ori_n80_), .Y(ori_ori_n537_));
  AN2        o0509(.A(ori_ori_n330_), .B(ori_ori_n312_), .Y(ori_ori_n538_));
  NA2        o0510(.A(ori_ori_n538_), .B(ori_ori_n537_), .Y(ori_ori_n539_));
  OA210      o0511(.A0(ori_ori_n539_), .A1(ori_ori_n535_), .B0(ori_ori_n534_), .Y(ori_ori_n540_));
  OAI220     o0512(.A0(ori_ori_n390_), .A1(ori_ori_n389_), .B0(ori_ori_n509_), .B1(ori_ori_n508_), .Y(ori_ori_n541_));
  NO2        o0513(.A(ori_ori_n226_), .B(ori_ori_n106_), .Y(ori_ori_n542_));
  NA2        o0514(.A(ori_ori_n391_), .B(ori_ori_n542_), .Y(ori_ori_n543_));
  INV        o0515(.A(ori_ori_n543_), .Y(ori_ori_n544_));
  NO2        o0516(.A(ori_ori_n273_), .B(n), .Y(ori_ori_n545_));
  NO2        o0517(.A(ori_ori_n417_), .B(ori_ori_n545_), .Y(ori_ori_n546_));
  NA2        o0518(.A(ori_ori_n541_), .B(f), .Y(ori_ori_n547_));
  NAi32      o0519(.An(d), .Bn(a), .C(b), .Y(ori_ori_n548_));
  NO2        o0520(.A(ori_ori_n548_), .B(ori_ori_n49_), .Y(ori_ori_n549_));
  NA2        o0521(.A(h), .B(f), .Y(ori_ori_n550_));
  NO2        o0522(.A(ori_ori_n550_), .B(ori_ori_n91_), .Y(ori_ori_n551_));
  NO3        o0523(.A(ori_ori_n171_), .B(ori_ori_n168_), .C(g), .Y(ori_ori_n552_));
  AOI220     o0524(.A0(ori_ori_n552_), .A1(ori_ori_n58_), .B0(ori_ori_n551_), .B1(ori_ori_n549_), .Y(ori_ori_n553_));
  OAI210     o0525(.A0(ori_ori_n547_), .A1(ori_ori_n546_), .B0(ori_ori_n553_), .Y(ori_ori_n554_));
  AN3        o0526(.A(j), .B(h), .C(g), .Y(ori_ori_n555_));
  NO2        o0527(.A(ori_ori_n141_), .B(c), .Y(ori_ori_n556_));
  NA3        o0528(.A(ori_ori_n556_), .B(ori_ori_n555_), .C(ori_ori_n441_), .Y(ori_ori_n557_));
  NA3        o0529(.A(f), .B(d), .C(b), .Y(ori_ori_n558_));
  NO4        o0530(.A(ori_ori_n558_), .B(ori_ori_n171_), .C(ori_ori_n168_), .D(g), .Y(ori_ori_n559_));
  NAi21      o0531(.An(ori_ori_n559_), .B(ori_ori_n557_), .Y(ori_ori_n560_));
  NO4        o0532(.A(ori_ori_n560_), .B(ori_ori_n554_), .C(ori_ori_n544_), .D(ori_ori_n540_), .Y(ori_ori_n561_));
  AN4        o0533(.A(ori_ori_n561_), .B(ori_ori_n532_), .C(ori_ori_n518_), .D(ori_ori_n512_), .Y(ori_ori_n562_));
  INV        o0534(.A(k), .Y(ori_ori_n563_));
  NA3        o0535(.A(l), .B(ori_ori_n563_), .C(i), .Y(ori_ori_n564_));
  INV        o0536(.A(ori_ori_n564_), .Y(ori_ori_n565_));
  NAi32      o0537(.An(h), .Bn(f), .C(g), .Y(ori_ori_n566_));
  NAi41      o0538(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n567_));
  OAI210     o0539(.A0(ori_ori_n516_), .A1(n), .B0(ori_ori_n567_), .Y(ori_ori_n568_));
  NA2        o0540(.A(ori_ori_n568_), .B(m), .Y(ori_ori_n569_));
  NAi31      o0541(.An(h), .B(g), .C(f), .Y(ori_ori_n570_));
  NO3        o0542(.A(ori_ori_n566_), .B(ori_ori_n68_), .C(ori_ori_n69_), .Y(ori_ori_n571_));
  NO4        o0543(.A(ori_ori_n570_), .B(ori_ori_n525_), .C(ori_ori_n144_), .D(ori_ori_n69_), .Y(ori_ori_n572_));
  OR2        o0544(.A(ori_ori_n572_), .B(ori_ori_n571_), .Y(ori_ori_n573_));
  NAi31      o0545(.An(f), .B(h), .C(g), .Y(ori_ori_n574_));
  NOi32      o0546(.An(b), .Bn(a), .C(c), .Y(ori_ori_n575_));
  NOi32      o0547(.An(d), .Bn(a), .C(e), .Y(ori_ori_n576_));
  NA2        o0548(.A(ori_ori_n576_), .B(ori_ori_n109_), .Y(ori_ori_n577_));
  NO2        o0549(.A(n), .B(c), .Y(ori_ori_n578_));
  NA3        o0550(.A(ori_ori_n578_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n579_));
  NA2        o0551(.A(ori_ori_n579_), .B(ori_ori_n577_), .Y(ori_ori_n580_));
  NOi32      o0552(.An(e), .Bn(a), .C(d), .Y(ori_ori_n581_));
  AOI210     o0553(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n581_), .Y(ori_ori_n582_));
  INV        o0554(.A(ori_ori_n533_), .Y(ori_ori_n583_));
  NA2        o0555(.A(ori_ori_n583_), .B(ori_ori_n580_), .Y(ori_ori_n584_));
  OAI210     o0556(.A0(ori_ori_n244_), .A1(ori_ori_n83_), .B0(ori_ori_n584_), .Y(ori_ori_n585_));
  AOI210     o0557(.A0(ori_ori_n573_), .A1(ori_ori_n565_), .B0(ori_ori_n585_), .Y(ori_ori_n586_));
  NO3        o0558(.A(ori_ori_n310_), .B(ori_ori_n60_), .C(n), .Y(ori_ori_n587_));
  NA3        o0559(.A(ori_ori_n494_), .B(ori_ori_n166_), .C(ori_ori_n165_), .Y(ori_ori_n588_));
  NA2        o0560(.A(ori_ori_n443_), .B(ori_ori_n226_), .Y(ori_ori_n589_));
  OR2        o0561(.A(ori_ori_n589_), .B(ori_ori_n588_), .Y(ori_ori_n590_));
  NA2        o0562(.A(ori_ori_n590_), .B(ori_ori_n587_), .Y(ori_ori_n591_));
  NO2        o0563(.A(ori_ori_n591_), .B(ori_ori_n83_), .Y(ori_ori_n592_));
  NA3        o0564(.A(ori_ori_n535_), .B(ori_ori_n332_), .C(ori_ori_n46_), .Y(ori_ori_n593_));
  NOi32      o0565(.An(e), .Bn(c), .C(f), .Y(ori_ori_n594_));
  NOi21      o0566(.An(f), .B(g), .Y(ori_ori_n595_));
  NO2        o0567(.A(ori_ori_n595_), .B(ori_ori_n206_), .Y(ori_ori_n596_));
  AOI220     o0568(.A0(ori_ori_n596_), .A1(ori_ori_n384_), .B0(ori_ori_n594_), .B1(ori_ori_n170_), .Y(ori_ori_n597_));
  NA3        o0569(.A(ori_ori_n597_), .B(ori_ori_n593_), .C(ori_ori_n173_), .Y(ori_ori_n598_));
  AOI210     o0570(.A0(ori_ori_n520_), .A1(ori_ori_n388_), .B0(ori_ori_n293_), .Y(ori_ori_n599_));
  NA2        o0571(.A(ori_ori_n599_), .B(ori_ori_n261_), .Y(ori_ori_n600_));
  NOi21      o0572(.An(j), .B(l), .Y(ori_ori_n601_));
  NAi21      o0573(.An(k), .B(h), .Y(ori_ori_n602_));
  NO2        o0574(.A(ori_ori_n602_), .B(ori_ori_n259_), .Y(ori_ori_n603_));
  NA2        o0575(.A(ori_ori_n603_), .B(ori_ori_n601_), .Y(ori_ori_n604_));
  OR2        o0576(.A(ori_ori_n604_), .B(ori_ori_n569_), .Y(ori_ori_n605_));
  NOi31      o0577(.An(m), .B(n), .C(k), .Y(ori_ori_n606_));
  NA2        o0578(.A(ori_ori_n601_), .B(ori_ori_n606_), .Y(ori_ori_n607_));
  AOI210     o0579(.A0(ori_ori_n388_), .A1(ori_ori_n364_), .B0(ori_ori_n293_), .Y(ori_ori_n608_));
  NAi21      o0580(.An(ori_ori_n607_), .B(ori_ori_n608_), .Y(ori_ori_n609_));
  NO2        o0581(.A(ori_ori_n273_), .B(ori_ori_n49_), .Y(ori_ori_n610_));
  NO2        o0582(.A(ori_ori_n304_), .B(ori_ori_n574_), .Y(ori_ori_n611_));
  NO2        o0583(.A(ori_ori_n516_), .B(ori_ori_n49_), .Y(ori_ori_n612_));
  AOI220     o0584(.A0(ori_ori_n612_), .A1(ori_ori_n611_), .B0(ori_ori_n610_), .B1(ori_ori_n551_), .Y(ori_ori_n613_));
  NA4        o0585(.A(ori_ori_n613_), .B(ori_ori_n609_), .C(ori_ori_n605_), .D(ori_ori_n600_), .Y(ori_ori_n614_));
  NA2        o0586(.A(ori_ori_n105_), .B(ori_ori_n36_), .Y(ori_ori_n615_));
  NO2        o0587(.A(k), .B(ori_ori_n209_), .Y(ori_ori_n616_));
  INV        o0588(.A(ori_ori_n353_), .Y(ori_ori_n617_));
  NO2        o0589(.A(ori_ori_n617_), .B(n), .Y(ori_ori_n618_));
  NAi31      o0590(.An(ori_ori_n615_), .B(ori_ori_n618_), .C(ori_ori_n616_), .Y(ori_ori_n619_));
  NO2        o0591(.A(ori_ori_n514_), .B(ori_ori_n171_), .Y(ori_ori_n620_));
  NA3        o0592(.A(ori_ori_n536_), .B(ori_ori_n267_), .C(ori_ori_n139_), .Y(ori_ori_n621_));
  NA2        o0593(.A(ori_ori_n490_), .B(ori_ori_n155_), .Y(ori_ori_n622_));
  NO3        o0594(.A(ori_ori_n385_), .B(ori_ori_n622_), .C(ori_ori_n83_), .Y(ori_ori_n623_));
  AOI210     o0595(.A0(ori_ori_n621_), .A1(ori_ori_n620_), .B0(ori_ori_n623_), .Y(ori_ori_n624_));
  AN3        o0596(.A(f), .B(d), .C(b), .Y(ori_ori_n625_));
  OAI210     o0597(.A0(ori_ori_n625_), .A1(ori_ori_n125_), .B0(n), .Y(ori_ori_n626_));
  NA3        o0598(.A(ori_ori_n490_), .B(ori_ori_n155_), .C(ori_ori_n209_), .Y(ori_ori_n627_));
  AOI210     o0599(.A0(ori_ori_n626_), .A1(ori_ori_n228_), .B0(ori_ori_n627_), .Y(ori_ori_n628_));
  NAi31      o0600(.An(m), .B(n), .C(k), .Y(ori_ori_n629_));
  OR2        o0601(.A(ori_ori_n128_), .B(ori_ori_n60_), .Y(ori_ori_n630_));
  OAI210     o0602(.A0(ori_ori_n630_), .A1(ori_ori_n629_), .B0(ori_ori_n246_), .Y(ori_ori_n631_));
  OAI210     o0603(.A0(ori_ori_n631_), .A1(ori_ori_n628_), .B0(j), .Y(ori_ori_n632_));
  NA3        o0604(.A(ori_ori_n632_), .B(ori_ori_n624_), .C(ori_ori_n619_), .Y(ori_ori_n633_));
  NO4        o0605(.A(ori_ori_n633_), .B(ori_ori_n614_), .C(ori_ori_n598_), .D(ori_ori_n592_), .Y(ori_ori_n634_));
  NAi31      o0606(.An(g), .B(h), .C(f), .Y(ori_ori_n635_));
  OR3        o0607(.A(ori_ori_n635_), .B(ori_ori_n273_), .C(n), .Y(ori_ori_n636_));
  OA210      o0608(.A0(ori_ori_n516_), .A1(n), .B0(ori_ori_n567_), .Y(ori_ori_n637_));
  NA3        o0609(.A(ori_ori_n406_), .B(ori_ori_n116_), .C(ori_ori_n80_), .Y(ori_ori_n638_));
  OAI210     o0610(.A0(ori_ori_n637_), .A1(ori_ori_n87_), .B0(ori_ori_n638_), .Y(ori_ori_n639_));
  NOi21      o0611(.An(ori_ori_n636_), .B(ori_ori_n639_), .Y(ori_ori_n640_));
  NO2        o0612(.A(ori_ori_n640_), .B(ori_ori_n510_), .Y(ori_ori_n641_));
  NO3        o0613(.A(g), .B(ori_ori_n208_), .C(ori_ori_n56_), .Y(ori_ori_n642_));
  NAi21      o0614(.An(h), .B(j), .Y(ori_ori_n643_));
  NA2        o0615(.A(ori_ori_n384_), .B(ori_ori_n642_), .Y(ori_ori_n644_));
  OR2        o0616(.A(ori_ori_n68_), .B(ori_ori_n69_), .Y(ori_ori_n645_));
  NA2        o0617(.A(ori_ori_n575_), .B(ori_ori_n334_), .Y(ori_ori_n646_));
  OA220      o0618(.A0(ori_ori_n607_), .A1(ori_ori_n646_), .B0(ori_ori_n604_), .B1(ori_ori_n645_), .Y(ori_ori_n647_));
  NA3        o0619(.A(ori_ori_n507_), .B(ori_ori_n96_), .C(ori_ori_n95_), .Y(ori_ori_n648_));
  AN2        o0620(.A(h), .B(f), .Y(ori_ori_n649_));
  NA2        o0621(.A(ori_ori_n649_), .B(ori_ori_n37_), .Y(ori_ori_n650_));
  NA2        o0622(.A(ori_ori_n96_), .B(ori_ori_n46_), .Y(ori_ori_n651_));
  OAI220     o0623(.A0(ori_ori_n651_), .A1(ori_ori_n323_), .B0(ori_ori_n650_), .B1(ori_ori_n448_), .Y(ori_ori_n652_));
  AOI210     o0624(.A0(ori_ori_n548_), .A1(ori_ori_n416_), .B0(ori_ori_n49_), .Y(ori_ori_n653_));
  INV        o0625(.A(ori_ori_n652_), .Y(ori_ori_n654_));
  NA4        o0626(.A(ori_ori_n654_), .B(ori_ori_n648_), .C(ori_ori_n647_), .D(ori_ori_n644_), .Y(ori_ori_n655_));
  NA2        o0627(.A(ori_ori_n127_), .B(ori_ori_n49_), .Y(ori_ori_n656_));
  AOI220     o0628(.A0(ori_ori_n656_), .A1(ori_ori_n513_), .B0(ori_ori_n353_), .B1(ori_ori_n109_), .Y(ori_ori_n657_));
  OA220      o0629(.A0(ori_ori_n657_), .A1(ori_ori_n533_), .B0(ori_ori_n351_), .B1(ori_ori_n107_), .Y(ori_ori_n658_));
  INV        o0630(.A(ori_ori_n658_), .Y(ori_ori_n659_));
  NO3        o0631(.A(ori_ori_n395_), .B(ori_ori_n187_), .C(ori_ori_n186_), .Y(ori_ori_n660_));
  NA2        o0632(.A(ori_ori_n660_), .B(ori_ori_n226_), .Y(ori_ori_n661_));
  NA3        o0633(.A(ori_ori_n661_), .B(ori_ori_n250_), .C(j), .Y(ori_ori_n662_));
  NO3        o0634(.A(ori_ori_n443_), .B(ori_ori_n168_), .C(i), .Y(ori_ori_n663_));
  NA2        o0635(.A(ori_ori_n447_), .B(ori_ori_n80_), .Y(ori_ori_n664_));
  NA2        o0636(.A(ori_ori_n662_), .B(ori_ori_n393_), .Y(ori_ori_n665_));
  NO4        o0637(.A(ori_ori_n665_), .B(ori_ori_n659_), .C(ori_ori_n655_), .D(ori_ori_n641_), .Y(ori_ori_n666_));
  NA4        o0638(.A(ori_ori_n666_), .B(ori_ori_n634_), .C(ori_ori_n586_), .D(ori_ori_n562_), .Y(ori08));
  NO2        o0639(.A(k), .B(h), .Y(ori_ori_n668_));
  AO210      o0640(.A0(ori_ori_n248_), .A1(ori_ori_n433_), .B0(ori_ori_n668_), .Y(ori_ori_n669_));
  NO2        o0641(.A(ori_ori_n669_), .B(ori_ori_n291_), .Y(ori_ori_n670_));
  NA2        o0642(.A(ori_ori_n594_), .B(ori_ori_n80_), .Y(ori_ori_n671_));
  NA2        o0643(.A(ori_ori_n671_), .B(ori_ori_n443_), .Y(ori_ori_n672_));
  AOI210     o0644(.A0(ori_ori_n672_), .A1(ori_ori_n670_), .B0(ori_ori_n475_), .Y(ori_ori_n673_));
  NA2        o0645(.A(ori_ori_n80_), .B(ori_ori_n106_), .Y(ori_ori_n674_));
  NO2        o0646(.A(ori_ori_n674_), .B(ori_ori_n57_), .Y(ori_ori_n675_));
  NO4        o0647(.A(ori_ori_n371_), .B(ori_ori_n108_), .C(j), .D(ori_ori_n209_), .Y(ori_ori_n676_));
  NA2        o0648(.A(ori_ori_n558_), .B(ori_ori_n228_), .Y(ori_ori_n677_));
  AOI220     o0649(.A0(ori_ori_n677_), .A1(ori_ori_n340_), .B0(ori_ori_n676_), .B1(ori_ori_n675_), .Y(ori_ori_n678_));
  AOI210     o0650(.A0(ori_ori_n558_), .A1(ori_ori_n151_), .B0(ori_ori_n80_), .Y(ori_ori_n679_));
  NA4        o0651(.A(ori_ori_n211_), .B(ori_ori_n134_), .C(ori_ori_n45_), .D(h), .Y(ori_ori_n680_));
  AN2        o0652(.A(l), .B(k), .Y(ori_ori_n681_));
  NA4        o0653(.A(ori_ori_n681_), .B(ori_ori_n105_), .C(ori_ori_n69_), .D(ori_ori_n209_), .Y(ori_ori_n682_));
  OAI210     o0654(.A0(ori_ori_n680_), .A1(g), .B0(ori_ori_n682_), .Y(ori_ori_n683_));
  NA2        o0655(.A(ori_ori_n683_), .B(ori_ori_n679_), .Y(ori_ori_n684_));
  NA4        o0656(.A(ori_ori_n684_), .B(ori_ori_n678_), .C(ori_ori_n673_), .D(ori_ori_n342_), .Y(ori_ori_n685_));
  AN2        o0657(.A(ori_ori_n517_), .B(ori_ori_n92_), .Y(ori_ori_n686_));
  NO4        o0658(.A(ori_ori_n168_), .B(ori_ori_n383_), .C(ori_ori_n108_), .D(g), .Y(ori_ori_n687_));
  AOI210     o0659(.A0(ori_ori_n687_), .A1(ori_ori_n677_), .B0(ori_ori_n502_), .Y(ori_ori_n688_));
  NO2        o0660(.A(ori_ori_n38_), .B(ori_ori_n208_), .Y(ori_ori_n689_));
  AOI220     o0661(.A0(ori_ori_n596_), .A1(ori_ori_n339_), .B0(ori_ori_n689_), .B1(ori_ori_n545_), .Y(ori_ori_n690_));
  NAi31      o0662(.An(ori_ori_n686_), .B(ori_ori_n690_), .C(ori_ori_n688_), .Y(ori_ori_n691_));
  OAI210     o0663(.A0(ori_ori_n536_), .A1(ori_ori_n47_), .B0(ori_ori_n630_), .Y(ori_ori_n692_));
  NO2        o0664(.A(ori_ori_n469_), .B(ori_ori_n127_), .Y(ori_ori_n693_));
  NA2        o0665(.A(ori_ori_n693_), .B(ori_ori_n692_), .Y(ori_ori_n694_));
  NO3        o0666(.A(ori_ori_n310_), .B(ori_ori_n126_), .C(ori_ori_n41_), .Y(ori_ori_n695_));
  NAi21      o0667(.An(ori_ori_n695_), .B(ori_ori_n682_), .Y(ori_ori_n696_));
  NA2        o0668(.A(ori_ori_n669_), .B(ori_ori_n129_), .Y(ori_ori_n697_));
  AOI220     o0669(.A0(ori_ori_n697_), .A1(ori_ori_n394_), .B0(ori_ori_n696_), .B1(ori_ori_n72_), .Y(ori_ori_n698_));
  NA2        o0670(.A(ori_ori_n694_), .B(ori_ori_n698_), .Y(ori_ori_n699_));
  NA2        o0671(.A(ori_ori_n353_), .B(ori_ori_n43_), .Y(ori_ori_n700_));
  NA3        o0672(.A(ori_ori_n661_), .B(ori_ori_n325_), .C(ori_ori_n375_), .Y(ori_ori_n701_));
  NA3        o0673(.A(m), .B(l), .C(k), .Y(ori_ori_n702_));
  AOI210     o0674(.A0(ori_ori_n638_), .A1(ori_ori_n636_), .B0(ori_ori_n702_), .Y(ori_ori_n703_));
  NA3        o0675(.A(ori_ori_n109_), .B(k), .C(ori_ori_n83_), .Y(ori_ori_n704_));
  INV        o0676(.A(ori_ori_n703_), .Y(ori_ori_n705_));
  NA3        o0677(.A(ori_ori_n705_), .B(ori_ori_n701_), .C(ori_ori_n700_), .Y(ori_ori_n706_));
  NO4        o0678(.A(ori_ori_n706_), .B(ori_ori_n699_), .C(ori_ori_n691_), .D(ori_ori_n685_), .Y(ori_ori_n707_));
  NA2        o0679(.A(ori_ori_n596_), .B(ori_ori_n384_), .Y(ori_ori_n708_));
  NA2        o0680(.A(ori_ori_n708_), .B(ori_ori_n247_), .Y(ori_ori_n709_));
  NA2        o0681(.A(ori_ori_n681_), .B(ori_ori_n69_), .Y(ori_ori_n710_));
  NO4        o0682(.A(ori_ori_n660_), .B(ori_ori_n168_), .C(n), .D(i), .Y(ori_ori_n711_));
  NOi21      o0683(.An(h), .B(j), .Y(ori_ori_n712_));
  NA2        o0684(.A(ori_ori_n712_), .B(f), .Y(ori_ori_n713_));
  NO2        o0685(.A(ori_ori_n713_), .B(ori_ori_n241_), .Y(ori_ori_n714_));
  NO3        o0686(.A(ori_ori_n714_), .B(ori_ori_n711_), .C(ori_ori_n663_), .Y(ori_ori_n715_));
  NO2        o0687(.A(ori_ori_n715_), .B(ori_ori_n710_), .Y(ori_ori_n716_));
  AOI210     o0688(.A0(ori_ori_n709_), .A1(l), .B0(ori_ori_n716_), .Y(ori_ori_n717_));
  NO2        o0689(.A(j), .B(i), .Y(ori_ori_n718_));
  NA3        o0690(.A(ori_ori_n718_), .B(ori_ori_n76_), .C(l), .Y(ori_ori_n719_));
  NA2        o0691(.A(ori_ori_n718_), .B(ori_ori_n33_), .Y(ori_ori_n720_));
  OR2        o0692(.A(ori_ori_n719_), .B(ori_ori_n569_), .Y(ori_ori_n721_));
  NO3        o0693(.A(ori_ori_n146_), .B(ori_ori_n49_), .C(ori_ori_n106_), .Y(ori_ori_n722_));
  NO3        o0694(.A(ori_ori_n525_), .B(ori_ori_n144_), .C(ori_ori_n69_), .Y(ori_ori_n723_));
  NO3        o0695(.A(ori_ori_n469_), .B(ori_ori_n425_), .C(j), .Y(ori_ori_n724_));
  AOI210     o0696(.A0(ori_ori_n513_), .A1(n), .B0(ori_ori_n535_), .Y(ori_ori_n725_));
  NA2        o0697(.A(ori_ori_n725_), .B(ori_ori_n538_), .Y(ori_ori_n726_));
  NO3        o0698(.A(ori_ori_n168_), .B(ori_ori_n383_), .C(ori_ori_n108_), .Y(ori_ori_n727_));
  AOI220     o0699(.A0(ori_ori_n727_), .A1(ori_ori_n242_), .B0(ori_ori_n589_), .B1(ori_ori_n302_), .Y(ori_ori_n728_));
  NAi31      o0700(.An(ori_ori_n582_), .B(ori_ori_n89_), .C(ori_ori_n80_), .Y(ori_ori_n729_));
  NA2        o0701(.A(ori_ori_n729_), .B(ori_ori_n728_), .Y(ori_ori_n730_));
  NO2        o0702(.A(ori_ori_n291_), .B(ori_ori_n129_), .Y(ori_ori_n731_));
  AOI220     o0703(.A0(ori_ori_n731_), .A1(ori_ori_n596_), .B0(ori_ori_n695_), .B1(ori_ori_n679_), .Y(ori_ori_n732_));
  NO2        o0704(.A(ori_ori_n702_), .B(ori_ori_n87_), .Y(ori_ori_n733_));
  NA2        o0705(.A(ori_ori_n724_), .B(ori_ori_n653_), .Y(ori_ori_n734_));
  NA2        o0706(.A(ori_ori_n734_), .B(ori_ori_n732_), .Y(ori_ori_n735_));
  OR2        o0707(.A(ori_ori_n735_), .B(ori_ori_n730_), .Y(ori_ori_n736_));
  NA3        o0708(.A(ori_ori_n725_), .B(ori_ori_n538_), .C(ori_ori_n537_), .Y(ori_ori_n737_));
  NA4        o0709(.A(ori_ori_n737_), .B(ori_ori_n211_), .C(ori_ori_n433_), .D(ori_ori_n34_), .Y(ori_ori_n738_));
  NO4        o0710(.A(ori_ori_n469_), .B(ori_ori_n421_), .C(j), .D(f), .Y(ori_ori_n739_));
  OAI220     o0711(.A0(ori_ori_n680_), .A1(ori_ori_n671_), .B0(ori_ori_n323_), .B1(ori_ori_n38_), .Y(ori_ori_n740_));
  AOI210     o0712(.A0(ori_ori_n739_), .A1(ori_ori_n254_), .B0(ori_ori_n740_), .Y(ori_ori_n741_));
  NA3        o0713(.A(ori_ori_n528_), .B(ori_ori_n288_), .C(h), .Y(ori_ori_n742_));
  NO2        o0714(.A(ori_ori_n88_), .B(ori_ori_n47_), .Y(ori_ori_n743_));
  OAI220     o0715(.A0(ori_ori_n742_), .A1(ori_ori_n579_), .B0(ori_ori_n719_), .B1(ori_ori_n645_), .Y(ori_ori_n744_));
  AOI210     o0716(.A0(ori_ori_n743_), .A1(ori_ori_n618_), .B0(ori_ori_n744_), .Y(ori_ori_n745_));
  NA3        o0717(.A(ori_ori_n745_), .B(ori_ori_n741_), .C(ori_ori_n738_), .Y(ori_ori_n746_));
  OR2        o0718(.A(ori_ori_n733_), .B(ori_ori_n92_), .Y(ori_ori_n747_));
  AOI220     o0719(.A0(ori_ori_n747_), .A1(ori_ori_n233_), .B0(ori_ori_n724_), .B1(ori_ori_n610_), .Y(ori_ori_n748_));
  NO2        o0720(.A(ori_ori_n637_), .B(ori_ori_n69_), .Y(ori_ori_n749_));
  AOI210     o0721(.A0(ori_ori_n739_), .A1(ori_ori_n749_), .B0(ori_ori_n327_), .Y(ori_ori_n750_));
  OAI210     o0722(.A0(ori_ori_n702_), .A1(ori_ori_n635_), .B0(ori_ori_n501_), .Y(ori_ori_n751_));
  NA3        o0723(.A(ori_ori_n245_), .B(ori_ori_n59_), .C(b), .Y(ori_ori_n752_));
  AOI220     o0724(.A0(ori_ori_n578_), .A1(ori_ori_n29_), .B0(ori_ori_n447_), .B1(ori_ori_n80_), .Y(ori_ori_n753_));
  NA2        o0725(.A(ori_ori_n753_), .B(ori_ori_n752_), .Y(ori_ori_n754_));
  NA2        o0726(.A(ori_ori_n754_), .B(ori_ori_n751_), .Y(ori_ori_n755_));
  NA3        o0727(.A(ori_ori_n755_), .B(ori_ori_n750_), .C(ori_ori_n748_), .Y(ori_ori_n756_));
  NOi41      o0728(.An(ori_ori_n721_), .B(ori_ori_n756_), .C(ori_ori_n746_), .D(ori_ori_n736_), .Y(ori_ori_n757_));
  NO3        o0729(.A(ori_ori_n333_), .B(ori_ori_n293_), .C(ori_ori_n108_), .Y(ori_ori_n758_));
  NA2        o0730(.A(ori_ori_n758_), .B(ori_ori_n726_), .Y(ori_ori_n759_));
  NO3        o0731(.A(ori_ori_n508_), .B(ori_ori_n90_), .C(h), .Y(ori_ori_n760_));
  NA2        o0732(.A(ori_ori_n760_), .B(ori_ori_n675_), .Y(ori_ori_n761_));
  NA3        o0733(.A(ori_ori_n761_), .B(ori_ori_n759_), .C(ori_ori_n396_), .Y(ori_ori_n762_));
  OR2        o0734(.A(ori_ori_n635_), .B(ori_ori_n88_), .Y(ori_ori_n763_));
  NOi31      o0735(.An(b), .B(d), .C(a), .Y(ori_ori_n764_));
  NO2        o0736(.A(ori_ori_n764_), .B(ori_ori_n576_), .Y(ori_ori_n765_));
  NO2        o0737(.A(ori_ori_n765_), .B(n), .Y(ori_ori_n766_));
  NOi21      o0738(.An(ori_ori_n753_), .B(ori_ori_n766_), .Y(ori_ori_n767_));
  OAI220     o0739(.A0(ori_ori_n767_), .A1(ori_ori_n763_), .B0(ori_ori_n742_), .B1(ori_ori_n577_), .Y(ori_ori_n768_));
  NO2        o0740(.A(ori_ori_n536_), .B(ori_ori_n80_), .Y(ori_ori_n769_));
  NO3        o0741(.A(ori_ori_n595_), .B(ori_ori_n320_), .C(ori_ori_n112_), .Y(ori_ori_n770_));
  NOi21      o0742(.An(ori_ori_n770_), .B(ori_ori_n156_), .Y(ori_ori_n771_));
  AOI210     o0743(.A0(ori_ori_n758_), .A1(ori_ori_n769_), .B0(ori_ori_n771_), .Y(ori_ori_n772_));
  OAI210     o0744(.A0(ori_ori_n680_), .A1(ori_ori_n385_), .B0(ori_ori_n772_), .Y(ori_ori_n773_));
  NO2        o0745(.A(ori_ori_n660_), .B(n), .Y(ori_ori_n774_));
  AOI220     o0746(.A0(ori_ori_n731_), .A1(ori_ori_n642_), .B0(ori_ori_n774_), .B1(ori_ori_n670_), .Y(ori_ori_n775_));
  NO2        o0747(.A(ori_ori_n317_), .B(ori_ori_n232_), .Y(ori_ori_n776_));
  OAI210     o0748(.A0(ori_ori_n92_), .A1(ori_ori_n89_), .B0(ori_ori_n776_), .Y(ori_ori_n777_));
  INV        o0749(.A(ori_ori_n777_), .Y(ori_ori_n778_));
  OAI210     o0750(.A0(ori_ori_n572_), .A1(ori_ori_n571_), .B0(ori_ori_n354_), .Y(ori_ori_n779_));
  NAi31      o0751(.An(ori_ori_n778_), .B(ori_ori_n779_), .C(ori_ori_n775_), .Y(ori_ori_n780_));
  NO4        o0752(.A(ori_ori_n780_), .B(ori_ori_n773_), .C(ori_ori_n768_), .D(ori_ori_n762_), .Y(ori_ori_n781_));
  NA4        o0753(.A(ori_ori_n781_), .B(ori_ori_n757_), .C(ori_ori_n717_), .D(ori_ori_n707_), .Y(ori09));
  INV        o0754(.A(ori_ori_n117_), .Y(ori_ori_n783_));
  NA2        o0755(.A(f), .B(e), .Y(ori_ori_n784_));
  NO2        o0756(.A(ori_ori_n221_), .B(ori_ori_n108_), .Y(ori_ori_n785_));
  NA4        o0757(.A(ori_ori_n304_), .B(ori_ori_n455_), .C(ori_ori_n257_), .D(ori_ori_n114_), .Y(ori_ori_n786_));
  AOI210     o0758(.A0(ori_ori_n786_), .A1(g), .B0(ori_ori_n452_), .Y(ori_ori_n787_));
  NO2        o0759(.A(ori_ori_n787_), .B(ori_ori_n784_), .Y(ori_ori_n788_));
  NA2        o0760(.A(ori_ori_n427_), .B(e), .Y(ori_ori_n789_));
  NO2        o0761(.A(ori_ori_n789_), .B(ori_ori_n494_), .Y(ori_ori_n790_));
  AOI210     o0762(.A0(ori_ori_n788_), .A1(ori_ori_n783_), .B0(ori_ori_n790_), .Y(ori_ori_n791_));
  NO2        o0763(.A(ori_ori_n199_), .B(ori_ori_n208_), .Y(ori_ori_n792_));
  NA3        o0764(.A(m), .B(l), .C(i), .Y(ori_ori_n793_));
  OAI220     o0765(.A0(ori_ori_n570_), .A1(ori_ori_n793_), .B0(ori_ori_n346_), .B1(ori_ori_n509_), .Y(ori_ori_n794_));
  NA4        o0766(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(g), .D(f), .Y(ori_ori_n795_));
  NAi21      o0767(.An(ori_ori_n794_), .B(ori_ori_n795_), .Y(ori_ori_n796_));
  OR2        o0768(.A(ori_ori_n796_), .B(ori_ori_n792_), .Y(ori_ori_n797_));
  NA3        o0769(.A(ori_ori_n763_), .B(ori_ori_n547_), .C(ori_ori_n501_), .Y(ori_ori_n798_));
  OA210      o0770(.A0(ori_ori_n798_), .A1(ori_ori_n797_), .B0(ori_ori_n766_), .Y(ori_ori_n799_));
  INV        o0771(.A(ori_ori_n330_), .Y(ori_ori_n800_));
  NO2        o0772(.A(ori_ori_n122_), .B(ori_ori_n120_), .Y(ori_ori_n801_));
  INV        o0773(.A(ori_ori_n332_), .Y(ori_ori_n802_));
  AOI210     o0774(.A0(ori_ori_n802_), .A1(ori_ori_n801_), .B0(ori_ori_n574_), .Y(ori_ori_n803_));
  NA2        o0775(.A(ori_ori_n752_), .B(ori_ori_n323_), .Y(ori_ori_n804_));
  NA2        o0776(.A(ori_ori_n334_), .B(ori_ori_n336_), .Y(ori_ori_n805_));
  OAI210     o0777(.A0(ori_ori_n199_), .A1(ori_ori_n208_), .B0(ori_ori_n805_), .Y(ori_ori_n806_));
  AOI220     o0778(.A0(ori_ori_n806_), .A1(ori_ori_n804_), .B0(ori_ori_n803_), .B1(ori_ori_n800_), .Y(ori_ori_n807_));
  NA2        o0779(.A(ori_ori_n669_), .B(ori_ori_n129_), .Y(ori_ori_n808_));
  NA3        o0780(.A(ori_ori_n808_), .B(ori_ori_n184_), .C(ori_ori_n31_), .Y(ori_ori_n809_));
  NA4        o0781(.A(ori_ori_n809_), .B(ori_ori_n807_), .C(ori_ori_n597_), .D(ori_ori_n78_), .Y(ori_ori_n810_));
  NO2        o0782(.A(ori_ori_n566_), .B(ori_ori_n481_), .Y(ori_ori_n811_));
  NA2        o0783(.A(ori_ori_n811_), .B(ori_ori_n184_), .Y(ori_ori_n812_));
  NOi21      o0784(.An(f), .B(d), .Y(ori_ori_n813_));
  NA2        o0785(.A(ori_ori_n813_), .B(m), .Y(ori_ori_n814_));
  NO2        o0786(.A(ori_ori_n814_), .B(ori_ori_n52_), .Y(ori_ori_n815_));
  NOi32      o0787(.An(g), .Bn(f), .C(d), .Y(ori_ori_n816_));
  NA4        o0788(.A(ori_ori_n816_), .B(ori_ori_n578_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n817_));
  NOi21      o0789(.An(ori_ori_n305_), .B(ori_ori_n817_), .Y(ori_ori_n818_));
  AOI210     o0790(.A0(ori_ori_n815_), .A1(ori_ori_n526_), .B0(ori_ori_n818_), .Y(ori_ori_n819_));
  NA2        o0791(.A(ori_ori_n304_), .B(ori_ori_n257_), .Y(ori_ori_n820_));
  AN2        o0792(.A(f), .B(d), .Y(ori_ori_n821_));
  NA3        o0793(.A(ori_ori_n460_), .B(ori_ori_n821_), .C(ori_ori_n80_), .Y(ori_ori_n822_));
  NO3        o0794(.A(ori_ori_n822_), .B(ori_ori_n69_), .C(ori_ori_n209_), .Y(ori_ori_n823_));
  NA2        o0795(.A(ori_ori_n820_), .B(ori_ori_n823_), .Y(ori_ori_n824_));
  NAi41      o0796(.An(ori_ori_n474_), .B(ori_ori_n824_), .C(ori_ori_n819_), .D(ori_ori_n812_), .Y(ori_ori_n825_));
  NO2        o0797(.A(ori_ori_n629_), .B(ori_ori_n320_), .Y(ori_ori_n826_));
  NA2        o0798(.A(ori_ori_n576_), .B(ori_ori_n80_), .Y(ori_ori_n827_));
  NO2        o0799(.A(ori_ori_n805_), .B(ori_ori_n827_), .Y(ori_ori_n828_));
  NOi31      o0800(.An(ori_ori_n219_), .B(ori_ori_n828_), .C(ori_ori_n300_), .Y(ori_ori_n829_));
  NA2        o0801(.A(c), .B(ori_ori_n111_), .Y(ori_ori_n830_));
  NO2        o0802(.A(ori_ori_n830_), .B(ori_ori_n400_), .Y(ori_ori_n831_));
  NA3        o0803(.A(ori_ori_n831_), .B(ori_ori_n492_), .C(f), .Y(ori_ori_n832_));
  OR2        o0804(.A(ori_ori_n635_), .B(ori_ori_n522_), .Y(ori_ori_n833_));
  INV        o0805(.A(ori_ori_n833_), .Y(ori_ori_n834_));
  NA2        o0806(.A(ori_ori_n765_), .B(ori_ori_n107_), .Y(ori_ori_n835_));
  NA2        o0807(.A(ori_ori_n835_), .B(ori_ori_n834_), .Y(ori_ori_n836_));
  NA3        o0808(.A(ori_ori_n836_), .B(ori_ori_n832_), .C(ori_ori_n829_), .Y(ori_ori_n837_));
  NO4        o0809(.A(ori_ori_n837_), .B(ori_ori_n825_), .C(ori_ori_n810_), .D(ori_ori_n799_), .Y(ori_ori_n838_));
  NA2        o0810(.A(ori_ori_n108_), .B(j), .Y(ori_ori_n839_));
  NO2        o0811(.A(ori_ori_n323_), .B(ori_ori_n795_), .Y(ori_ori_n840_));
  NO2        o0812(.A(ori_ori_n129_), .B(ori_ori_n127_), .Y(ori_ori_n841_));
  NO2        o0813(.A(ori_ori_n226_), .B(ori_ori_n220_), .Y(ori_ori_n842_));
  AOI220     o0814(.A0(ori_ori_n842_), .A1(ori_ori_n223_), .B0(ori_ori_n298_), .B1(ori_ori_n841_), .Y(ori_ori_n843_));
  INV        o0815(.A(ori_ori_n843_), .Y(ori_ori_n844_));
  NA2        o0816(.A(e), .B(d), .Y(ori_ori_n845_));
  OAI220     o0817(.A0(ori_ori_n845_), .A1(c), .B0(ori_ori_n317_), .B1(d), .Y(ori_ori_n846_));
  NA3        o0818(.A(ori_ori_n846_), .B(ori_ori_n436_), .C(ori_ori_n490_), .Y(ori_ori_n847_));
  AOI210     o0819(.A0(ori_ori_n497_), .A1(ori_ori_n175_), .B0(ori_ori_n226_), .Y(ori_ori_n848_));
  AOI210     o0820(.A0(ori_ori_n596_), .A1(ori_ori_n339_), .B0(ori_ori_n848_), .Y(ori_ori_n849_));
  NA2        o0821(.A(ori_ori_n281_), .B(ori_ori_n160_), .Y(ori_ori_n850_));
  NA2        o0822(.A(ori_ori_n823_), .B(ori_ori_n850_), .Y(ori_ori_n851_));
  NA3        o0823(.A(ori_ori_n851_), .B(ori_ori_n849_), .C(ori_ori_n847_), .Y(ori_ori_n852_));
  NO3        o0824(.A(ori_ori_n852_), .B(ori_ori_n844_), .C(ori_ori_n840_), .Y(ori_ori_n853_));
  NA2        o0825(.A(ori_ori_n800_), .B(ori_ori_n31_), .Y(ori_ori_n854_));
  AO210      o0826(.A0(ori_ori_n854_), .A1(ori_ori_n671_), .B0(ori_ori_n212_), .Y(ori_ori_n855_));
  OAI220     o0827(.A0(ori_ori_n595_), .A1(ori_ori_n60_), .B0(ori_ori_n293_), .B1(j), .Y(ori_ori_n856_));
  AOI220     o0828(.A0(ori_ori_n856_), .A1(ori_ori_n826_), .B0(ori_ori_n587_), .B1(ori_ori_n594_), .Y(ori_ori_n857_));
  OAI210     o0829(.A0(ori_ori_n789_), .A1(ori_ori_n165_), .B0(ori_ori_n857_), .Y(ori_ori_n858_));
  OAI210     o0830(.A0(ori_ori_n785_), .A1(ori_ori_n850_), .B0(ori_ori_n816_), .Y(ori_ori_n859_));
  NO2        o0831(.A(ori_ori_n859_), .B(ori_ori_n579_), .Y(ori_ori_n860_));
  AN2        o0832(.A(ori_ori_n804_), .B(ori_ori_n794_), .Y(ori_ori_n861_));
  NOi31      o0833(.An(ori_ori_n526_), .B(ori_ori_n814_), .C(ori_ori_n289_), .Y(ori_ori_n862_));
  NO4        o0834(.A(ori_ori_n862_), .B(ori_ori_n861_), .C(ori_ori_n860_), .D(ori_ori_n858_), .Y(ori_ori_n863_));
  AO220      o0835(.A0(ori_ori_n436_), .A1(ori_ori_n712_), .B0(ori_ori_n170_), .B1(f), .Y(ori_ori_n864_));
  OAI210     o0836(.A0(ori_ori_n864_), .A1(ori_ori_n439_), .B0(ori_ori_n846_), .Y(ori_ori_n865_));
  NO2        o0837(.A(ori_ori_n425_), .B(ori_ori_n66_), .Y(ori_ori_n866_));
  OAI210     o0838(.A0(ori_ori_n798_), .A1(ori_ori_n866_), .B0(ori_ori_n675_), .Y(ori_ori_n867_));
  AN4        o0839(.A(ori_ori_n867_), .B(ori_ori_n865_), .C(ori_ori_n863_), .D(ori_ori_n855_), .Y(ori_ori_n868_));
  NA4        o0840(.A(ori_ori_n868_), .B(ori_ori_n853_), .C(ori_ori_n838_), .D(ori_ori_n791_), .Y(ori12));
  NO2        o0841(.A(ori_ori_n434_), .B(c), .Y(ori_ori_n870_));
  NO4        o0842(.A(ori_ori_n426_), .B(ori_ori_n248_), .C(ori_ori_n563_), .D(ori_ori_n209_), .Y(ori_ori_n871_));
  NA2        o0843(.A(ori_ori_n871_), .B(ori_ori_n870_), .Y(ori_ori_n872_));
  NA2        o0844(.A(ori_ori_n526_), .B(ori_ori_n866_), .Y(ori_ori_n873_));
  NO2        o0845(.A(ori_ori_n434_), .B(ori_ori_n111_), .Y(ori_ori_n874_));
  NO2        o0846(.A(ori_ori_n801_), .B(ori_ori_n346_), .Y(ori_ori_n875_));
  NO2        o0847(.A(ori_ori_n635_), .B(ori_ori_n371_), .Y(ori_ori_n876_));
  AOI220     o0848(.A0(ori_ori_n876_), .A1(ori_ori_n524_), .B0(ori_ori_n875_), .B1(ori_ori_n874_), .Y(ori_ori_n877_));
  NA3        o0849(.A(ori_ori_n877_), .B(ori_ori_n873_), .C(ori_ori_n872_), .Y(ori_ori_n878_));
  AOI210     o0850(.A0(ori_ori_n229_), .A1(ori_ori_n329_), .B0(ori_ori_n196_), .Y(ori_ori_n879_));
  OR2        o0851(.A(ori_ori_n879_), .B(ori_ori_n871_), .Y(ori_ori_n880_));
  AOI210     o0852(.A0(ori_ori_n326_), .A1(ori_ori_n381_), .B0(ori_ori_n209_), .Y(ori_ori_n881_));
  OAI210     o0853(.A0(ori_ori_n881_), .A1(ori_ori_n880_), .B0(ori_ori_n395_), .Y(ori_ori_n882_));
  NO2        o0854(.A(ori_ori_n615_), .B(ori_ori_n259_), .Y(ori_ori_n883_));
  NO2        o0855(.A(ori_ori_n570_), .B(ori_ori_n793_), .Y(ori_ori_n884_));
  AOI220     o0856(.A0(ori_ori_n884_), .A1(ori_ori_n545_), .B0(ori_ori_n776_), .B1(ori_ori_n883_), .Y(ori_ori_n885_));
  NA2        o0857(.A(ori_ori_n885_), .B(ori_ori_n882_), .Y(ori_ori_n886_));
  OR2        o0858(.A(ori_ori_n318_), .B(ori_ori_n874_), .Y(ori_ori_n887_));
  NA2        o0859(.A(ori_ori_n887_), .B(ori_ori_n347_), .Y(ori_ori_n888_));
  NA4        o0860(.A(ori_ori_n427_), .B(ori_ori_n423_), .C(ori_ori_n176_), .D(g), .Y(ori_ori_n889_));
  NA2        o0861(.A(ori_ori_n889_), .B(ori_ori_n888_), .Y(ori_ori_n890_));
  NO3        o0862(.A(ori_ori_n640_), .B(ori_ori_n88_), .C(ori_ori_n45_), .Y(ori_ori_n891_));
  NO4        o0863(.A(ori_ori_n891_), .B(ori_ori_n890_), .C(ori_ori_n886_), .D(ori_ori_n878_), .Y(ori_ori_n892_));
  NO2        o0864(.A(ori_ori_n361_), .B(ori_ori_n360_), .Y(ori_ori_n893_));
  INV        o0865(.A(ori_ori_n68_), .Y(ori_ori_n894_));
  NA2        o0866(.A(ori_ori_n536_), .B(ori_ori_n139_), .Y(ori_ori_n895_));
  NOi21      o0867(.An(ori_ori_n34_), .B(ori_ori_n629_), .Y(ori_ori_n896_));
  AOI220     o0868(.A0(ori_ori_n896_), .A1(ori_ori_n895_), .B0(ori_ori_n894_), .B1(ori_ori_n893_), .Y(ori_ori_n897_));
  OAI210     o0869(.A0(ori_ori_n246_), .A1(ori_ori_n45_), .B0(ori_ori_n897_), .Y(ori_ori_n898_));
  INV        o0870(.A(ori_ori_n314_), .Y(ori_ori_n899_));
  NO2        o0871(.A(ori_ori_n49_), .B(ori_ori_n45_), .Y(ori_ori_n900_));
  NO2        o0872(.A(ori_ori_n488_), .B(ori_ori_n293_), .Y(ori_ori_n901_));
  INV        o0873(.A(ori_ori_n901_), .Y(ori_ori_n902_));
  NO2        o0874(.A(ori_ori_n902_), .B(ori_ori_n139_), .Y(ori_ori_n903_));
  INV        o0875(.A(ori_ori_n358_), .Y(ori_ori_n904_));
  NO4        o0876(.A(ori_ori_n904_), .B(ori_ori_n903_), .C(ori_ori_n899_), .D(ori_ori_n898_), .Y(ori_ori_n905_));
  NA2        o0877(.A(ori_ori_n339_), .B(g), .Y(ori_ori_n906_));
  NA2        o0878(.A(ori_ori_n158_), .B(i), .Y(ori_ori_n907_));
  NA2        o0879(.A(ori_ori_n46_), .B(i), .Y(ori_ori_n908_));
  OAI220     o0880(.A0(ori_ori_n908_), .A1(ori_ori_n195_), .B0(ori_ori_n907_), .B1(ori_ori_n88_), .Y(ori_ori_n909_));
  INV        o0881(.A(ori_ori_n909_), .Y(ori_ori_n910_));
  NA2        o0882(.A(ori_ori_n536_), .B(ori_ori_n373_), .Y(ori_ori_n911_));
  AOI210     o0883(.A0(ori_ori_n911_), .A1(n), .B0(ori_ori_n535_), .Y(ori_ori_n912_));
  OAI220     o0884(.A0(ori_ori_n912_), .A1(ori_ori_n906_), .B0(ori_ori_n910_), .B1(ori_ori_n323_), .Y(ori_ori_n913_));
  NO2        o0885(.A(ori_ori_n635_), .B(ori_ori_n481_), .Y(ori_ori_n914_));
  NA3        o0886(.A(ori_ori_n334_), .B(ori_ori_n601_), .C(i), .Y(ori_ori_n915_));
  OAI210     o0887(.A0(ori_ori_n425_), .A1(ori_ori_n304_), .B0(ori_ori_n915_), .Y(ori_ori_n916_));
  OAI220     o0888(.A0(ori_ori_n916_), .A1(ori_ori_n914_), .B0(ori_ori_n653_), .B1(ori_ori_n723_), .Y(ori_ori_n917_));
  NA2        o0889(.A(ori_ori_n581_), .B(ori_ori_n109_), .Y(ori_ori_n918_));
  OR3        o0890(.A(ori_ori_n304_), .B(ori_ori_n421_), .C(f), .Y(ori_ori_n919_));
  NA3        o0891(.A(ori_ori_n601_), .B(ori_ori_n76_), .C(i), .Y(ori_ori_n920_));
  OA220      o0892(.A0(ori_ori_n920_), .A1(ori_ori_n918_), .B0(ori_ori_n919_), .B1(ori_ori_n569_), .Y(ori_ori_n921_));
  NA3        o0893(.A(ori_ori_n319_), .B(ori_ori_n113_), .C(g), .Y(ori_ori_n922_));
  AOI210     o0894(.A0(ori_ori_n650_), .A1(ori_ori_n922_), .B0(m), .Y(ori_ori_n923_));
  OAI210     o0895(.A0(ori_ori_n923_), .A1(ori_ori_n875_), .B0(ori_ori_n318_), .Y(ori_ori_n924_));
  NA2        o0896(.A(ori_ori_n664_), .B(ori_ori_n827_), .Y(ori_ori_n925_));
  INV        o0897(.A(ori_ori_n795_), .Y(ori_ori_n926_));
  NA2        o0898(.A(ori_ori_n217_), .B(ori_ori_n73_), .Y(ori_ori_n927_));
  NA3        o0899(.A(ori_ori_n927_), .B(ori_ori_n920_), .C(ori_ori_n919_), .Y(ori_ori_n928_));
  AOI220     o0900(.A0(ori_ori_n928_), .A1(ori_ori_n254_), .B0(ori_ori_n926_), .B1(ori_ori_n925_), .Y(ori_ori_n929_));
  NA4        o0901(.A(ori_ori_n929_), .B(ori_ori_n924_), .C(ori_ori_n921_), .D(ori_ori_n917_), .Y(ori_ori_n930_));
  NO2        o0902(.A(ori_ori_n371_), .B(ori_ori_n87_), .Y(ori_ori_n931_));
  OAI210     o0903(.A0(ori_ori_n931_), .A1(ori_ori_n883_), .B0(ori_ori_n233_), .Y(ori_ori_n932_));
  NA2        o0904(.A(ori_ori_n639_), .B(ori_ori_n84_), .Y(ori_ori_n933_));
  NO2        o0905(.A(ori_ori_n442_), .B(ori_ori_n209_), .Y(ori_ori_n934_));
  AOI220     o0906(.A0(ori_ori_n934_), .A1(ori_ori_n374_), .B0(ori_ori_n887_), .B1(ori_ori_n213_), .Y(ori_ori_n935_));
  NA2        o0907(.A(ori_ori_n568_), .B(ori_ori_n86_), .Y(ori_ori_n936_));
  NA4        o0908(.A(ori_ori_n936_), .B(ori_ori_n935_), .C(ori_ori_n933_), .D(ori_ori_n932_), .Y(ori_ori_n937_));
  OAI210     o0909(.A0(ori_ori_n926_), .A1(ori_ori_n884_), .B0(ori_ori_n524_), .Y(ori_ori_n938_));
  NA2        o0910(.A(ori_ori_n923_), .B(ori_ori_n874_), .Y(ori_ori_n939_));
  NO3        o0911(.A(ori_ori_n839_), .B(ori_ori_n49_), .C(ori_ori_n45_), .Y(ori_ori_n940_));
  AOI220     o0912(.A0(ori_ori_n940_), .A1(ori_ori_n599_), .B0(ori_ori_n620_), .B1(ori_ori_n513_), .Y(ori_ori_n941_));
  NA3        o0913(.A(ori_ori_n941_), .B(ori_ori_n939_), .C(ori_ori_n938_), .Y(ori_ori_n942_));
  NO4        o0914(.A(ori_ori_n942_), .B(ori_ori_n937_), .C(ori_ori_n930_), .D(ori_ori_n913_), .Y(ori_ori_n943_));
  NAi31      o0915(.An(ori_ori_n135_), .B(ori_ori_n411_), .C(n), .Y(ori_ori_n944_));
  NO2        o0916(.A(ori_ori_n120_), .B(ori_ori_n332_), .Y(ori_ori_n945_));
  NO2        o0917(.A(ori_ori_n945_), .B(ori_ori_n944_), .Y(ori_ori_n946_));
  NO3        o0918(.A(ori_ori_n268_), .B(ori_ori_n135_), .C(ori_ori_n400_), .Y(ori_ori_n947_));
  AOI210     o0919(.A0(ori_ori_n947_), .A1(ori_ori_n482_), .B0(ori_ori_n946_), .Y(ori_ori_n948_));
  NA2        o0920(.A(ori_ori_n475_), .B(i), .Y(ori_ori_n949_));
  NA2        o0921(.A(ori_ori_n949_), .B(ori_ori_n948_), .Y(ori_ori_n950_));
  NA2        o0922(.A(ori_ori_n226_), .B(ori_ori_n166_), .Y(ori_ori_n951_));
  NO3        o0923(.A(ori_ori_n302_), .B(ori_ori_n427_), .C(ori_ori_n170_), .Y(ori_ori_n952_));
  NOi31      o0924(.An(ori_ori_n951_), .B(ori_ori_n952_), .C(ori_ori_n209_), .Y(ori_ori_n953_));
  NAi21      o0925(.An(ori_ori_n536_), .B(ori_ori_n934_), .Y(ori_ori_n954_));
  NA2        o0926(.A(ori_ori_n466_), .B(g), .Y(ori_ori_n955_));
  NA2        o0927(.A(ori_ori_n955_), .B(ori_ori_n954_), .Y(ori_ori_n956_));
  OAI220     o0928(.A0(ori_ori_n944_), .A1(ori_ori_n229_), .B0(ori_ori_n915_), .B1(ori_ori_n577_), .Y(ori_ori_n957_));
  NO2        o0929(.A(ori_ori_n636_), .B(ori_ori_n371_), .Y(ori_ori_n958_));
  NA2        o0930(.A(ori_ori_n879_), .B(ori_ori_n870_), .Y(ori_ori_n959_));
  OAI220     o0931(.A0(ori_ori_n876_), .A1(ori_ori_n884_), .B0(ori_ori_n526_), .B1(ori_ori_n417_), .Y(ori_ori_n960_));
  NA3        o0932(.A(ori_ori_n960_), .B(ori_ori_n959_), .C(ori_ori_n593_), .Y(ori_ori_n961_));
  OAI210     o0933(.A0(ori_ori_n879_), .A1(ori_ori_n871_), .B0(ori_ori_n951_), .Y(ori_ori_n962_));
  NA3        o0934(.A(ori_ori_n911_), .B(ori_ori_n471_), .C(ori_ori_n46_), .Y(ori_ori_n963_));
  INV        o0935(.A(ori_ori_n322_), .Y(ori_ori_n964_));
  NA4        o0936(.A(ori_ori_n964_), .B(ori_ori_n963_), .C(ori_ori_n962_), .D(ori_ori_n269_), .Y(ori_ori_n965_));
  OR4        o0937(.A(ori_ori_n965_), .B(ori_ori_n961_), .C(ori_ori_n958_), .D(ori_ori_n957_), .Y(ori_ori_n966_));
  NO4        o0938(.A(ori_ori_n966_), .B(ori_ori_n956_), .C(ori_ori_n953_), .D(ori_ori_n950_), .Y(ori_ori_n967_));
  NA4        o0939(.A(ori_ori_n967_), .B(ori_ori_n943_), .C(ori_ori_n905_), .D(ori_ori_n892_), .Y(ori13));
  NAi32      o0940(.An(d), .Bn(c), .C(e), .Y(ori_ori_n969_));
  AN2        o0941(.A(d), .B(c), .Y(ori_ori_n970_));
  NA2        o0942(.A(ori_ori_n970_), .B(ori_ori_n111_), .Y(ori_ori_n971_));
  NO3        o0943(.A(m), .B(i), .C(h), .Y(ori_ori_n972_));
  NA3        o0944(.A(k), .B(j), .C(i), .Y(ori_ori_n973_));
  NO2        o0945(.A(f), .B(c), .Y(ori_ori_n974_));
  NOi21      o0946(.An(ori_ori_n974_), .B(ori_ori_n426_), .Y(ori_ori_n975_));
  AN3        o0947(.A(g), .B(f), .C(c), .Y(ori_ori_n976_));
  NA3        o0948(.A(l), .B(k), .C(j), .Y(ori_ori_n977_));
  NA2        o0949(.A(i), .B(h), .Y(ori_ori_n978_));
  NO3        o0950(.A(ori_ori_n978_), .B(ori_ori_n977_), .C(ori_ori_n127_), .Y(ori_ori_n979_));
  NO3        o0951(.A(ori_ori_n136_), .B(ori_ori_n280_), .C(ori_ori_n209_), .Y(ori_ori_n980_));
  NA3        o0952(.A(c), .B(b), .C(a), .Y(ori_ori_n981_));
  NO2        o0953(.A(ori_ori_n509_), .B(ori_ori_n574_), .Y(ori_ori_n982_));
  NA4        o0954(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(g), .D(ori_ori_n208_), .Y(ori_ori_n983_));
  NA4        o0955(.A(ori_ori_n555_), .B(m), .C(ori_ori_n108_), .D(ori_ori_n208_), .Y(ori_ori_n984_));
  NA3        o0956(.A(ori_ori_n984_), .B(ori_ori_n362_), .C(ori_ori_n983_), .Y(ori_ori_n985_));
  NO2        o0957(.A(ori_ori_n985_), .B(ori_ori_n982_), .Y(ori_ori_n986_));
  NOi41      o0958(.An(ori_ori_n763_), .B(ori_ori_n806_), .C(ori_ori_n796_), .D(ori_ori_n689_), .Y(ori_ori_n987_));
  OAI220     o0959(.A0(ori_ori_n987_), .A1(ori_ori_n664_), .B0(ori_ori_n986_), .B1(ori_ori_n567_), .Y(ori_ori_n988_));
  NOi31      o0960(.An(m), .B(n), .C(f), .Y(ori_ori_n989_));
  NA2        o0961(.A(ori_ori_n989_), .B(ori_ori_n51_), .Y(ori_ori_n990_));
  NA2        o0962(.A(ori_ori_n490_), .B(l), .Y(ori_ori_n991_));
  NO2        o0963(.A(ori_ori_n280_), .B(a), .Y(ori_ori_n992_));
  NO2        o0964(.A(ori_ori_n83_), .B(g), .Y(ori_ori_n993_));
  NO3        o0965(.A(ori_ori_n988_), .B(ori_ori_n778_), .C(ori_ori_n544_), .Y(ori_ori_n994_));
  NA2        o0966(.A(c), .B(b), .Y(ori_ori_n995_));
  NO2        o0967(.A(ori_ori_n674_), .B(ori_ori_n995_), .Y(ori_ori_n996_));
  OAI210     o0968(.A0(ori_ori_n814_), .A1(ori_ori_n787_), .B0(ori_ori_n405_), .Y(ori_ori_n997_));
  OAI210     o0969(.A0(ori_ori_n997_), .A1(ori_ori_n815_), .B0(ori_ori_n996_), .Y(ori_ori_n998_));
  NAi21      o0970(.An(ori_ori_n413_), .B(ori_ori_n996_), .Y(ori_ori_n999_));
  NA3        o0971(.A(ori_ori_n417_), .B(ori_ori_n541_), .C(f), .Y(ori_ori_n1000_));
  NA2        o0972(.A(ori_ori_n530_), .B(ori_ori_n992_), .Y(ori_ori_n1001_));
  NA3        o0973(.A(ori_ori_n1001_), .B(ori_ori_n1000_), .C(ori_ori_n999_), .Y(ori_ori_n1002_));
  NA2        o0974(.A(ori_ori_n257_), .B(ori_ori_n114_), .Y(ori_ori_n1003_));
  OAI210     o0975(.A0(ori_ori_n1003_), .A1(ori_ori_n283_), .B0(g), .Y(ori_ori_n1004_));
  NAi21      o0976(.An(f), .B(d), .Y(ori_ori_n1005_));
  NO2        o0977(.A(ori_ori_n1005_), .B(ori_ori_n981_), .Y(ori_ori_n1006_));
  INV        o0978(.A(ori_ori_n1006_), .Y(ori_ori_n1007_));
  NO2        o0979(.A(ori_ori_n1004_), .B(ori_ori_n1007_), .Y(ori_ori_n1008_));
  AOI210     o0980(.A0(ori_ori_n1008_), .A1(ori_ori_n109_), .B0(ori_ori_n1002_), .Y(ori_ori_n1009_));
  NA2        o0981(.A(ori_ori_n452_), .B(ori_ori_n451_), .Y(ori_ori_n1010_));
  NO2        o0982(.A(ori_ori_n177_), .B(ori_ori_n232_), .Y(ori_ori_n1011_));
  NA2        o0983(.A(ori_ori_n1011_), .B(m), .Y(ori_ori_n1012_));
  NA2        o0984(.A(ori_ori_n991_), .B(ori_ori_n455_), .Y(ori_ori_n1013_));
  OAI210     o0985(.A0(ori_ori_n1013_), .A1(ori_ori_n305_), .B0(ori_ori_n453_), .Y(ori_ori_n1014_));
  AOI210     o0986(.A0(ori_ori_n1014_), .A1(ori_ori_n1010_), .B0(ori_ori_n1012_), .Y(ori_ori_n1015_));
  NA2        o0987(.A(ori_ori_n430_), .B(ori_ori_n1006_), .Y(ori_ori_n1016_));
  NO2        o0988(.A(ori_ori_n365_), .B(ori_ori_n364_), .Y(ori_ori_n1017_));
  NA2        o0989(.A(ori_ori_n1011_), .B(ori_ori_n419_), .Y(ori_ori_n1018_));
  NAi31      o0990(.An(ori_ori_n1017_), .B(ori_ori_n1018_), .C(ori_ori_n1016_), .Y(ori_ori_n1019_));
  NO2        o0991(.A(ori_ori_n1019_), .B(ori_ori_n1015_), .Y(ori_ori_n1020_));
  NA4        o0992(.A(ori_ori_n1020_), .B(ori_ori_n1009_), .C(ori_ori_n998_), .D(ori_ori_n994_), .Y(ori00));
  AOI210     o0993(.A0(ori_ori_n292_), .A1(ori_ori_n209_), .B0(ori_ori_n272_), .Y(ori_ori_n1022_));
  NO2        o0994(.A(ori_ori_n1022_), .B(ori_ori_n558_), .Y(ori_ori_n1023_));
  NA2        o0995(.A(ori_ori_n492_), .B(f), .Y(ori_ori_n1024_));
  OAI210     o0996(.A0(ori_ori_n945_), .A1(ori_ori_n40_), .B0(ori_ori_n622_), .Y(ori_ori_n1025_));
  NA3        o0997(.A(ori_ori_n1025_), .B(ori_ori_n253_), .C(n), .Y(ori_ori_n1026_));
  AOI210     o0998(.A0(ori_ori_n1026_), .A1(ori_ori_n1024_), .B0(ori_ori_n971_), .Y(ori_ori_n1027_));
  NO3        o0999(.A(ori_ori_n1027_), .B(ori_ori_n686_), .C(ori_ori_n1023_), .Y(ori_ori_n1028_));
  NA3        o1000(.A(d), .B(ori_ori_n56_), .C(b), .Y(ori_ori_n1029_));
  INV        o1001(.A(ori_ori_n557_), .Y(ori_ori_n1030_));
  NO3        o1002(.A(ori_ori_n1030_), .B(ori_ori_n1017_), .C(ori_ori_n862_), .Y(ori_ori_n1031_));
  NO4        o1003(.A(ori_ori_n472_), .B(ori_ori_n348_), .C(ori_ori_n995_), .D(ori_ori_n59_), .Y(ori_ori_n1032_));
  NA3        o1004(.A(ori_ori_n375_), .B(ori_ori_n216_), .C(g), .Y(ori_ori_n1033_));
  OA220      o1005(.A0(ori_ori_n1033_), .A1(ori_ori_n1029_), .B0(ori_ori_n376_), .B1(ori_ori_n128_), .Y(ori_ori_n1034_));
  NO2        o1006(.A(h), .B(g), .Y(ori_ori_n1035_));
  OAI220     o1007(.A0(ori_ori_n509_), .A1(ori_ori_n574_), .B0(ori_ori_n88_), .B1(ori_ori_n87_), .Y(ori_ori_n1036_));
  NA2        o1008(.A(ori_ori_n1036_), .B(ori_ori_n517_), .Y(ori_ori_n1037_));
  AOI220     o1009(.A0(ori_ori_n311_), .A1(ori_ori_n242_), .B0(ori_ori_n172_), .B1(ori_ori_n143_), .Y(ori_ori_n1038_));
  NA3        o1010(.A(ori_ori_n1038_), .B(ori_ori_n1037_), .C(ori_ori_n1034_), .Y(ori_ori_n1039_));
  NO3        o1011(.A(ori_ori_n1039_), .B(ori_ori_n1032_), .C(ori_ori_n263_), .Y(ori_ori_n1040_));
  INV        o1012(.A(ori_ori_n316_), .Y(ori_ori_n1041_));
  AOI210     o1013(.A0(ori_ori_n242_), .A1(ori_ori_n339_), .B0(ori_ori_n559_), .Y(ori_ori_n1042_));
  NA3        o1014(.A(ori_ori_n1042_), .B(ori_ori_n1041_), .C(ori_ori_n149_), .Y(ori_ori_n1043_));
  NO2        o1015(.A(ori_ori_n1043_), .B(ori_ori_n500_), .Y(ori_ori_n1044_));
  AN3        o1016(.A(ori_ori_n1044_), .B(ori_ori_n1040_), .C(ori_ori_n1031_), .Y(ori_ori_n1045_));
  NA2        o1017(.A(ori_ori_n517_), .B(ori_ori_n98_), .Y(ori_ori_n1046_));
  NA3        o1018(.A(ori_ori_n989_), .B(ori_ori_n581_), .C(ori_ori_n449_), .Y(ori_ori_n1047_));
  NA3        o1019(.A(ori_ori_n1047_), .B(ori_ori_n1046_), .C(ori_ori_n236_), .Y(ori_ori_n1048_));
  NA2        o1020(.A(ori_ori_n985_), .B(ori_ori_n517_), .Y(ori_ori_n1049_));
  NA4        o1021(.A(ori_ori_n625_), .B(ori_ori_n201_), .C(ori_ori_n216_), .D(ori_ori_n158_), .Y(ori_ori_n1050_));
  NA2        o1022(.A(ori_ori_n1050_), .B(ori_ori_n1049_), .Y(ori_ori_n1051_));
  OAI210     o1023(.A0(ori_ori_n448_), .A1(ori_ori_n115_), .B0(ori_ori_n817_), .Y(ori_ori_n1052_));
  NA2        o1024(.A(ori_ori_n1052_), .B(ori_ori_n1013_), .Y(ori_ori_n1053_));
  NO2        o1025(.A(ori_ori_n212_), .B(ori_ori_n209_), .Y(ori_ori_n1054_));
  NA2        o1026(.A(n), .B(e), .Y(ori_ori_n1055_));
  NO2        o1027(.A(ori_ori_n1055_), .B(ori_ori_n141_), .Y(ori_ori_n1056_));
  AOI220     o1028(.A0(ori_ori_n1056_), .A1(ori_ori_n270_), .B0(ori_ori_n800_), .B1(ori_ori_n1054_), .Y(ori_ori_n1057_));
  OAI210     o1029(.A0(ori_ori_n349_), .A1(ori_ori_n306_), .B0(ori_ori_n432_), .Y(ori_ori_n1058_));
  NA3        o1030(.A(ori_ori_n1058_), .B(ori_ori_n1057_), .C(ori_ori_n1053_), .Y(ori_ori_n1059_));
  NA2        o1031(.A(ori_ori_n1056_), .B(ori_ori_n803_), .Y(ori_ori_n1060_));
  AOI220     o1032(.A0(ori_ori_n896_), .A1(ori_ori_n556_), .B0(ori_ori_n625_), .B1(ori_ori_n239_), .Y(ori_ori_n1061_));
  NO2        o1033(.A(ori_ori_n64_), .B(h), .Y(ori_ori_n1062_));
  NA3        o1034(.A(ori_ori_n1061_), .B(ori_ori_n1060_), .C(ori_ori_n819_), .Y(ori_ori_n1063_));
  NO4        o1035(.A(ori_ori_n1063_), .B(ori_ori_n1059_), .C(ori_ori_n1051_), .D(ori_ori_n1048_), .Y(ori_ori_n1064_));
  NA2        o1036(.A(ori_ori_n788_), .B(ori_ori_n722_), .Y(ori_ori_n1065_));
  NA4        o1037(.A(ori_ori_n1065_), .B(ori_ori_n1064_), .C(ori_ori_n1045_), .D(ori_ori_n1028_), .Y(ori01));
  NO2        o1038(.A(ori_ori_n463_), .B(ori_ori_n278_), .Y(ori_ori_n1067_));
  NA2        o1039(.A(ori_ori_n386_), .B(i), .Y(ori_ori_n1068_));
  NA3        o1040(.A(ori_ori_n1068_), .B(ori_ori_n1067_), .C(ori_ori_n959_), .Y(ori_ori_n1069_));
  NA2        o1041(.A(ori_ori_n568_), .B(ori_ori_n86_), .Y(ori_ori_n1070_));
  NA2        o1042(.A(ori_ori_n536_), .B(ori_ori_n267_), .Y(ori_ori_n1071_));
  NA2        o1043(.A(ori_ori_n901_), .B(ori_ori_n1071_), .Y(ori_ori_n1072_));
  NA4        o1044(.A(ori_ori_n1072_), .B(ori_ori_n1070_), .C(ori_ori_n857_), .D(ori_ori_n324_), .Y(ori_ori_n1073_));
  NA2        o1045(.A(ori_ori_n45_), .B(f), .Y(ori_ori_n1074_));
  NA2        o1046(.A(ori_ori_n681_), .B(ori_ori_n93_), .Y(ori_ori_n1075_));
  NO2        o1047(.A(ori_ori_n1075_), .B(ori_ori_n1074_), .Y(ori_ori_n1076_));
  OAI210     o1048(.A0(ori_ori_n742_), .A1(ori_ori_n577_), .B0(ori_ori_n1050_), .Y(ori_ori_n1077_));
  AOI210     o1049(.A0(ori_ori_n1076_), .A1(ori_ori_n610_), .B0(ori_ori_n1077_), .Y(ori_ori_n1078_));
  OR2        o1050(.A(ori_ori_n637_), .B(ori_ori_n362_), .Y(ori_ori_n1079_));
  NAi41      o1051(.An(ori_ori_n157_), .B(ori_ori_n1079_), .C(ori_ori_n1078_), .D(ori_ori_n843_), .Y(ori_ori_n1080_));
  NO2        o1052(.A(ori_ori_n652_), .B(ori_ori_n495_), .Y(ori_ori_n1081_));
  NA4        o1053(.A(ori_ori_n681_), .B(ori_ori_n93_), .C(ori_ori_n45_), .D(ori_ori_n208_), .Y(ori_ori_n1082_));
  OA220      o1054(.A0(ori_ori_n1082_), .A1(ori_ori_n645_), .B0(ori_ori_n190_), .B1(ori_ori_n188_), .Y(ori_ori_n1083_));
  NA3        o1055(.A(ori_ori_n1083_), .B(ori_ori_n1081_), .C(ori_ori_n131_), .Y(ori_ori_n1084_));
  NO4        o1056(.A(ori_ori_n1084_), .B(ori_ori_n1080_), .C(ori_ori_n1073_), .D(ori_ori_n1069_), .Y(ori_ori_n1085_));
  INV        o1057(.A(ori_ori_n1033_), .Y(ori_ori_n1086_));
  OAI210     o1058(.A0(ori_ori_n1086_), .A1(ori_ori_n295_), .B0(ori_ori_n513_), .Y(ori_ori_n1087_));
  AOI210     o1059(.A0(ori_ori_n199_), .A1(ori_ori_n85_), .B0(ori_ori_n208_), .Y(ori_ori_n1088_));
  OAI210     o1060(.A0(ori_ori_n766_), .A1(ori_ori_n417_), .B0(ori_ori_n1088_), .Y(ori_ori_n1089_));
  AN3        o1061(.A(m), .B(l), .C(k), .Y(ori_ori_n1090_));
  OAI210     o1062(.A0(ori_ori_n350_), .A1(ori_ori_n34_), .B0(ori_ori_n1090_), .Y(ori_ori_n1091_));
  OR2        o1063(.A(ori_ori_n1091_), .B(ori_ori_n323_), .Y(ori_ori_n1092_));
  NA3        o1064(.A(ori_ori_n1092_), .B(ori_ori_n1089_), .C(ori_ori_n1087_), .Y(ori_ori_n1093_));
  NA2        o1065(.A(ori_ori_n573_), .B(ori_ori_n113_), .Y(ori_ori_n1094_));
  INV        o1066(.A(ori_ori_n1094_), .Y(ori_ori_n1095_));
  NA2        o1067(.A(ori_ori_n277_), .B(ori_ori_n190_), .Y(ori_ori_n1096_));
  NA2        o1068(.A(ori_ori_n1096_), .B(ori_ori_n642_), .Y(ori_ori_n1097_));
  NA2        o1069(.A(ori_ori_n1076_), .B(ori_ori_n653_), .Y(ori_ori_n1098_));
  NA3        o1070(.A(ori_ori_n1098_), .B(ori_ori_n1097_), .C(ori_ori_n745_), .Y(ori_ori_n1099_));
  NO3        o1071(.A(ori_ori_n1099_), .B(ori_ori_n1095_), .C(ori_ori_n1093_), .Y(ori_ori_n1100_));
  NA3        o1072(.A(ori_ori_n578_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n1101_));
  NO2        o1073(.A(ori_ori_n1101_), .B(ori_ori_n199_), .Y(ori_ori_n1102_));
  AOI210     o1074(.A0(ori_ori_n489_), .A1(ori_ori_n58_), .B0(ori_ori_n1102_), .Y(ori_ori_n1103_));
  OR3        o1075(.A(ori_ori_n1075_), .B(ori_ori_n579_), .C(ori_ori_n1074_), .Y(ori_ori_n1104_));
  NO2        o1076(.A(ori_ori_n1082_), .B(ori_ori_n918_), .Y(ori_ori_n1105_));
  NO2        o1077(.A(ori_ori_n202_), .B(ori_ori_n107_), .Y(ori_ori_n1106_));
  NO2        o1078(.A(ori_ori_n1106_), .B(ori_ori_n1105_), .Y(ori_ori_n1107_));
  NA4        o1079(.A(ori_ori_n1107_), .B(ori_ori_n1104_), .C(ori_ori_n1103_), .D(ori_ori_n721_), .Y(ori_ori_n1108_));
  NO2        o1080(.A(ori_ori_n907_), .B(ori_ori_n228_), .Y(ori_ori_n1109_));
  NO2        o1081(.A(ori_ori_n908_), .B(ori_ori_n538_), .Y(ori_ori_n1110_));
  OAI210     o1082(.A0(ori_ori_n1110_), .A1(ori_ori_n1109_), .B0(ori_ori_n332_), .Y(ori_ori_n1111_));
  NA2        o1083(.A(ori_ori_n551_), .B(ori_ori_n549_), .Y(ori_ori_n1112_));
  NO3        o1084(.A(ori_ori_n75_), .B(ori_ori_n293_), .C(ori_ori_n45_), .Y(ori_ori_n1113_));
  NA2        o1085(.A(ori_ori_n1113_), .B(ori_ori_n535_), .Y(ori_ori_n1114_));
  NA3        o1086(.A(ori_ori_n1114_), .B(ori_ori_n1112_), .C(ori_ori_n647_), .Y(ori_ori_n1115_));
  OR2        o1087(.A(ori_ori_n1033_), .B(ori_ori_n1029_), .Y(ori_ori_n1116_));
  NO2        o1088(.A(ori_ori_n362_), .B(ori_ori_n68_), .Y(ori_ori_n1117_));
  INV        o1089(.A(ori_ori_n1117_), .Y(ori_ori_n1118_));
  NA2        o1090(.A(ori_ori_n1113_), .B(ori_ori_n769_), .Y(ori_ori_n1119_));
  NA4        o1091(.A(ori_ori_n1119_), .B(ori_ori_n1118_), .C(ori_ori_n1116_), .D(ori_ori_n378_), .Y(ori_ori_n1120_));
  NOi41      o1092(.An(ori_ori_n1111_), .B(ori_ori_n1120_), .C(ori_ori_n1115_), .D(ori_ori_n1108_), .Y(ori_ori_n1121_));
  NO2        o1093(.A(ori_ori_n126_), .B(ori_ori_n45_), .Y(ori_ori_n1122_));
  NO2        o1094(.A(ori_ori_n45_), .B(ori_ori_n40_), .Y(ori_ori_n1123_));
  AO220      o1095(.A0(ori_ori_n1123_), .A1(ori_ori_n596_), .B0(ori_ori_n1122_), .B1(ori_ori_n679_), .Y(ori_ori_n1124_));
  NA2        o1096(.A(ori_ori_n1124_), .B(ori_ori_n332_), .Y(ori_ori_n1125_));
  INV        o1097(.A(ori_ori_n128_), .Y(ori_ori_n1126_));
  NO3        o1098(.A(ori_ori_n978_), .B(ori_ori_n171_), .C(ori_ori_n83_), .Y(ori_ori_n1127_));
  NA2        o1099(.A(ori_ori_n1127_), .B(ori_ori_n1126_), .Y(ori_ori_n1128_));
  NA2        o1100(.A(ori_ori_n1128_), .B(ori_ori_n1125_), .Y(ori_ori_n1129_));
  NO2        o1101(.A(ori_ori_n589_), .B(ori_ori_n588_), .Y(ori_ori_n1130_));
  NO4        o1102(.A(ori_ori_n978_), .B(ori_ori_n1130_), .C(ori_ori_n169_), .D(ori_ori_n83_), .Y(ori_ori_n1131_));
  NO3        o1103(.A(ori_ori_n1131_), .B(ori_ori_n1129_), .C(ori_ori_n614_), .Y(ori_ori_n1132_));
  NA4        o1104(.A(ori_ori_n1132_), .B(ori_ori_n1121_), .C(ori_ori_n1100_), .D(ori_ori_n1085_), .Y(ori06));
  NO2        o1105(.A(ori_ori_n220_), .B(ori_ori_n100_), .Y(ori_ori_n1134_));
  OAI210     o1106(.A0(ori_ori_n1134_), .A1(ori_ori_n1127_), .B0(ori_ori_n374_), .Y(ori_ori_n1135_));
  NO3        o1107(.A(ori_ori_n575_), .B(ori_ori_n764_), .C(ori_ori_n576_), .Y(ori_ori_n1136_));
  OR2        o1108(.A(ori_ori_n1136_), .B(ori_ori_n833_), .Y(ori_ori_n1137_));
  NA3        o1109(.A(ori_ori_n1137_), .B(ori_ori_n1135_), .C(ori_ori_n1111_), .Y(ori_ori_n1138_));
  NO3        o1110(.A(ori_ori_n1138_), .B(ori_ori_n1115_), .C(ori_ori_n252_), .Y(ori_ori_n1139_));
  NO2        o1111(.A(ori_ori_n293_), .B(ori_ori_n45_), .Y(ori_ori_n1140_));
  AOI210     o1112(.A0(ori_ori_n1140_), .A1(ori_ori_n535_), .B0(ori_ori_n1109_), .Y(ori_ori_n1141_));
  AOI210     o1113(.A0(ori_ori_n1140_), .A1(ori_ori_n539_), .B0(ori_ori_n1124_), .Y(ori_ori_n1142_));
  AOI210     o1114(.A0(ori_ori_n1142_), .A1(ori_ori_n1141_), .B0(ori_ori_n329_), .Y(ori_ori_n1143_));
  OAI210     o1115(.A0(ori_ori_n85_), .A1(ori_ori_n40_), .B0(ori_ori_n651_), .Y(ori_ori_n1144_));
  NA2        o1116(.A(ori_ori_n1144_), .B(ori_ori_n618_), .Y(ori_ori_n1145_));
  NO2        o1117(.A(ori_ori_n497_), .B(ori_ori_n166_), .Y(ori_ori_n1146_));
  NOi21      o1118(.An(ori_ori_n130_), .B(ori_ori_n45_), .Y(ori_ori_n1147_));
  NO2        o1119(.A(ori_ori_n582_), .B(ori_ori_n990_), .Y(ori_ori_n1148_));
  NO3        o1120(.A(ori_ori_n1148_), .B(ori_ori_n1147_), .C(ori_ori_n1146_), .Y(ori_ori_n1149_));
  NA2        o1121(.A(ori_ori_n1149_), .B(ori_ori_n1145_), .Y(ori_ori_n1150_));
  NO2        o1122(.A(ori_ori_n713_), .B(ori_ori_n360_), .Y(ori_ori_n1151_));
  NO2        o1123(.A(ori_ori_n653_), .B(ori_ori_n610_), .Y(ori_ori_n1152_));
  NOi21      o1124(.An(ori_ori_n1151_), .B(ori_ori_n1152_), .Y(ori_ori_n1153_));
  AN2        o1125(.A(ori_ori_n896_), .B(ori_ori_n621_), .Y(ori_ori_n1154_));
  NO4        o1126(.A(ori_ori_n1154_), .B(ori_ori_n1153_), .C(ori_ori_n1150_), .D(ori_ori_n1143_), .Y(ori_ori_n1155_));
  NO2        o1127(.A(ori_ori_n704_), .B(ori_ori_n47_), .Y(ori_ori_n1156_));
  NA2        o1128(.A(ori_ori_n353_), .B(ori_ori_n1156_), .Y(ori_ori_n1157_));
  NO3        o1129(.A(ori_ori_n238_), .B(ori_ori_n100_), .C(ori_ori_n280_), .Y(ori_ori_n1158_));
  OAI220     o1130(.A0(ori_ori_n671_), .A1(ori_ori_n243_), .B0(ori_ori_n494_), .B1(ori_ori_n497_), .Y(ori_ori_n1159_));
  INV        o1131(.A(k), .Y(ori_ori_n1160_));
  NO3        o1132(.A(ori_ori_n1160_), .B(ori_ori_n574_), .C(j), .Y(ori_ori_n1161_));
  NOi21      o1133(.An(ori_ori_n1161_), .B(ori_ori_n645_), .Y(ori_ori_n1162_));
  NO3        o1134(.A(ori_ori_n1162_), .B(ori_ori_n1159_), .C(ori_ori_n1158_), .Y(ori_ori_n1163_));
  NA4        o1135(.A(ori_ori_n753_), .B(ori_ori_n752_), .C(ori_ori_n424_), .D(ori_ori_n827_), .Y(ori_ori_n1164_));
  NAi31      o1136(.An(ori_ori_n713_), .B(ori_ori_n1164_), .C(ori_ori_n198_), .Y(ori_ori_n1165_));
  NA4        o1137(.A(ori_ori_n1165_), .B(ori_ori_n1163_), .C(ori_ori_n1157_), .D(ori_ori_n1061_), .Y(ori_ori_n1166_));
  AOI210     o1138(.A0(ori_ori_n551_), .A1(ori_ori_n432_), .B0(ori_ori_n366_), .Y(ori_ori_n1167_));
  NA2        o1139(.A(ori_ori_n1161_), .B(ori_ori_n749_), .Y(ori_ori_n1168_));
  NA2        o1140(.A(ori_ori_n1168_), .B(ori_ori_n1167_), .Y(ori_ori_n1169_));
  AN2        o1141(.A(ori_ori_n871_), .B(ori_ori_n870_), .Y(ori_ori_n1170_));
  NO3        o1142(.A(ori_ori_n1170_), .B(ori_ori_n485_), .C(ori_ori_n466_), .Y(ori_ori_n1171_));
  NA2        o1143(.A(ori_ori_n1171_), .B(ori_ori_n1119_), .Y(ori_ori_n1172_));
  NAi21      o1144(.An(j), .B(i), .Y(ori_ori_n1173_));
  NO4        o1145(.A(ori_ori_n1130_), .B(ori_ori_n1173_), .C(ori_ori_n426_), .D(ori_ori_n230_), .Y(ori_ori_n1174_));
  NO4        o1146(.A(ori_ori_n1174_), .B(ori_ori_n1172_), .C(ori_ori_n1169_), .D(ori_ori_n1166_), .Y(ori_ori_n1175_));
  NA4        o1147(.A(ori_ori_n1175_), .B(ori_ori_n1155_), .C(ori_ori_n1139_), .D(ori_ori_n1132_), .Y(ori07));
  NAi32      o1148(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1177_));
  NO3        o1149(.A(ori_ori_n1177_), .B(g), .C(f), .Y(ori_ori_n1178_));
  NAi21      o1150(.An(f), .B(c), .Y(ori_ori_n1179_));
  OR2        o1151(.A(e), .B(d), .Y(ori_ori_n1180_));
  NOi31      o1152(.An(n), .B(m), .C(b), .Y(ori_ori_n1181_));
  NOi41      o1153(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1182_));
  NO2        o1154(.A(ori_ori_n973_), .B(ori_ori_n301_), .Y(ori_ori_n1183_));
  NA2        o1155(.A(ori_ori_n523_), .B(ori_ori_n76_), .Y(ori_ori_n1184_));
  NA2        o1156(.A(ori_ori_n1062_), .B(ori_ori_n287_), .Y(ori_ori_n1185_));
  NA2        o1157(.A(ori_ori_n1185_), .B(ori_ori_n1184_), .Y(ori_ori_n1186_));
  NO2        o1158(.A(ori_ori_n1186_), .B(ori_ori_n1178_), .Y(ori_ori_n1187_));
  NO3        o1159(.A(e), .B(d), .C(c), .Y(ori_ori_n1188_));
  NO2        o1160(.A(ori_ori_n127_), .B(ori_ori_n209_), .Y(ori_ori_n1189_));
  NA2        o1161(.A(ori_ori_n1189_), .B(ori_ori_n1188_), .Y(ori_ori_n1190_));
  INV        o1162(.A(ori_ori_n1190_), .Y(ori_ori_n1191_));
  NA3        o1163(.A(ori_ori_n668_), .B(ori_ori_n656_), .C(ori_ori_n108_), .Y(ori_ori_n1192_));
  NO2        o1164(.A(ori_ori_n1192_), .B(ori_ori_n45_), .Y(ori_ori_n1193_));
  NO2        o1165(.A(l), .B(k), .Y(ori_ori_n1194_));
  NO3        o1166(.A(ori_ori_n426_), .B(d), .C(c), .Y(ori_ori_n1195_));
  NO2        o1167(.A(ori_ori_n1193_), .B(ori_ori_n1191_), .Y(ori_ori_n1196_));
  NO2        o1168(.A(g), .B(c), .Y(ori_ori_n1197_));
  NO2        o1169(.A(ori_ori_n434_), .B(a), .Y(ori_ori_n1198_));
  NA2        o1170(.A(ori_ori_n1198_), .B(ori_ori_n109_), .Y(ori_ori_n1199_));
  NA2        o1171(.A(ori_ori_n132_), .B(ori_ori_n216_), .Y(ori_ori_n1200_));
  NO2        o1172(.A(ori_ori_n1200_), .B(ori_ori_n1289_), .Y(ori_ori_n1201_));
  NO2        o1173(.A(ori_ori_n720_), .B(ori_ori_n182_), .Y(ori_ori_n1202_));
  NOi31      o1174(.An(m), .B(n), .C(b), .Y(ori_ori_n1203_));
  NOi31      o1175(.An(f), .B(d), .C(c), .Y(ori_ori_n1204_));
  NA2        o1176(.A(ori_ori_n1204_), .B(ori_ori_n1203_), .Y(ori_ori_n1205_));
  INV        o1177(.A(ori_ori_n1205_), .Y(ori_ori_n1206_));
  NO3        o1178(.A(ori_ori_n1206_), .B(ori_ori_n1202_), .C(ori_ori_n1201_), .Y(ori_ori_n1207_));
  NA2        o1179(.A(ori_ori_n976_), .B(ori_ori_n450_), .Y(ori_ori_n1208_));
  NO2        o1180(.A(ori_ori_n1208_), .B(ori_ori_n426_), .Y(ori_ori_n1209_));
  NO3        o1181(.A(ori_ori_n41_), .B(i), .C(h), .Y(ori_ori_n1210_));
  NO2        o1182(.A(ori_ori_n972_), .B(ori_ori_n1209_), .Y(ori_ori_n1211_));
  AN3        o1183(.A(ori_ori_n1211_), .B(ori_ori_n1207_), .C(ori_ori_n1199_), .Y(ori_ori_n1212_));
  NA2        o1184(.A(ori_ori_n1181_), .B(ori_ori_n372_), .Y(ori_ori_n1213_));
  INV        o1185(.A(ori_ori_n1213_), .Y(ori_ori_n1214_));
  INV        o1186(.A(ori_ori_n979_), .Y(ori_ori_n1215_));
  NAi21      o1187(.An(ori_ori_n1214_), .B(ori_ori_n1215_), .Y(ori_ori_n1216_));
  NO4        o1188(.A(ori_ori_n127_), .B(g), .C(f), .D(e), .Y(ori_ori_n1217_));
  NA2        o1189(.A(ori_ori_n1182_), .B(ori_ori_n1194_), .Y(ori_ori_n1218_));
  INV        o1190(.A(ori_ori_n1218_), .Y(ori_ori_n1219_));
  OR3        o1191(.A(ori_ori_n522_), .B(ori_ori_n521_), .C(ori_ori_n108_), .Y(ori_ori_n1220_));
  NA2        o1192(.A(ori_ori_n989_), .B(ori_ori_n400_), .Y(ori_ori_n1221_));
  NO2        o1193(.A(ori_ori_n1221_), .B(ori_ori_n423_), .Y(ori_ori_n1222_));
  AO210      o1194(.A0(ori_ori_n1222_), .A1(ori_ori_n111_), .B0(ori_ori_n1219_), .Y(ori_ori_n1223_));
  NO2        o1195(.A(ori_ori_n1223_), .B(ori_ori_n1216_), .Y(ori_ori_n1224_));
  NA4        o1196(.A(ori_ori_n1224_), .B(ori_ori_n1212_), .C(ori_ori_n1196_), .D(ori_ori_n1187_), .Y(ori_ori_n1225_));
  NO2        o1197(.A(ori_ori_n995_), .B(ori_ori_n106_), .Y(ori_ori_n1226_));
  NO2        o1198(.A(ori_ori_n383_), .B(j), .Y(ori_ori_n1227_));
  NA2        o1199(.A(ori_ori_n1210_), .B(ori_ori_n989_), .Y(ori_ori_n1228_));
  NA2        o1200(.A(ori_ori_n975_), .B(ori_ori_n145_), .Y(ori_ori_n1229_));
  NA2        o1201(.A(ori_ori_n1229_), .B(ori_ori_n1228_), .Y(ori_ori_n1230_));
  NA2        o1202(.A(ori_ori_n1227_), .B(ori_ori_n154_), .Y(ori_ori_n1231_));
  INV        o1203(.A(ori_ori_n1231_), .Y(ori_ori_n1232_));
  NO2        o1204(.A(ori_ori_n1232_), .B(ori_ori_n1230_), .Y(ori_ori_n1233_));
  INV        o1205(.A(ori_ori_n49_), .Y(ori_ori_n1234_));
  NA2        o1206(.A(ori_ori_n1234_), .B(ori_ori_n1035_), .Y(ori_ori_n1235_));
  INV        o1207(.A(ori_ori_n1235_), .Y(ori_ori_n1236_));
  NO2        o1208(.A(ori_ori_n643_), .B(ori_ori_n171_), .Y(ori_ori_n1237_));
  NO2        o1209(.A(ori_ori_n1237_), .B(ori_ori_n1236_), .Y(ori_ori_n1238_));
  NO3        o1210(.A(ori_ori_n981_), .B(ori_ori_n1180_), .C(ori_ori_n49_), .Y(ori_ori_n1239_));
  NA3        o1211(.A(ori_ori_n1226_), .B(ori_ori_n450_), .C(f), .Y(ori_ori_n1240_));
  INV        o1212(.A(ori_ori_n174_), .Y(ori_ori_n1241_));
  NO2        o1213(.A(ori_ori_n1288_), .B(ori_ori_n1240_), .Y(ori_ori_n1242_));
  NO2        o1214(.A(ori_ori_n1173_), .B(ori_ori_n169_), .Y(ori_ori_n1243_));
  NOi21      o1215(.An(d), .B(f), .Y(ori_ori_n1244_));
  NA2        o1216(.A(h), .B(ori_ori_n1243_), .Y(ori_ori_n1245_));
  INV        o1217(.A(ori_ori_n1245_), .Y(ori_ori_n1246_));
  NO2        o1218(.A(ori_ori_n1246_), .B(ori_ori_n1242_), .Y(ori_ori_n1247_));
  NA3        o1219(.A(ori_ori_n1247_), .B(ori_ori_n1238_), .C(ori_ori_n1233_), .Y(ori_ori_n1248_));
  NA2        o1220(.A(h), .B(ori_ori_n1183_), .Y(ori_ori_n1249_));
  OAI210     o1221(.A0(ori_ori_n1217_), .A1(ori_ori_n1181_), .B0(ori_ori_n830_), .Y(ori_ori_n1250_));
  NO2        o1222(.A(ori_ori_n969_), .B(ori_ori_n127_), .Y(ori_ori_n1251_));
  NA2        o1223(.A(ori_ori_n1251_), .B(ori_ori_n595_), .Y(ori_ori_n1252_));
  NA3        o1224(.A(ori_ori_n1252_), .B(ori_ori_n1250_), .C(ori_ori_n1249_), .Y(ori_ori_n1253_));
  NA2        o1225(.A(ori_ori_n1197_), .B(ori_ori_n1244_), .Y(ori_ori_n1254_));
  NO2        o1226(.A(ori_ori_n1254_), .B(m), .Y(ori_ori_n1255_));
  NO2        o1227(.A(ori_ori_n146_), .B(ori_ori_n176_), .Y(ori_ori_n1256_));
  OAI210     o1228(.A0(ori_ori_n1256_), .A1(ori_ori_n106_), .B0(ori_ori_n1203_), .Y(ori_ori_n1257_));
  INV        o1229(.A(ori_ori_n1257_), .Y(ori_ori_n1258_));
  NO3        o1230(.A(ori_ori_n1258_), .B(ori_ori_n1255_), .C(ori_ori_n1253_), .Y(ori_ori_n1259_));
  NO2        o1231(.A(ori_ori_n1179_), .B(e), .Y(ori_ori_n1260_));
  NA2        o1232(.A(ori_ori_n1260_), .B(ori_ori_n398_), .Y(ori_ori_n1261_));
  BUFFER     o1233(.A(ori_ori_n127_), .Y(ori_ori_n1262_));
  NO2        o1234(.A(ori_ori_n1262_), .B(ori_ori_n1261_), .Y(ori_ori_n1263_));
  NO2        o1235(.A(ori_ori_n1220_), .B(ori_ori_n346_), .Y(ori_ori_n1264_));
  NO2        o1236(.A(ori_ori_n1264_), .B(ori_ori_n1263_), .Y(ori_ori_n1265_));
  NO2        o1237(.A(ori_ori_n1195_), .B(ori_ori_n1239_), .Y(ori_ori_n1266_));
  INV        o1238(.A(ori_ori_n993_), .Y(ori_ori_n1267_));
  OAI210     o1239(.A0(ori_ori_n1267_), .A1(ori_ori_n65_), .B0(ori_ori_n1266_), .Y(ori_ori_n1268_));
  OR2        o1240(.A(h), .B(ori_ori_n521_), .Y(ori_ori_n1269_));
  NO2        o1241(.A(ori_ori_n1269_), .B(ori_ori_n169_), .Y(ori_ori_n1270_));
  NA2        o1242(.A(ori_ori_n980_), .B(ori_ori_n216_), .Y(ori_ori_n1271_));
  NO2        o1243(.A(ori_ori_n49_), .B(l), .Y(ori_ori_n1272_));
  INV        o1244(.A(ori_ori_n468_), .Y(ori_ori_n1273_));
  NA2        o1245(.A(ori_ori_n1273_), .B(ori_ori_n1272_), .Y(ori_ori_n1274_));
  NA2        o1246(.A(ori_ori_n1274_), .B(ori_ori_n1271_), .Y(ori_ori_n1275_));
  NO3        o1247(.A(ori_ori_n1275_), .B(ori_ori_n1270_), .C(ori_ori_n1268_), .Y(ori_ori_n1276_));
  NA3        o1248(.A(ori_ori_n1276_), .B(ori_ori_n1265_), .C(ori_ori_n1259_), .Y(ori_ori_n1277_));
  NA3        o1249(.A(ori_ori_n900_), .B(ori_ori_n132_), .C(ori_ori_n46_), .Y(ori_ori_n1278_));
  INV        o1250(.A(ori_ori_n1260_), .Y(ori_ori_n1279_));
  NO2        o1251(.A(ori_ori_n1279_), .B(ori_ori_n1241_), .Y(ori_ori_n1280_));
  INV        o1252(.A(ori_ori_n1280_), .Y(ori_ori_n1281_));
  NO2        o1253(.A(ori_ori_n1221_), .B(d), .Y(ori_ori_n1282_));
  INV        o1254(.A(ori_ori_n1282_), .Y(ori_ori_n1283_));
  NA3        o1255(.A(ori_ori_n1283_), .B(ori_ori_n1281_), .C(ori_ori_n1278_), .Y(ori_ori_n1284_));
  OR4        o1256(.A(ori_ori_n1284_), .B(ori_ori_n1277_), .C(ori_ori_n1248_), .D(ori_ori_n1225_), .Y(ori04));
  INV        o1257(.A(ori_ori_n109_), .Y(ori_ori_n1288_));
  INV        o1258(.A(h), .Y(ori_ori_n1289_));
  ZERO       o1259(.Y(ori02));
  ZERO       o1260(.Y(ori03));
  ZERO       o1261(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  INV        m0023(.A(mai_mai_n51_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO4        m0025(.A(mai_mai_n53_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n54_));
  AOI210     m0026(.A0(mai_mai_n54_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NA3        m0031(.A(g), .B(mai_mai_n59_), .C(a), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(h), .Y(mai_mai_n61_));
  NAi31      m0033(.An(i), .B(l), .C(j), .Y(mai_mai_n62_));
  OAI220     m0034(.A0(mai_mai_n62_), .A1(mai_mai_n49_), .B0(mai_mai_n61_), .B1(mai_mai_n44_), .Y(mai_mai_n63_));
  NAi31      m0035(.An(mai_mai_n60_), .B(mai_mai_n63_), .C(mai_mai_n58_), .Y(mai_mai_n64_));
  NAi41      m0036(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n65_));
  NA2        m0037(.A(g), .B(f), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi21      m0039(.An(i), .B(j), .Y(mai_mai_n68_));
  NAi32      m0040(.An(n), .Bn(k), .C(m), .Y(mai_mai_n69_));
  NO2        m0041(.A(mai_mai_n69_), .B(mai_mai_n68_), .Y(mai_mai_n70_));
  NAi31      m0042(.An(l), .B(m), .C(k), .Y(mai_mai_n71_));
  NAi41      m0043(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n72_));
  NA2        m0044(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n73_));
  INV        m0045(.A(m), .Y(mai_mai_n74_));
  NOi21      m0046(.An(k), .B(l), .Y(mai_mai_n75_));
  NA2        m0047(.A(mai_mai_n75_), .B(mai_mai_n74_), .Y(mai_mai_n76_));
  AN4        m0048(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n77_));
  NAi32      m0049(.An(m), .Bn(k), .C(j), .Y(mai_mai_n78_));
  NOi32      m0050(.An(h), .Bn(g), .C(f), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n73_), .B(mai_mai_n64_), .Y(mai_mai_n80_));
  INV        m0052(.A(n), .Y(mai_mai_n81_));
  NOi32      m0053(.An(e), .Bn(b), .C(d), .Y(mai_mai_n82_));
  NA2        m0054(.A(mai_mai_n82_), .B(mai_mai_n81_), .Y(mai_mai_n83_));
  INV        m0055(.A(j), .Y(mai_mai_n84_));
  AN3        m0056(.A(m), .B(k), .C(i), .Y(mai_mai_n85_));
  NA3        m0057(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(g), .Y(mai_mai_n86_));
  NAi32      m0058(.An(g), .Bn(f), .C(h), .Y(mai_mai_n87_));
  NAi31      m0059(.An(j), .B(m), .C(l), .Y(mai_mai_n88_));
  NA2        m0060(.A(m), .B(l), .Y(mai_mai_n89_));
  NAi31      m0061(.An(k), .B(j), .C(g), .Y(mai_mai_n90_));
  AN2        m0062(.A(j), .B(g), .Y(mai_mai_n91_));
  NOi32      m0063(.An(m), .Bn(l), .C(i), .Y(mai_mai_n92_));
  NOi21      m0064(.An(g), .B(i), .Y(mai_mai_n93_));
  NOi32      m0065(.An(m), .Bn(j), .C(k), .Y(mai_mai_n94_));
  NAi41      m0066(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n95_));
  AN2        m0067(.A(e), .B(b), .Y(mai_mai_n96_));
  NOi31      m0068(.An(c), .B(h), .C(f), .Y(mai_mai_n97_));
  NA2        m0069(.A(mai_mai_n97_), .B(mai_mai_n96_), .Y(mai_mai_n98_));
  NO2        m0070(.A(mai_mai_n98_), .B(mai_mai_n95_), .Y(mai_mai_n99_));
  NOi21      m0071(.An(g), .B(f), .Y(mai_mai_n100_));
  NOi21      m0072(.An(i), .B(h), .Y(mai_mai_n101_));
  NA3        m0073(.A(mai_mai_n101_), .B(mai_mai_n100_), .C(mai_mai_n36_), .Y(mai_mai_n102_));
  INV        m0074(.A(a), .Y(mai_mai_n103_));
  NA2        m0075(.A(mai_mai_n96_), .B(mai_mai_n103_), .Y(mai_mai_n104_));
  INV        m0076(.A(l), .Y(mai_mai_n105_));
  NOi21      m0077(.An(m), .B(n), .Y(mai_mai_n106_));
  AN2        m0078(.A(k), .B(h), .Y(mai_mai_n107_));
  NO2        m0079(.A(mai_mai_n102_), .B(mai_mai_n83_), .Y(mai_mai_n108_));
  INV        m0080(.A(b), .Y(mai_mai_n109_));
  NA2        m0081(.A(l), .B(j), .Y(mai_mai_n110_));
  AN2        m0082(.A(k), .B(i), .Y(mai_mai_n111_));
  NA2        m0083(.A(mai_mai_n111_), .B(mai_mai_n110_), .Y(mai_mai_n112_));
  NA2        m0084(.A(g), .B(e), .Y(mai_mai_n113_));
  NOi32      m0085(.An(c), .Bn(a), .C(d), .Y(mai_mai_n114_));
  NA2        m0086(.A(mai_mai_n114_), .B(mai_mai_n106_), .Y(mai_mai_n115_));
  NO4        m0087(.A(mai_mai_n115_), .B(mai_mai_n113_), .C(mai_mai_n112_), .D(mai_mai_n109_), .Y(mai_mai_n116_));
  NO3        m0088(.A(mai_mai_n116_), .B(mai_mai_n108_), .C(mai_mai_n99_), .Y(mai_mai_n117_));
  INV        m0089(.A(mai_mai_n117_), .Y(mai_mai_n118_));
  NOi31      m0090(.An(k), .B(m), .C(j), .Y(mai_mai_n119_));
  NOi31      m0091(.An(k), .B(m), .C(i), .Y(mai_mai_n120_));
  NOi32      m0092(.An(f), .Bn(b), .C(e), .Y(mai_mai_n121_));
  NAi21      m0093(.An(g), .B(h), .Y(mai_mai_n122_));
  NAi21      m0094(.An(m), .B(n), .Y(mai_mai_n123_));
  NAi21      m0095(.An(j), .B(k), .Y(mai_mai_n124_));
  NO3        m0096(.A(mai_mai_n124_), .B(mai_mai_n123_), .C(mai_mai_n122_), .Y(mai_mai_n125_));
  NAi31      m0097(.An(j), .B(k), .C(h), .Y(mai_mai_n126_));
  NA2        m0098(.A(mai_mai_n125_), .B(mai_mai_n121_), .Y(mai_mai_n127_));
  NO2        m0099(.A(k), .B(j), .Y(mai_mai_n128_));
  AN2        m0100(.A(k), .B(j), .Y(mai_mai_n129_));
  NAi21      m0101(.An(c), .B(b), .Y(mai_mai_n130_));
  NA2        m0102(.A(f), .B(d), .Y(mai_mai_n131_));
  NAi31      m0103(.An(f), .B(e), .C(b), .Y(mai_mai_n132_));
  NA2        m0104(.A(d), .B(b), .Y(mai_mai_n133_));
  NAi21      m0105(.An(e), .B(f), .Y(mai_mai_n134_));
  NO2        m0106(.A(mai_mai_n134_), .B(mai_mai_n133_), .Y(mai_mai_n135_));
  NA2        m0107(.A(b), .B(a), .Y(mai_mai_n136_));
  NAi21      m0108(.An(e), .B(g), .Y(mai_mai_n137_));
  NAi21      m0109(.An(c), .B(d), .Y(mai_mai_n138_));
  NAi31      m0110(.An(l), .B(k), .C(h), .Y(mai_mai_n139_));
  NO2        m0111(.A(mai_mai_n123_), .B(mai_mai_n139_), .Y(mai_mai_n140_));
  INV        m0112(.A(mai_mai_n127_), .Y(mai_mai_n141_));
  NAi31      m0113(.An(e), .B(f), .C(b), .Y(mai_mai_n142_));
  NOi21      m0114(.An(g), .B(d), .Y(mai_mai_n143_));
  NO2        m0115(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n144_));
  NOi21      m0116(.An(h), .B(i), .Y(mai_mai_n145_));
  NOi21      m0117(.An(k), .B(m), .Y(mai_mai_n146_));
  NA3        m0118(.A(mai_mai_n146_), .B(mai_mai_n145_), .C(n), .Y(mai_mai_n147_));
  NOi21      m0119(.An(mai_mai_n144_), .B(mai_mai_n147_), .Y(mai_mai_n148_));
  NOi21      m0120(.An(h), .B(g), .Y(mai_mai_n149_));
  NO2        m0121(.A(mai_mai_n131_), .B(mai_mai_n130_), .Y(mai_mai_n150_));
  NA2        m0122(.A(mai_mai_n150_), .B(mai_mai_n149_), .Y(mai_mai_n151_));
  NAi31      m0123(.An(l), .B(j), .C(h), .Y(mai_mai_n152_));
  NOi32      m0124(.An(n), .Bn(k), .C(m), .Y(mai_mai_n153_));
  NA2        m0125(.A(l), .B(i), .Y(mai_mai_n154_));
  NA2        m0126(.A(mai_mai_n154_), .B(mai_mai_n153_), .Y(mai_mai_n155_));
  NO2        m0127(.A(mai_mai_n155_), .B(mai_mai_n151_), .Y(mai_mai_n156_));
  NAi31      m0128(.An(d), .B(f), .C(c), .Y(mai_mai_n157_));
  NAi31      m0129(.An(e), .B(f), .C(c), .Y(mai_mai_n158_));
  NA2        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NA2        m0131(.A(j), .B(h), .Y(mai_mai_n160_));
  OR3        m0132(.A(n), .B(m), .C(k), .Y(mai_mai_n161_));
  NO2        m0133(.A(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  NAi32      m0134(.An(m), .Bn(k), .C(n), .Y(mai_mai_n163_));
  NO2        m0135(.A(mai_mai_n163_), .B(mai_mai_n160_), .Y(mai_mai_n164_));
  AOI220     m0136(.A0(mai_mai_n164_), .A1(mai_mai_n144_), .B0(mai_mai_n162_), .B1(mai_mai_n159_), .Y(mai_mai_n165_));
  NO2        m0137(.A(n), .B(m), .Y(mai_mai_n166_));
  NA2        m0138(.A(mai_mai_n166_), .B(mai_mai_n50_), .Y(mai_mai_n167_));
  NAi21      m0139(.An(f), .B(e), .Y(mai_mai_n168_));
  NA2        m0140(.A(d), .B(c), .Y(mai_mai_n169_));
  NO2        m0141(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  NOi21      m0142(.An(mai_mai_n170_), .B(mai_mai_n167_), .Y(mai_mai_n171_));
  NAi21      m0143(.An(d), .B(c), .Y(mai_mai_n172_));
  NAi31      m0144(.An(m), .B(n), .C(b), .Y(mai_mai_n173_));
  NA2        m0145(.A(k), .B(i), .Y(mai_mai_n174_));
  NAi21      m0146(.An(h), .B(f), .Y(mai_mai_n175_));
  NO2        m0147(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  NO2        m0148(.A(mai_mai_n173_), .B(mai_mai_n138_), .Y(mai_mai_n177_));
  NA2        m0149(.A(mai_mai_n177_), .B(mai_mai_n176_), .Y(mai_mai_n178_));
  NOi32      m0150(.An(f), .Bn(c), .C(d), .Y(mai_mai_n179_));
  NOi32      m0151(.An(f), .Bn(c), .C(e), .Y(mai_mai_n180_));
  NO2        m0152(.A(mai_mai_n180_), .B(mai_mai_n179_), .Y(mai_mai_n181_));
  NO3        m0153(.A(n), .B(m), .C(j), .Y(mai_mai_n182_));
  NA2        m0154(.A(mai_mai_n182_), .B(mai_mai_n107_), .Y(mai_mai_n183_));
  AO210      m0155(.A0(mai_mai_n183_), .A1(mai_mai_n167_), .B0(mai_mai_n181_), .Y(mai_mai_n184_));
  NAi41      m0156(.An(mai_mai_n171_), .B(mai_mai_n184_), .C(mai_mai_n178_), .D(mai_mai_n165_), .Y(mai_mai_n185_));
  OR4        m0157(.A(mai_mai_n185_), .B(mai_mai_n156_), .C(mai_mai_n148_), .D(mai_mai_n141_), .Y(mai_mai_n186_));
  NO4        m0158(.A(mai_mai_n186_), .B(mai_mai_n118_), .C(mai_mai_n80_), .D(mai_mai_n55_), .Y(mai_mai_n187_));
  NA3        m0159(.A(m), .B(mai_mai_n105_), .C(j), .Y(mai_mai_n188_));
  NAi31      m0160(.An(n), .B(h), .C(g), .Y(mai_mai_n189_));
  NO2        m0161(.A(mai_mai_n189_), .B(mai_mai_n188_), .Y(mai_mai_n190_));
  NOi32      m0162(.An(m), .Bn(k), .C(l), .Y(mai_mai_n191_));
  NA3        m0163(.A(mai_mai_n191_), .B(mai_mai_n84_), .C(g), .Y(mai_mai_n192_));
  NO2        m0164(.A(mai_mai_n192_), .B(n), .Y(mai_mai_n193_));
  NOi21      m0165(.An(k), .B(j), .Y(mai_mai_n194_));
  NA4        m0166(.A(mai_mai_n194_), .B(mai_mai_n106_), .C(i), .D(g), .Y(mai_mai_n195_));
  AN2        m0167(.A(i), .B(g), .Y(mai_mai_n196_));
  NA3        m0168(.A(mai_mai_n75_), .B(mai_mai_n196_), .C(mai_mai_n106_), .Y(mai_mai_n197_));
  NA2        m0169(.A(mai_mai_n197_), .B(mai_mai_n195_), .Y(mai_mai_n198_));
  NO2        m0170(.A(mai_mai_n198_), .B(mai_mai_n193_), .Y(mai_mai_n199_));
  NAi41      m0171(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n200_));
  INV        m0172(.A(mai_mai_n200_), .Y(mai_mai_n201_));
  INV        m0173(.A(f), .Y(mai_mai_n202_));
  INV        m0174(.A(g), .Y(mai_mai_n203_));
  NOi31      m0175(.An(i), .B(j), .C(h), .Y(mai_mai_n204_));
  NOi21      m0176(.An(l), .B(m), .Y(mai_mai_n205_));
  NA2        m0177(.A(mai_mai_n205_), .B(mai_mai_n204_), .Y(mai_mai_n206_));
  NO2        m0178(.A(mai_mai_n199_), .B(mai_mai_n32_), .Y(mai_mai_n207_));
  NOi21      m0179(.An(n), .B(m), .Y(mai_mai_n208_));
  NOi32      m0180(.An(l), .Bn(i), .C(j), .Y(mai_mai_n209_));
  NA2        m0181(.A(mai_mai_n209_), .B(mai_mai_n208_), .Y(mai_mai_n210_));
  OR2        m0182(.A(mai_mai_n210_), .B(mai_mai_n98_), .Y(mai_mai_n211_));
  NAi21      m0183(.An(j), .B(h), .Y(mai_mai_n212_));
  XN2        m0184(.A(i), .B(h), .Y(mai_mai_n213_));
  NA2        m0185(.A(mai_mai_n213_), .B(mai_mai_n212_), .Y(mai_mai_n214_));
  NOi31      m0186(.An(k), .B(n), .C(m), .Y(mai_mai_n215_));
  NOi31      m0187(.An(mai_mai_n215_), .B(mai_mai_n169_), .C(mai_mai_n168_), .Y(mai_mai_n216_));
  NA2        m0188(.A(mai_mai_n216_), .B(mai_mai_n214_), .Y(mai_mai_n217_));
  NAi31      m0189(.An(f), .B(e), .C(c), .Y(mai_mai_n218_));
  NO4        m0190(.A(mai_mai_n218_), .B(mai_mai_n161_), .C(mai_mai_n160_), .D(mai_mai_n59_), .Y(mai_mai_n219_));
  NA4        m0191(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n220_));
  NAi32      m0192(.An(m), .Bn(i), .C(k), .Y(mai_mai_n221_));
  NO3        m0193(.A(mai_mai_n221_), .B(mai_mai_n87_), .C(mai_mai_n220_), .Y(mai_mai_n222_));
  INV        m0194(.A(k), .Y(mai_mai_n223_));
  NO2        m0195(.A(mai_mai_n222_), .B(mai_mai_n219_), .Y(mai_mai_n224_));
  NAi21      m0196(.An(n), .B(a), .Y(mai_mai_n225_));
  NO2        m0197(.A(mai_mai_n225_), .B(mai_mai_n133_), .Y(mai_mai_n226_));
  NAi41      m0198(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n227_));
  NO2        m0199(.A(mai_mai_n227_), .B(e), .Y(mai_mai_n228_));
  NO3        m0200(.A(mai_mai_n134_), .B(mai_mai_n90_), .C(mai_mai_n89_), .Y(mai_mai_n229_));
  OAI210     m0201(.A0(mai_mai_n229_), .A1(mai_mai_n228_), .B0(mai_mai_n226_), .Y(mai_mai_n230_));
  AN4        m0202(.A(mai_mai_n230_), .B(mai_mai_n224_), .C(mai_mai_n217_), .D(mai_mai_n211_), .Y(mai_mai_n231_));
  OR2        m0203(.A(h), .B(g), .Y(mai_mai_n232_));
  NO2        m0204(.A(mai_mai_n232_), .B(mai_mai_n95_), .Y(mai_mai_n233_));
  NA2        m0205(.A(mai_mai_n233_), .B(mai_mai_n121_), .Y(mai_mai_n234_));
  NA2        m0206(.A(mai_mai_n146_), .B(mai_mai_n101_), .Y(mai_mai_n235_));
  NO2        m0207(.A(n), .B(a), .Y(mai_mai_n236_));
  NAi31      m0208(.An(mai_mai_n227_), .B(mai_mai_n236_), .C(mai_mai_n96_), .Y(mai_mai_n237_));
  NAi21      m0209(.An(h), .B(i), .Y(mai_mai_n238_));
  NA2        m0210(.A(mai_mai_n166_), .B(k), .Y(mai_mai_n239_));
  NO2        m0211(.A(mai_mai_n239_), .B(mai_mai_n238_), .Y(mai_mai_n240_));
  NA2        m0212(.A(mai_mai_n240_), .B(mai_mai_n179_), .Y(mai_mai_n241_));
  NA3        m0213(.A(mai_mai_n241_), .B(mai_mai_n237_), .C(mai_mai_n234_), .Y(mai_mai_n242_));
  NOi21      m0214(.An(g), .B(e), .Y(mai_mai_n243_));
  NO2        m0215(.A(mai_mai_n72_), .B(mai_mai_n74_), .Y(mai_mai_n244_));
  NA2        m0216(.A(mai_mai_n244_), .B(mai_mai_n243_), .Y(mai_mai_n245_));
  NOi32      m0217(.An(l), .Bn(j), .C(i), .Y(mai_mai_n246_));
  AOI210     m0218(.A0(mai_mai_n75_), .A1(mai_mai_n84_), .B0(mai_mai_n246_), .Y(mai_mai_n247_));
  NAi21      m0219(.An(f), .B(g), .Y(mai_mai_n248_));
  NO2        m0220(.A(mai_mai_n248_), .B(mai_mai_n65_), .Y(mai_mai_n249_));
  NO2        m0221(.A(mai_mai_n69_), .B(mai_mai_n110_), .Y(mai_mai_n250_));
  NO2        m0222(.A(mai_mai_n247_), .B(mai_mai_n245_), .Y(mai_mai_n251_));
  NO3        m0223(.A(mai_mai_n124_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n252_));
  NOi41      m0224(.An(mai_mai_n231_), .B(mai_mai_n251_), .C(mai_mai_n242_), .D(mai_mai_n207_), .Y(mai_mai_n253_));
  NO4        m0225(.A(mai_mai_n190_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n254_));
  NO2        m0226(.A(mai_mai_n254_), .B(mai_mai_n104_), .Y(mai_mai_n255_));
  NA3        m0227(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n256_));
  NAi21      m0228(.An(h), .B(g), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n235_), .B(mai_mai_n248_), .Y(mai_mai_n258_));
  NAi31      m0230(.An(g), .B(k), .C(h), .Y(mai_mai_n259_));
  NO3        m0231(.A(mai_mai_n123_), .B(mai_mai_n259_), .C(l), .Y(mai_mai_n260_));
  NAi31      m0232(.An(e), .B(d), .C(a), .Y(mai_mai_n261_));
  NA2        m0233(.A(mai_mai_n260_), .B(mai_mai_n121_), .Y(mai_mai_n262_));
  INV        m0234(.A(mai_mai_n262_), .Y(mai_mai_n263_));
  NA4        m0235(.A(mai_mai_n146_), .B(mai_mai_n79_), .C(mai_mai_n77_), .D(mai_mai_n110_), .Y(mai_mai_n264_));
  NA3        m0236(.A(mai_mai_n146_), .B(mai_mai_n145_), .C(mai_mai_n81_), .Y(mai_mai_n265_));
  NO2        m0237(.A(mai_mai_n265_), .B(mai_mai_n181_), .Y(mai_mai_n266_));
  NOi21      m0238(.An(mai_mai_n264_), .B(mai_mai_n266_), .Y(mai_mai_n267_));
  NA3        m0239(.A(e), .B(c), .C(b), .Y(mai_mai_n268_));
  NO2        m0240(.A(mai_mai_n60_), .B(mai_mai_n268_), .Y(mai_mai_n269_));
  NAi32      m0241(.An(k), .Bn(i), .C(j), .Y(mai_mai_n270_));
  NAi31      m0242(.An(h), .B(l), .C(i), .Y(mai_mai_n271_));
  NA3        m0243(.A(mai_mai_n271_), .B(mai_mai_n270_), .C(mai_mai_n152_), .Y(mai_mai_n272_));
  NOi21      m0244(.An(mai_mai_n272_), .B(mai_mai_n49_), .Y(mai_mai_n273_));
  OAI210     m0245(.A0(mai_mai_n249_), .A1(mai_mai_n269_), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  NAi21      m0246(.An(l), .B(k), .Y(mai_mai_n275_));
  NO2        m0247(.A(mai_mai_n275_), .B(mai_mai_n49_), .Y(mai_mai_n276_));
  NOi21      m0248(.An(l), .B(j), .Y(mai_mai_n277_));
  NA2        m0249(.A(mai_mai_n149_), .B(mai_mai_n277_), .Y(mai_mai_n278_));
  NA3        m0250(.A(mai_mai_n111_), .B(mai_mai_n110_), .C(g), .Y(mai_mai_n279_));
  OR3        m0251(.A(mai_mai_n72_), .B(mai_mai_n74_), .C(e), .Y(mai_mai_n280_));
  AOI210     m0252(.A0(mai_mai_n279_), .A1(mai_mai_n278_), .B0(mai_mai_n280_), .Y(mai_mai_n281_));
  INV        m0253(.A(mai_mai_n281_), .Y(mai_mai_n282_));
  NAi32      m0254(.An(j), .Bn(h), .C(i), .Y(mai_mai_n283_));
  NAi21      m0255(.An(m), .B(l), .Y(mai_mai_n284_));
  NO3        m0256(.A(mai_mai_n284_), .B(mai_mai_n283_), .C(mai_mai_n81_), .Y(mai_mai_n285_));
  NA2        m0257(.A(h), .B(g), .Y(mai_mai_n286_));
  NA2        m0258(.A(mai_mai_n285_), .B(mai_mai_n150_), .Y(mai_mai_n287_));
  NA4        m0259(.A(mai_mai_n287_), .B(mai_mai_n282_), .C(mai_mai_n274_), .D(mai_mai_n267_), .Y(mai_mai_n288_));
  NO2        m0260(.A(mai_mai_n132_), .B(d), .Y(mai_mai_n289_));
  NA2        m0261(.A(mai_mai_n289_), .B(mai_mai_n53_), .Y(mai_mai_n290_));
  NO2        m0262(.A(mai_mai_n98_), .B(mai_mai_n95_), .Y(mai_mai_n291_));
  NAi32      m0263(.An(n), .Bn(m), .C(l), .Y(mai_mai_n292_));
  NO2        m0264(.A(mai_mai_n292_), .B(mai_mai_n283_), .Y(mai_mai_n293_));
  NA2        m0265(.A(mai_mai_n293_), .B(mai_mai_n170_), .Y(mai_mai_n294_));
  NO2        m0266(.A(mai_mai_n115_), .B(mai_mai_n109_), .Y(mai_mai_n295_));
  NAi31      m0267(.An(k), .B(l), .C(j), .Y(mai_mai_n296_));
  OAI210     m0268(.A0(mai_mai_n275_), .A1(j), .B0(mai_mai_n296_), .Y(mai_mai_n297_));
  NOi21      m0269(.An(mai_mai_n297_), .B(mai_mai_n113_), .Y(mai_mai_n298_));
  NA2        m0270(.A(mai_mai_n298_), .B(mai_mai_n295_), .Y(mai_mai_n299_));
  NA3        m0271(.A(mai_mai_n299_), .B(mai_mai_n294_), .C(mai_mai_n290_), .Y(mai_mai_n300_));
  NO4        m0272(.A(mai_mai_n300_), .B(mai_mai_n288_), .C(mai_mai_n263_), .D(mai_mai_n255_), .Y(mai_mai_n301_));
  NA2        m0273(.A(mai_mai_n240_), .B(mai_mai_n180_), .Y(mai_mai_n302_));
  NAi21      m0274(.An(m), .B(k), .Y(mai_mai_n303_));
  NO2        m0275(.A(mai_mai_n213_), .B(mai_mai_n303_), .Y(mai_mai_n304_));
  NAi41      m0276(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n305_), .B(mai_mai_n137_), .Y(mai_mai_n306_));
  NA2        m0278(.A(mai_mai_n306_), .B(mai_mai_n304_), .Y(mai_mai_n307_));
  NAi31      m0279(.An(i), .B(l), .C(h), .Y(mai_mai_n308_));
  NA2        m0280(.A(e), .B(c), .Y(mai_mai_n309_));
  NO3        m0281(.A(mai_mai_n309_), .B(n), .C(d), .Y(mai_mai_n310_));
  NOi21      m0282(.An(f), .B(h), .Y(mai_mai_n311_));
  NA2        m0283(.A(mai_mai_n311_), .B(mai_mai_n111_), .Y(mai_mai_n312_));
  NO2        m0284(.A(mai_mai_n312_), .B(mai_mai_n203_), .Y(mai_mai_n313_));
  NAi31      m0285(.An(d), .B(e), .C(b), .Y(mai_mai_n314_));
  NO2        m0286(.A(mai_mai_n123_), .B(mai_mai_n314_), .Y(mai_mai_n315_));
  NA2        m0287(.A(mai_mai_n315_), .B(mai_mai_n313_), .Y(mai_mai_n316_));
  NA3        m0288(.A(mai_mai_n316_), .B(mai_mai_n307_), .C(mai_mai_n302_), .Y(mai_mai_n317_));
  NA2        m0289(.A(mai_mai_n236_), .B(mai_mai_n96_), .Y(mai_mai_n318_));
  OR2        m0290(.A(mai_mai_n318_), .B(mai_mai_n192_), .Y(mai_mai_n319_));
  NOi31      m0291(.An(l), .B(n), .C(m), .Y(mai_mai_n320_));
  NA2        m0292(.A(mai_mai_n320_), .B(mai_mai_n204_), .Y(mai_mai_n321_));
  NO2        m0293(.A(mai_mai_n321_), .B(mai_mai_n181_), .Y(mai_mai_n322_));
  NAi21      m0294(.An(mai_mai_n322_), .B(mai_mai_n319_), .Y(mai_mai_n323_));
  NAi32      m0295(.An(m), .Bn(j), .C(k), .Y(mai_mai_n324_));
  NAi41      m0296(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n325_));
  OAI210     m0297(.A0(mai_mai_n200_), .A1(mai_mai_n324_), .B0(mai_mai_n325_), .Y(mai_mai_n326_));
  NOi31      m0298(.An(j), .B(m), .C(k), .Y(mai_mai_n327_));
  NO2        m0299(.A(mai_mai_n119_), .B(mai_mai_n327_), .Y(mai_mai_n328_));
  AN3        m0300(.A(h), .B(g), .C(f), .Y(mai_mai_n329_));
  NAi31      m0301(.An(mai_mai_n328_), .B(mai_mai_n329_), .C(mai_mai_n326_), .Y(mai_mai_n330_));
  NOi32      m0302(.An(m), .Bn(j), .C(l), .Y(mai_mai_n331_));
  NO2        m0303(.A(mai_mai_n331_), .B(mai_mai_n92_), .Y(mai_mai_n332_));
  NO2        m0304(.A(mai_mai_n284_), .B(mai_mai_n283_), .Y(mai_mai_n333_));
  NO2        m0305(.A(mai_mai_n206_), .B(g), .Y(mai_mai_n334_));
  NO2        m0306(.A(mai_mai_n142_), .B(mai_mai_n81_), .Y(mai_mai_n335_));
  INV        m0307(.A(mai_mai_n78_), .Y(mai_mai_n336_));
  NA3        m0308(.A(mai_mai_n336_), .B(mai_mai_n329_), .C(mai_mai_n201_), .Y(mai_mai_n337_));
  NA2        m0309(.A(mai_mai_n337_), .B(mai_mai_n330_), .Y(mai_mai_n338_));
  NA3        m0310(.A(h), .B(g), .C(f), .Y(mai_mai_n339_));
  NO2        m0311(.A(mai_mai_n339_), .B(mai_mai_n76_), .Y(mai_mai_n340_));
  NA2        m0312(.A(mai_mai_n325_), .B(mai_mai_n200_), .Y(mai_mai_n341_));
  NA2        m0313(.A(mai_mai_n149_), .B(e), .Y(mai_mai_n342_));
  NO2        m0314(.A(mai_mai_n342_), .B(mai_mai_n41_), .Y(mai_mai_n343_));
  AOI220     m0315(.A0(mai_mai_n343_), .A1(mai_mai_n295_), .B0(mai_mai_n341_), .B1(mai_mai_n340_), .Y(mai_mai_n344_));
  NOi32      m0316(.An(j), .Bn(g), .C(i), .Y(mai_mai_n345_));
  NA3        m0317(.A(mai_mai_n345_), .B(mai_mai_n275_), .C(mai_mai_n106_), .Y(mai_mai_n346_));
  AO210      m0318(.A0(mai_mai_n104_), .A1(mai_mai_n32_), .B0(mai_mai_n346_), .Y(mai_mai_n347_));
  NOi32      m0319(.An(e), .Bn(b), .C(a), .Y(mai_mai_n348_));
  AN2        m0320(.A(l), .B(j), .Y(mai_mai_n349_));
  NA3        m0321(.A(mai_mai_n197_), .B(mai_mai_n195_), .C(mai_mai_n35_), .Y(mai_mai_n350_));
  NA2        m0322(.A(mai_mai_n350_), .B(mai_mai_n348_), .Y(mai_mai_n351_));
  NO2        m0323(.A(mai_mai_n314_), .B(n), .Y(mai_mai_n352_));
  NA2        m0324(.A(mai_mai_n196_), .B(k), .Y(mai_mai_n353_));
  NA3        m0325(.A(m), .B(mai_mai_n105_), .C(mai_mai_n202_), .Y(mai_mai_n354_));
  NA4        m0326(.A(mai_mai_n191_), .B(mai_mai_n84_), .C(g), .D(mai_mai_n202_), .Y(mai_mai_n355_));
  INV        m0327(.A(mai_mai_n355_), .Y(mai_mai_n356_));
  NAi41      m0328(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n51_), .B(mai_mai_n106_), .Y(mai_mai_n358_));
  NA2        m0330(.A(mai_mai_n356_), .B(mai_mai_n352_), .Y(mai_mai_n359_));
  NA4        m0331(.A(mai_mai_n359_), .B(mai_mai_n351_), .C(mai_mai_n347_), .D(mai_mai_n344_), .Y(mai_mai_n360_));
  NO4        m0332(.A(mai_mai_n360_), .B(mai_mai_n338_), .C(mai_mai_n323_), .D(mai_mai_n317_), .Y(mai_mai_n361_));
  NA4        m0333(.A(mai_mai_n361_), .B(mai_mai_n301_), .C(mai_mai_n253_), .D(mai_mai_n187_), .Y(mai10));
  NA3        m0334(.A(m), .B(k), .C(i), .Y(mai_mai_n363_));
  NO3        m0335(.A(mai_mai_n363_), .B(j), .C(mai_mai_n203_), .Y(mai_mai_n364_));
  NOi21      m0336(.An(e), .B(f), .Y(mai_mai_n365_));
  NO4        m0337(.A(mai_mai_n138_), .B(mai_mai_n365_), .C(n), .D(mai_mai_n103_), .Y(mai_mai_n366_));
  NAi31      m0338(.An(b), .B(f), .C(c), .Y(mai_mai_n367_));
  INV        m0339(.A(mai_mai_n367_), .Y(mai_mai_n368_));
  NOi32      m0340(.An(k), .Bn(h), .C(j), .Y(mai_mai_n369_));
  NA2        m0341(.A(mai_mai_n369_), .B(mai_mai_n208_), .Y(mai_mai_n370_));
  NA2        m0342(.A(mai_mai_n147_), .B(mai_mai_n370_), .Y(mai_mai_n371_));
  AOI220     m0343(.A0(mai_mai_n371_), .A1(mai_mai_n368_), .B0(mai_mai_n366_), .B1(mai_mai_n364_), .Y(mai_mai_n372_));
  AN2        m0344(.A(j), .B(h), .Y(mai_mai_n373_));
  NO3        m0345(.A(n), .B(m), .C(k), .Y(mai_mai_n374_));
  NA2        m0346(.A(mai_mai_n374_), .B(mai_mai_n373_), .Y(mai_mai_n375_));
  NO3        m0347(.A(mai_mai_n375_), .B(mai_mai_n138_), .C(mai_mai_n202_), .Y(mai_mai_n376_));
  OR2        m0348(.A(m), .B(k), .Y(mai_mai_n377_));
  NO2        m0349(.A(mai_mai_n160_), .B(mai_mai_n377_), .Y(mai_mai_n378_));
  NA4        m0350(.A(n), .B(f), .C(c), .D(mai_mai_n109_), .Y(mai_mai_n379_));
  NOi21      m0351(.An(mai_mai_n378_), .B(mai_mai_n379_), .Y(mai_mai_n380_));
  NOi32      m0352(.An(d), .Bn(a), .C(c), .Y(mai_mai_n381_));
  NA2        m0353(.A(mai_mai_n381_), .B(mai_mai_n168_), .Y(mai_mai_n382_));
  NAi21      m0354(.An(i), .B(g), .Y(mai_mai_n383_));
  NAi31      m0355(.An(k), .B(m), .C(j), .Y(mai_mai_n384_));
  NO3        m0356(.A(mai_mai_n384_), .B(mai_mai_n383_), .C(n), .Y(mai_mai_n385_));
  NOi21      m0357(.An(mai_mai_n385_), .B(mai_mai_n382_), .Y(mai_mai_n386_));
  NO3        m0358(.A(mai_mai_n386_), .B(mai_mai_n380_), .C(mai_mai_n376_), .Y(mai_mai_n387_));
  NO2        m0359(.A(mai_mai_n379_), .B(mai_mai_n284_), .Y(mai_mai_n388_));
  NOi32      m0360(.An(f), .Bn(d), .C(c), .Y(mai_mai_n389_));
  AOI220     m0361(.A0(mai_mai_n389_), .A1(mai_mai_n293_), .B0(mai_mai_n388_), .B1(mai_mai_n204_), .Y(mai_mai_n390_));
  NA3        m0362(.A(mai_mai_n390_), .B(mai_mai_n387_), .C(mai_mai_n372_), .Y(mai_mai_n391_));
  NO2        m0363(.A(mai_mai_n59_), .B(mai_mai_n109_), .Y(mai_mai_n392_));
  NA2        m0364(.A(mai_mai_n236_), .B(mai_mai_n392_), .Y(mai_mai_n393_));
  INV        m0365(.A(e), .Y(mai_mai_n394_));
  NA2        m0366(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n395_));
  OAI220     m0367(.A0(mai_mai_n395_), .A1(mai_mai_n188_), .B0(mai_mai_n192_), .B1(mai_mai_n394_), .Y(mai_mai_n396_));
  AN2        m0368(.A(g), .B(e), .Y(mai_mai_n397_));
  NA3        m0369(.A(mai_mai_n397_), .B(mai_mai_n191_), .C(i), .Y(mai_mai_n398_));
  OAI210     m0370(.A0(mai_mai_n86_), .A1(mai_mai_n394_), .B0(mai_mai_n398_), .Y(mai_mai_n399_));
  NO2        m0371(.A(mai_mai_n399_), .B(mai_mai_n396_), .Y(mai_mai_n400_));
  NOi32      m0372(.An(h), .Bn(e), .C(g), .Y(mai_mai_n401_));
  NA3        m0373(.A(mai_mai_n401_), .B(mai_mai_n277_), .C(m), .Y(mai_mai_n402_));
  NOi21      m0374(.An(g), .B(h), .Y(mai_mai_n403_));
  AN3        m0375(.A(m), .B(l), .C(i), .Y(mai_mai_n404_));
  NA3        m0376(.A(mai_mai_n404_), .B(mai_mai_n403_), .C(e), .Y(mai_mai_n405_));
  AN3        m0377(.A(h), .B(g), .C(e), .Y(mai_mai_n406_));
  NA2        m0378(.A(mai_mai_n406_), .B(mai_mai_n92_), .Y(mai_mai_n407_));
  AN2        m0379(.A(mai_mai_n407_), .B(mai_mai_n402_), .Y(mai_mai_n408_));
  AOI210     m0380(.A0(mai_mai_n408_), .A1(mai_mai_n400_), .B0(mai_mai_n393_), .Y(mai_mai_n409_));
  NA3        m0381(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n410_));
  NO2        m0382(.A(mai_mai_n410_), .B(mai_mai_n393_), .Y(mai_mai_n411_));
  NA3        m0383(.A(mai_mai_n381_), .B(mai_mai_n168_), .C(mai_mai_n81_), .Y(mai_mai_n412_));
  NAi31      m0384(.An(b), .B(c), .C(a), .Y(mai_mai_n413_));
  NO2        m0385(.A(mai_mai_n413_), .B(n), .Y(mai_mai_n414_));
  NA2        m0386(.A(mai_mai_n51_), .B(m), .Y(mai_mai_n415_));
  NO2        m0387(.A(mai_mai_n415_), .B(mai_mai_n134_), .Y(mai_mai_n416_));
  NA2        m0388(.A(mai_mai_n416_), .B(mai_mai_n414_), .Y(mai_mai_n417_));
  INV        m0389(.A(mai_mai_n417_), .Y(mai_mai_n418_));
  NO4        m0390(.A(mai_mai_n418_), .B(mai_mai_n411_), .C(mai_mai_n409_), .D(mai_mai_n391_), .Y(mai_mai_n419_));
  NA2        m0391(.A(i), .B(g), .Y(mai_mai_n420_));
  NO3        m0392(.A(mai_mai_n261_), .B(mai_mai_n420_), .C(c), .Y(mai_mai_n421_));
  NOi21      m0393(.An(a), .B(n), .Y(mai_mai_n422_));
  NOi21      m0394(.An(d), .B(c), .Y(mai_mai_n423_));
  NA2        m0395(.A(mai_mai_n423_), .B(mai_mai_n422_), .Y(mai_mai_n424_));
  NA3        m0396(.A(i), .B(g), .C(f), .Y(mai_mai_n425_));
  OR2        m0397(.A(mai_mai_n425_), .B(mai_mai_n71_), .Y(mai_mai_n426_));
  NA3        m0398(.A(mai_mai_n404_), .B(mai_mai_n403_), .C(mai_mai_n168_), .Y(mai_mai_n427_));
  AOI210     m0399(.A0(mai_mai_n427_), .A1(mai_mai_n426_), .B0(mai_mai_n424_), .Y(mai_mai_n428_));
  AOI210     m0400(.A0(mai_mai_n421_), .A1(mai_mai_n276_), .B0(mai_mai_n428_), .Y(mai_mai_n429_));
  OR2        m0401(.A(n), .B(m), .Y(mai_mai_n430_));
  NO2        m0402(.A(mai_mai_n430_), .B(mai_mai_n139_), .Y(mai_mai_n431_));
  NO2        m0403(.A(mai_mai_n169_), .B(mai_mai_n134_), .Y(mai_mai_n432_));
  OAI210     m0404(.A0(mai_mai_n431_), .A1(mai_mai_n162_), .B0(mai_mai_n432_), .Y(mai_mai_n433_));
  INV        m0405(.A(mai_mai_n358_), .Y(mai_mai_n434_));
  NA3        m0406(.A(mai_mai_n434_), .B(mai_mai_n348_), .C(d), .Y(mai_mai_n435_));
  NO2        m0407(.A(mai_mai_n413_), .B(mai_mai_n49_), .Y(mai_mai_n436_));
  NO3        m0408(.A(mai_mai_n66_), .B(mai_mai_n105_), .C(e), .Y(mai_mai_n437_));
  NAi21      m0409(.An(k), .B(j), .Y(mai_mai_n438_));
  NA2        m0410(.A(mai_mai_n238_), .B(mai_mai_n438_), .Y(mai_mai_n439_));
  NA3        m0411(.A(mai_mai_n439_), .B(mai_mai_n437_), .C(mai_mai_n436_), .Y(mai_mai_n440_));
  NAi21      m0412(.An(e), .B(d), .Y(mai_mai_n441_));
  INV        m0413(.A(mai_mai_n441_), .Y(mai_mai_n442_));
  NO2        m0414(.A(mai_mai_n239_), .B(mai_mai_n202_), .Y(mai_mai_n443_));
  NA3        m0415(.A(mai_mai_n443_), .B(mai_mai_n442_), .C(mai_mai_n214_), .Y(mai_mai_n444_));
  NA4        m0416(.A(mai_mai_n444_), .B(mai_mai_n440_), .C(mai_mai_n435_), .D(mai_mai_n433_), .Y(mai_mai_n445_));
  NO2        m0417(.A(mai_mai_n321_), .B(mai_mai_n202_), .Y(mai_mai_n446_));
  NA2        m0418(.A(mai_mai_n446_), .B(mai_mai_n442_), .Y(mai_mai_n447_));
  NOi31      m0419(.An(n), .B(m), .C(k), .Y(mai_mai_n448_));
  AOI220     m0420(.A0(mai_mai_n448_), .A1(mai_mai_n373_), .B0(mai_mai_n208_), .B1(mai_mai_n50_), .Y(mai_mai_n449_));
  NAi31      m0421(.An(g), .B(f), .C(c), .Y(mai_mai_n450_));
  OR3        m0422(.A(mai_mai_n450_), .B(mai_mai_n449_), .C(e), .Y(mai_mai_n451_));
  NA3        m0423(.A(mai_mai_n451_), .B(mai_mai_n447_), .C(mai_mai_n294_), .Y(mai_mai_n452_));
  NOi41      m0424(.An(mai_mai_n429_), .B(mai_mai_n452_), .C(mai_mai_n445_), .D(mai_mai_n251_), .Y(mai_mai_n453_));
  NOi32      m0425(.An(c), .Bn(a), .C(b), .Y(mai_mai_n454_));
  NA2        m0426(.A(mai_mai_n454_), .B(mai_mai_n106_), .Y(mai_mai_n455_));
  INV        m0427(.A(mai_mai_n259_), .Y(mai_mai_n456_));
  AN2        m0428(.A(e), .B(d), .Y(mai_mai_n457_));
  NA2        m0429(.A(mai_mai_n457_), .B(mai_mai_n456_), .Y(mai_mai_n458_));
  INV        m0430(.A(mai_mai_n134_), .Y(mai_mai_n459_));
  NO2        m0431(.A(mai_mai_n122_), .B(mai_mai_n41_), .Y(mai_mai_n460_));
  NO2        m0432(.A(mai_mai_n66_), .B(e), .Y(mai_mai_n461_));
  NOi31      m0433(.An(j), .B(k), .C(i), .Y(mai_mai_n462_));
  NOi21      m0434(.An(mai_mai_n152_), .B(mai_mai_n462_), .Y(mai_mai_n463_));
  NA4        m0435(.A(mai_mai_n308_), .B(mai_mai_n463_), .C(mai_mai_n247_), .D(mai_mai_n112_), .Y(mai_mai_n464_));
  NA2        m0436(.A(mai_mai_n464_), .B(mai_mai_n461_), .Y(mai_mai_n465_));
  AOI210     m0437(.A0(mai_mai_n465_), .A1(mai_mai_n458_), .B0(mai_mai_n455_), .Y(mai_mai_n466_));
  NO2        m0438(.A(mai_mai_n198_), .B(mai_mai_n193_), .Y(mai_mai_n467_));
  NOi21      m0439(.An(a), .B(b), .Y(mai_mai_n468_));
  NA3        m0440(.A(e), .B(d), .C(c), .Y(mai_mai_n469_));
  NAi21      m0441(.An(mai_mai_n469_), .B(mai_mai_n468_), .Y(mai_mai_n470_));
  NO2        m0442(.A(mai_mai_n412_), .B(mai_mai_n192_), .Y(mai_mai_n471_));
  NOi21      m0443(.An(mai_mai_n470_), .B(mai_mai_n471_), .Y(mai_mai_n472_));
  AOI210     m0444(.A0(mai_mai_n254_), .A1(mai_mai_n467_), .B0(mai_mai_n472_), .Y(mai_mai_n473_));
  NO4        m0445(.A(mai_mai_n175_), .B(mai_mai_n95_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n474_));
  NA2        m0446(.A(mai_mai_n368_), .B(mai_mai_n140_), .Y(mai_mai_n475_));
  OR2        m0447(.A(k), .B(j), .Y(mai_mai_n476_));
  NA2        m0448(.A(l), .B(k), .Y(mai_mai_n477_));
  AOI210     m0449(.A0(mai_mai_n221_), .A1(mai_mai_n324_), .B0(mai_mai_n81_), .Y(mai_mai_n478_));
  INV        m0450(.A(mai_mai_n264_), .Y(mai_mai_n479_));
  NA2        m0451(.A(mai_mai_n381_), .B(mai_mai_n106_), .Y(mai_mai_n480_));
  NO4        m0452(.A(mai_mai_n480_), .B(mai_mai_n90_), .C(mai_mai_n105_), .D(e), .Y(mai_mai_n481_));
  NO3        m0453(.A(mai_mai_n412_), .B(mai_mai_n88_), .C(mai_mai_n122_), .Y(mai_mai_n482_));
  NO3        m0454(.A(mai_mai_n482_), .B(mai_mai_n481_), .C(mai_mai_n479_), .Y(mai_mai_n483_));
  NA2        m0455(.A(mai_mai_n483_), .B(mai_mai_n475_), .Y(mai_mai_n484_));
  NO4        m0456(.A(mai_mai_n484_), .B(mai_mai_n474_), .C(mai_mai_n473_), .D(mai_mai_n466_), .Y(mai_mai_n485_));
  NA2        m0457(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n486_));
  NOi21      m0458(.An(d), .B(e), .Y(mai_mai_n487_));
  NAi31      m0459(.An(j), .B(l), .C(i), .Y(mai_mai_n488_));
  OAI210     m0460(.A0(mai_mai_n488_), .A1(mai_mai_n123_), .B0(mai_mai_n95_), .Y(mai_mai_n489_));
  NO3        m0461(.A(mai_mai_n382_), .B(mai_mai_n332_), .C(mai_mai_n189_), .Y(mai_mai_n490_));
  NO2        m0462(.A(mai_mai_n382_), .B(mai_mai_n358_), .Y(mai_mai_n491_));
  NO4        m0463(.A(mai_mai_n491_), .B(mai_mai_n490_), .C(mai_mai_n171_), .D(mai_mai_n291_), .Y(mai_mai_n492_));
  NA3        m0464(.A(mai_mai_n492_), .B(mai_mai_n486_), .C(mai_mai_n231_), .Y(mai_mai_n493_));
  OAI210     m0465(.A0(mai_mai_n120_), .A1(mai_mai_n119_), .B0(n), .Y(mai_mai_n494_));
  NO2        m0466(.A(mai_mai_n494_), .B(mai_mai_n122_), .Y(mai_mai_n495_));
  OA210      m0467(.A0(mai_mai_n233_), .A1(mai_mai_n495_), .B0(mai_mai_n180_), .Y(mai_mai_n496_));
  XO2        m0468(.A(i), .B(h), .Y(mai_mai_n497_));
  NA3        m0469(.A(mai_mai_n497_), .B(mai_mai_n146_), .C(n), .Y(mai_mai_n498_));
  NAi41      m0470(.An(mai_mai_n285_), .B(mai_mai_n498_), .C(mai_mai_n449_), .D(mai_mai_n370_), .Y(mai_mai_n499_));
  NOi32      m0471(.An(mai_mai_n499_), .Bn(mai_mai_n461_), .C(mai_mai_n256_), .Y(mai_mai_n500_));
  NAi31      m0472(.An(c), .B(f), .C(d), .Y(mai_mai_n501_));
  AOI210     m0473(.A0(mai_mai_n265_), .A1(mai_mai_n183_), .B0(mai_mai_n501_), .Y(mai_mai_n502_));
  INV        m0474(.A(mai_mai_n502_), .Y(mai_mai_n503_));
  NA3        m0475(.A(mai_mai_n366_), .B(mai_mai_n92_), .C(mai_mai_n91_), .Y(mai_mai_n504_));
  NA2        m0476(.A(mai_mai_n215_), .B(mai_mai_n101_), .Y(mai_mai_n505_));
  AOI210     m0477(.A0(mai_mai_n505_), .A1(mai_mai_n167_), .B0(mai_mai_n501_), .Y(mai_mai_n506_));
  AOI210     m0478(.A0(mai_mai_n346_), .A1(mai_mai_n35_), .B0(mai_mai_n470_), .Y(mai_mai_n507_));
  NOi31      m0479(.An(mai_mai_n504_), .B(mai_mai_n507_), .C(mai_mai_n506_), .Y(mai_mai_n508_));
  AN2        m0480(.A(mai_mai_n273_), .B(mai_mai_n249_), .Y(mai_mai_n509_));
  NA3        m0481(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n510_));
  NO2        m0482(.A(mai_mai_n510_), .B(mai_mai_n424_), .Y(mai_mai_n511_));
  NO2        m0483(.A(mai_mai_n511_), .B(mai_mai_n281_), .Y(mai_mai_n512_));
  NAi41      m0484(.An(mai_mai_n509_), .B(mai_mai_n512_), .C(mai_mai_n508_), .D(mai_mai_n503_), .Y(mai_mai_n513_));
  NO4        m0485(.A(mai_mai_n513_), .B(mai_mai_n500_), .C(mai_mai_n496_), .D(mai_mai_n493_), .Y(mai_mai_n514_));
  NA4        m0486(.A(mai_mai_n514_), .B(mai_mai_n485_), .C(mai_mai_n453_), .D(mai_mai_n419_), .Y(mai11));
  NO2        m0487(.A(mai_mai_n72_), .B(f), .Y(mai_mai_n516_));
  NA2        m0488(.A(j), .B(g), .Y(mai_mai_n517_));
  NAi31      m0489(.An(i), .B(m), .C(l), .Y(mai_mai_n518_));
  NA3        m0490(.A(m), .B(k), .C(j), .Y(mai_mai_n519_));
  OAI220     m0491(.A0(mai_mai_n519_), .A1(mai_mai_n122_), .B0(mai_mai_n518_), .B1(mai_mai_n517_), .Y(mai_mai_n520_));
  NA2        m0492(.A(mai_mai_n520_), .B(mai_mai_n516_), .Y(mai_mai_n521_));
  NOi32      m0493(.An(e), .Bn(b), .C(f), .Y(mai_mai_n522_));
  NA2        m0494(.A(mai_mai_n246_), .B(mai_mai_n106_), .Y(mai_mai_n523_));
  NA2        m0495(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n524_));
  NAi31      m0496(.An(d), .B(e), .C(a), .Y(mai_mai_n525_));
  NO2        m0497(.A(mai_mai_n525_), .B(n), .Y(mai_mai_n526_));
  NAi41      m0498(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n527_));
  AN2        m0499(.A(mai_mai_n527_), .B(mai_mai_n357_), .Y(mai_mai_n528_));
  AOI210     m0500(.A0(mai_mai_n528_), .A1(mai_mai_n382_), .B0(mai_mai_n257_), .Y(mai_mai_n529_));
  NA2        m0501(.A(j), .B(i), .Y(mai_mai_n530_));
  NAi31      m0502(.An(n), .B(m), .C(k), .Y(mai_mai_n531_));
  NO3        m0503(.A(mai_mai_n531_), .B(mai_mai_n530_), .C(mai_mai_n105_), .Y(mai_mai_n532_));
  NO4        m0504(.A(n), .B(d), .C(mai_mai_n109_), .D(a), .Y(mai_mai_n533_));
  OR2        m0505(.A(n), .B(c), .Y(mai_mai_n534_));
  NO2        m0506(.A(mai_mai_n534_), .B(mai_mai_n136_), .Y(mai_mai_n535_));
  NO2        m0507(.A(mai_mai_n535_), .B(mai_mai_n533_), .Y(mai_mai_n536_));
  NOi32      m0508(.An(g), .Bn(f), .C(i), .Y(mai_mai_n537_));
  AOI220     m0509(.A0(mai_mai_n537_), .A1(mai_mai_n94_), .B0(mai_mai_n520_), .B1(f), .Y(mai_mai_n538_));
  NO2        m0510(.A(mai_mai_n259_), .B(mai_mai_n49_), .Y(mai_mai_n539_));
  NO2        m0511(.A(mai_mai_n538_), .B(mai_mai_n536_), .Y(mai_mai_n540_));
  AOI210     m0512(.A0(mai_mai_n532_), .A1(mai_mai_n529_), .B0(mai_mai_n540_), .Y(mai_mai_n541_));
  NA2        m0513(.A(mai_mai_n129_), .B(mai_mai_n34_), .Y(mai_mai_n542_));
  OAI220     m0514(.A0(mai_mai_n542_), .A1(m), .B0(mai_mai_n524_), .B1(mai_mai_n221_), .Y(mai_mai_n543_));
  NOi41      m0515(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n544_));
  NAi32      m0516(.An(e), .Bn(b), .C(c), .Y(mai_mai_n545_));
  OR2        m0517(.A(mai_mai_n545_), .B(mai_mai_n81_), .Y(mai_mai_n546_));
  AN2        m0518(.A(mai_mai_n325_), .B(mai_mai_n305_), .Y(mai_mai_n547_));
  NA2        m0519(.A(mai_mai_n547_), .B(mai_mai_n546_), .Y(mai_mai_n548_));
  OA210      m0520(.A0(mai_mai_n548_), .A1(mai_mai_n544_), .B0(mai_mai_n543_), .Y(mai_mai_n549_));
  OAI220     m0521(.A0(mai_mai_n384_), .A1(mai_mai_n383_), .B0(mai_mai_n518_), .B1(mai_mai_n517_), .Y(mai_mai_n550_));
  NAi31      m0522(.An(d), .B(c), .C(a), .Y(mai_mai_n551_));
  NO2        m0523(.A(mai_mai_n551_), .B(n), .Y(mai_mai_n552_));
  NA3        m0524(.A(mai_mai_n552_), .B(mai_mai_n550_), .C(e), .Y(mai_mai_n553_));
  NO3        m0525(.A(mai_mai_n62_), .B(mai_mai_n49_), .C(mai_mai_n203_), .Y(mai_mai_n554_));
  NO2        m0526(.A(mai_mai_n218_), .B(mai_mai_n103_), .Y(mai_mai_n555_));
  OAI210     m0527(.A0(mai_mai_n554_), .A1(mai_mai_n385_), .B0(mai_mai_n555_), .Y(mai_mai_n556_));
  NA2        m0528(.A(mai_mai_n556_), .B(mai_mai_n553_), .Y(mai_mai_n557_));
  INV        m0529(.A(mai_mai_n414_), .Y(mai_mai_n558_));
  NA2        m0530(.A(mai_mai_n550_), .B(f), .Y(mai_mai_n559_));
  NAi32      m0531(.An(d), .Bn(a), .C(b), .Y(mai_mai_n560_));
  NO2        m0532(.A(mai_mai_n559_), .B(mai_mai_n558_), .Y(mai_mai_n561_));
  AN3        m0533(.A(j), .B(h), .C(g), .Y(mai_mai_n562_));
  NO2        m0534(.A(mai_mai_n133_), .B(c), .Y(mai_mai_n563_));
  NA3        m0535(.A(mai_mai_n563_), .B(mai_mai_n562_), .C(mai_mai_n448_), .Y(mai_mai_n564_));
  NA3        m0536(.A(f), .B(d), .C(b), .Y(mai_mai_n565_));
  NO4        m0537(.A(mai_mai_n565_), .B(mai_mai_n163_), .C(mai_mai_n160_), .D(g), .Y(mai_mai_n566_));
  INV        m0538(.A(mai_mai_n564_), .Y(mai_mai_n567_));
  NO4        m0539(.A(mai_mai_n567_), .B(mai_mai_n561_), .C(mai_mai_n557_), .D(mai_mai_n549_), .Y(mai_mai_n568_));
  AN3        m0540(.A(mai_mai_n568_), .B(mai_mai_n541_), .C(mai_mai_n521_), .Y(mai_mai_n569_));
  INV        m0541(.A(k), .Y(mai_mai_n570_));
  NA3        m0542(.A(l), .B(mai_mai_n570_), .C(i), .Y(mai_mai_n571_));
  INV        m0543(.A(mai_mai_n571_), .Y(mai_mai_n572_));
  NA4        m0544(.A(mai_mai_n381_), .B(mai_mai_n403_), .C(mai_mai_n168_), .D(mai_mai_n106_), .Y(mai_mai_n573_));
  NAi32      m0545(.An(h), .Bn(f), .C(g), .Y(mai_mai_n574_));
  NAi41      m0546(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n575_));
  OAI210     m0547(.A0(mai_mai_n525_), .A1(n), .B0(mai_mai_n575_), .Y(mai_mai_n576_));
  NA2        m0548(.A(mai_mai_n576_), .B(m), .Y(mai_mai_n577_));
  NAi31      m0549(.An(h), .B(g), .C(f), .Y(mai_mai_n578_));
  OR3        m0550(.A(mai_mai_n578_), .B(mai_mai_n261_), .C(mai_mai_n49_), .Y(mai_mai_n579_));
  NA4        m0551(.A(mai_mai_n403_), .B(mai_mai_n114_), .C(mai_mai_n106_), .D(e), .Y(mai_mai_n580_));
  AN2        m0552(.A(mai_mai_n580_), .B(mai_mai_n579_), .Y(mai_mai_n581_));
  OA210      m0553(.A0(mai_mai_n577_), .A1(mai_mai_n574_), .B0(mai_mai_n581_), .Y(mai_mai_n582_));
  NO3        m0554(.A(mai_mai_n574_), .B(mai_mai_n72_), .C(mai_mai_n74_), .Y(mai_mai_n583_));
  NO4        m0555(.A(mai_mai_n578_), .B(mai_mai_n534_), .C(mai_mai_n136_), .D(mai_mai_n74_), .Y(mai_mai_n584_));
  OR2        m0556(.A(mai_mai_n584_), .B(mai_mai_n583_), .Y(mai_mai_n585_));
  NAi31      m0557(.An(mai_mai_n585_), .B(mai_mai_n582_), .C(mai_mai_n573_), .Y(mai_mai_n586_));
  NAi31      m0558(.An(f), .B(h), .C(g), .Y(mai_mai_n587_));
  NO4        m0559(.A(mai_mai_n296_), .B(mai_mai_n587_), .C(mai_mai_n72_), .D(mai_mai_n74_), .Y(mai_mai_n588_));
  NOi32      m0560(.An(b), .Bn(a), .C(c), .Y(mai_mai_n589_));
  NOi41      m0561(.An(mai_mai_n589_), .B(mai_mai_n339_), .C(mai_mai_n69_), .D(mai_mai_n110_), .Y(mai_mai_n590_));
  OR2        m0562(.A(mai_mai_n590_), .B(mai_mai_n588_), .Y(mai_mai_n591_));
  NOi32      m0563(.An(d), .Bn(a), .C(e), .Y(mai_mai_n592_));
  NO2        m0564(.A(n), .B(c), .Y(mai_mai_n593_));
  NA3        m0565(.A(mai_mai_n593_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n594_));
  NAi32      m0566(.An(n), .Bn(f), .C(m), .Y(mai_mai_n595_));
  NA2        m0567(.A(mai_mai_n595_), .B(mai_mai_n594_), .Y(mai_mai_n596_));
  NOi32      m0568(.An(e), .Bn(a), .C(d), .Y(mai_mai_n597_));
  AOI210     m0569(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n597_), .Y(mai_mai_n598_));
  AOI210     m0570(.A0(mai_mai_n598_), .A1(mai_mai_n202_), .B0(mai_mai_n542_), .Y(mai_mai_n599_));
  AOI210     m0571(.A0(mai_mai_n599_), .A1(mai_mai_n596_), .B0(mai_mai_n591_), .Y(mai_mai_n600_));
  INV        m0572(.A(mai_mai_n600_), .Y(mai_mai_n601_));
  AOI210     m0573(.A0(mai_mai_n586_), .A1(mai_mai_n572_), .B0(mai_mai_n601_), .Y(mai_mai_n602_));
  NO3        m0574(.A(mai_mai_n303_), .B(mai_mai_n61_), .C(n), .Y(mai_mai_n603_));
  NA3        m0575(.A(mai_mai_n501_), .B(mai_mai_n158_), .C(mai_mai_n157_), .Y(mai_mai_n604_));
  NA2        m0576(.A(mai_mai_n450_), .B(mai_mai_n218_), .Y(mai_mai_n605_));
  OR2        m0577(.A(mai_mai_n605_), .B(mai_mai_n604_), .Y(mai_mai_n606_));
  NA2        m0578(.A(mai_mai_n75_), .B(mai_mai_n106_), .Y(mai_mai_n607_));
  NO2        m0579(.A(mai_mai_n607_), .B(mai_mai_n45_), .Y(mai_mai_n608_));
  AOI220     m0580(.A0(mai_mai_n608_), .A1(mai_mai_n529_), .B0(mai_mai_n606_), .B1(mai_mai_n603_), .Y(mai_mai_n609_));
  NO2        m0581(.A(mai_mai_n609_), .B(mai_mai_n84_), .Y(mai_mai_n610_));
  NOi32      m0582(.An(e), .Bn(c), .C(f), .Y(mai_mai_n611_));
  NOi21      m0583(.An(f), .B(g), .Y(mai_mai_n612_));
  NO2        m0584(.A(mai_mai_n612_), .B(mai_mai_n200_), .Y(mai_mai_n613_));
  AOI220     m0585(.A0(mai_mai_n613_), .A1(mai_mai_n378_), .B0(mai_mai_n611_), .B1(mai_mai_n162_), .Y(mai_mai_n614_));
  NA2        m0586(.A(mai_mai_n614_), .B(mai_mai_n165_), .Y(mai_mai_n615_));
  AOI210     m0587(.A0(mai_mai_n528_), .A1(mai_mai_n382_), .B0(mai_mai_n286_), .Y(mai_mai_n616_));
  NAi21      m0588(.An(k), .B(h), .Y(mai_mai_n617_));
  NO2        m0589(.A(mai_mai_n617_), .B(mai_mai_n248_), .Y(mai_mai_n618_));
  NOi31      m0590(.An(m), .B(n), .C(k), .Y(mai_mai_n619_));
  NA2        m0591(.A(j), .B(mai_mai_n619_), .Y(mai_mai_n620_));
  AOI210     m0592(.A0(mai_mai_n382_), .A1(mai_mai_n357_), .B0(mai_mai_n286_), .Y(mai_mai_n621_));
  NAi21      m0593(.An(mai_mai_n620_), .B(mai_mai_n621_), .Y(mai_mai_n622_));
  NO2        m0594(.A(mai_mai_n525_), .B(mai_mai_n49_), .Y(mai_mai_n623_));
  INV        m0595(.A(mai_mai_n622_), .Y(mai_mai_n624_));
  NA2        m0596(.A(mai_mai_n101_), .B(mai_mai_n36_), .Y(mai_mai_n625_));
  INV        m0597(.A(mai_mai_n348_), .Y(mai_mai_n626_));
  NO2        m0598(.A(mai_mai_n626_), .B(n), .Y(mai_mai_n627_));
  NO2        m0599(.A(mai_mai_n524_), .B(mai_mai_n163_), .Y(mai_mai_n628_));
  NA3        m0600(.A(mai_mai_n545_), .B(mai_mai_n256_), .C(mai_mai_n132_), .Y(mai_mai_n629_));
  NA2        m0601(.A(mai_mai_n497_), .B(mai_mai_n146_), .Y(mai_mai_n630_));
  NO3        m0602(.A(mai_mai_n379_), .B(mai_mai_n630_), .C(mai_mai_n84_), .Y(mai_mai_n631_));
  AOI210     m0603(.A0(mai_mai_n629_), .A1(mai_mai_n628_), .B0(mai_mai_n631_), .Y(mai_mai_n632_));
  AN3        m0604(.A(f), .B(d), .C(b), .Y(mai_mai_n633_));
  OAI210     m0605(.A0(mai_mai_n633_), .A1(mai_mai_n121_), .B0(n), .Y(mai_mai_n634_));
  NA3        m0606(.A(mai_mai_n497_), .B(mai_mai_n146_), .C(mai_mai_n203_), .Y(mai_mai_n635_));
  AOI210     m0607(.A0(mai_mai_n634_), .A1(mai_mai_n220_), .B0(mai_mai_n635_), .Y(mai_mai_n636_));
  NAi31      m0608(.An(m), .B(n), .C(k), .Y(mai_mai_n637_));
  INV        m0609(.A(mai_mai_n237_), .Y(mai_mai_n638_));
  OAI210     m0610(.A0(mai_mai_n638_), .A1(mai_mai_n636_), .B0(j), .Y(mai_mai_n639_));
  NA2        m0611(.A(mai_mai_n639_), .B(mai_mai_n632_), .Y(mai_mai_n640_));
  NO4        m0612(.A(mai_mai_n640_), .B(mai_mai_n624_), .C(mai_mai_n615_), .D(mai_mai_n610_), .Y(mai_mai_n641_));
  NA2        m0613(.A(mai_mai_n366_), .B(mai_mai_n149_), .Y(mai_mai_n642_));
  NAi31      m0614(.An(g), .B(h), .C(f), .Y(mai_mai_n643_));
  OR3        m0615(.A(mai_mai_n643_), .B(mai_mai_n261_), .C(n), .Y(mai_mai_n644_));
  OA210      m0616(.A0(mai_mai_n525_), .A1(n), .B0(mai_mai_n575_), .Y(mai_mai_n645_));
  NA3        m0617(.A(mai_mai_n401_), .B(mai_mai_n114_), .C(mai_mai_n81_), .Y(mai_mai_n646_));
  OAI210     m0618(.A0(mai_mai_n645_), .A1(mai_mai_n87_), .B0(mai_mai_n646_), .Y(mai_mai_n647_));
  NOi21      m0619(.An(mai_mai_n644_), .B(mai_mai_n647_), .Y(mai_mai_n648_));
  AOI210     m0620(.A0(mai_mai_n648_), .A1(mai_mai_n642_), .B0(mai_mai_n519_), .Y(mai_mai_n649_));
  NO3        m0621(.A(g), .B(mai_mai_n202_), .C(mai_mai_n56_), .Y(mai_mai_n650_));
  NAi21      m0622(.An(h), .B(j), .Y(mai_mai_n651_));
  NO2        m0623(.A(mai_mai_n505_), .B(mai_mai_n84_), .Y(mai_mai_n652_));
  OAI210     m0624(.A0(mai_mai_n652_), .A1(mai_mai_n378_), .B0(mai_mai_n650_), .Y(mai_mai_n653_));
  AN2        m0625(.A(h), .B(f), .Y(mai_mai_n654_));
  NA2        m0626(.A(mai_mai_n654_), .B(mai_mai_n37_), .Y(mai_mai_n655_));
  NA2        m0627(.A(mai_mai_n94_), .B(mai_mai_n46_), .Y(mai_mai_n656_));
  NO2        m0628(.A(mai_mai_n656_), .B(mai_mai_n318_), .Y(mai_mai_n657_));
  AOI210     m0629(.A0(mai_mai_n560_), .A1(mai_mai_n413_), .B0(mai_mai_n49_), .Y(mai_mai_n658_));
  OAI220     m0630(.A0(mai_mai_n578_), .A1(mai_mai_n571_), .B0(mai_mai_n312_), .B1(mai_mai_n517_), .Y(mai_mai_n659_));
  AOI210     m0631(.A0(mai_mai_n659_), .A1(mai_mai_n658_), .B0(mai_mai_n657_), .Y(mai_mai_n660_));
  NA2        m0632(.A(mai_mai_n660_), .B(mai_mai_n653_), .Y(mai_mai_n661_));
  NO2        m0633(.A(mai_mai_n238_), .B(f), .Y(mai_mai_n662_));
  NO2        m0634(.A(mai_mai_n612_), .B(mai_mai_n61_), .Y(mai_mai_n663_));
  NO3        m0635(.A(mai_mai_n663_), .B(mai_mai_n662_), .C(mai_mai_n34_), .Y(mai_mai_n664_));
  NA2        m0636(.A(mai_mai_n315_), .B(mai_mai_n129_), .Y(mai_mai_n665_));
  NA2        m0637(.A(mai_mai_n123_), .B(mai_mai_n49_), .Y(mai_mai_n666_));
  NA2        m0638(.A(mai_mai_n666_), .B(mai_mai_n522_), .Y(mai_mai_n667_));
  OA220      m0639(.A0(mai_mai_n667_), .A1(mai_mai_n542_), .B0(mai_mai_n346_), .B1(mai_mai_n104_), .Y(mai_mai_n668_));
  OAI210     m0640(.A0(mai_mai_n665_), .A1(mai_mai_n664_), .B0(mai_mai_n668_), .Y(mai_mai_n669_));
  NO3        m0641(.A(mai_mai_n389_), .B(mai_mai_n180_), .C(mai_mai_n179_), .Y(mai_mai_n670_));
  NA2        m0642(.A(mai_mai_n670_), .B(mai_mai_n218_), .Y(mai_mai_n671_));
  NA3        m0643(.A(mai_mai_n671_), .B(mai_mai_n240_), .C(j), .Y(mai_mai_n672_));
  NA2        m0644(.A(mai_mai_n454_), .B(mai_mai_n81_), .Y(mai_mai_n673_));
  NO4        m0645(.A(mai_mai_n519_), .B(mai_mai_n673_), .C(mai_mai_n122_), .D(mai_mai_n202_), .Y(mai_mai_n674_));
  INV        m0646(.A(mai_mai_n674_), .Y(mai_mai_n675_));
  NA4        m0647(.A(mai_mai_n675_), .B(mai_mai_n672_), .C(mai_mai_n504_), .D(mai_mai_n387_), .Y(mai_mai_n676_));
  NO4        m0648(.A(mai_mai_n676_), .B(mai_mai_n669_), .C(mai_mai_n661_), .D(mai_mai_n649_), .Y(mai_mai_n677_));
  NA4        m0649(.A(mai_mai_n677_), .B(mai_mai_n641_), .C(mai_mai_n602_), .D(mai_mai_n569_), .Y(mai08));
  NO2        m0650(.A(k), .B(h), .Y(mai_mai_n679_));
  AO210      m0651(.A0(mai_mai_n238_), .A1(mai_mai_n438_), .B0(mai_mai_n679_), .Y(mai_mai_n680_));
  NO2        m0652(.A(mai_mai_n680_), .B(mai_mai_n284_), .Y(mai_mai_n681_));
  NA2        m0653(.A(mai_mai_n611_), .B(mai_mai_n81_), .Y(mai_mai_n682_));
  NA2        m0654(.A(mai_mai_n682_), .B(mai_mai_n450_), .Y(mai_mai_n683_));
  AOI210     m0655(.A0(mai_mai_n683_), .A1(mai_mai_n681_), .B0(mai_mai_n482_), .Y(mai_mai_n684_));
  NA2        m0656(.A(mai_mai_n81_), .B(mai_mai_n103_), .Y(mai_mai_n685_));
  NO2        m0657(.A(mai_mai_n685_), .B(mai_mai_n57_), .Y(mai_mai_n686_));
  NO3        m0658(.A(mai_mai_n363_), .B(mai_mai_n105_), .C(mai_mai_n203_), .Y(mai_mai_n687_));
  NA2        m0659(.A(mai_mai_n565_), .B(mai_mai_n220_), .Y(mai_mai_n688_));
  AOI220     m0660(.A0(mai_mai_n688_), .A1(mai_mai_n334_), .B0(mai_mai_n687_), .B1(mai_mai_n686_), .Y(mai_mai_n689_));
  AOI210     m0661(.A0(mai_mai_n565_), .A1(mai_mai_n142_), .B0(mai_mai_n81_), .Y(mai_mai_n690_));
  NA4        m0662(.A(mai_mai_n205_), .B(mai_mai_n129_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n691_));
  AN2        m0663(.A(l), .B(k), .Y(mai_mai_n692_));
  NA4        m0664(.A(mai_mai_n692_), .B(mai_mai_n101_), .C(mai_mai_n74_), .D(mai_mai_n203_), .Y(mai_mai_n693_));
  OAI210     m0665(.A0(mai_mai_n691_), .A1(g), .B0(mai_mai_n693_), .Y(mai_mai_n694_));
  NA2        m0666(.A(mai_mai_n694_), .B(mai_mai_n690_), .Y(mai_mai_n695_));
  NA3        m0667(.A(mai_mai_n695_), .B(mai_mai_n689_), .C(mai_mai_n684_), .Y(mai_mai_n696_));
  NO4        m0668(.A(mai_mai_n160_), .B(mai_mai_n377_), .C(mai_mai_n105_), .D(g), .Y(mai_mai_n697_));
  NO2        m0669(.A(mai_mai_n528_), .B(mai_mai_n35_), .Y(mai_mai_n698_));
  INV        m0670(.A(mai_mai_n698_), .Y(mai_mai_n699_));
  NO3        m0671(.A(mai_mai_n303_), .B(mai_mai_n122_), .C(mai_mai_n41_), .Y(mai_mai_n700_));
  INV        m0672(.A(mai_mai_n693_), .Y(mai_mai_n701_));
  NA2        m0673(.A(mai_mai_n680_), .B(mai_mai_n126_), .Y(mai_mai_n702_));
  AOI220     m0674(.A0(mai_mai_n702_), .A1(mai_mai_n388_), .B0(mai_mai_n701_), .B1(mai_mai_n77_), .Y(mai_mai_n703_));
  OAI210     m0675(.A0(mai_mai_n699_), .A1(mai_mai_n84_), .B0(mai_mai_n703_), .Y(mai_mai_n704_));
  NA2        m0676(.A(mai_mai_n348_), .B(mai_mai_n43_), .Y(mai_mai_n705_));
  NA3        m0677(.A(mai_mai_n671_), .B(mai_mai_n320_), .C(mai_mai_n369_), .Y(mai_mai_n706_));
  NA2        m0678(.A(mai_mai_n692_), .B(mai_mai_n208_), .Y(mai_mai_n707_));
  NO2        m0679(.A(mai_mai_n707_), .B(mai_mai_n314_), .Y(mai_mai_n708_));
  AOI210     m0680(.A0(mai_mai_n708_), .A1(mai_mai_n662_), .B0(mai_mai_n481_), .Y(mai_mai_n709_));
  NA3        m0681(.A(m), .B(l), .C(k), .Y(mai_mai_n710_));
  AOI210     m0682(.A0(mai_mai_n646_), .A1(mai_mai_n644_), .B0(mai_mai_n710_), .Y(mai_mai_n711_));
  NO2        m0683(.A(mai_mai_n527_), .B(mai_mai_n257_), .Y(mai_mai_n712_));
  NOi21      m0684(.An(mai_mai_n712_), .B(mai_mai_n523_), .Y(mai_mai_n713_));
  NA4        m0685(.A(mai_mai_n106_), .B(l), .C(k), .D(mai_mai_n84_), .Y(mai_mai_n714_));
  NA3        m0686(.A(mai_mai_n114_), .B(mai_mai_n397_), .C(i), .Y(mai_mai_n715_));
  NO2        m0687(.A(mai_mai_n715_), .B(mai_mai_n714_), .Y(mai_mai_n716_));
  NO3        m0688(.A(mai_mai_n716_), .B(mai_mai_n713_), .C(mai_mai_n711_), .Y(mai_mai_n717_));
  NA4        m0689(.A(mai_mai_n717_), .B(mai_mai_n709_), .C(mai_mai_n706_), .D(mai_mai_n705_), .Y(mai_mai_n718_));
  NO4        m0690(.A(mai_mai_n718_), .B(mai_mai_n704_), .C(mai_mai_n511_), .D(mai_mai_n696_), .Y(mai_mai_n719_));
  NA2        m0691(.A(mai_mai_n613_), .B(mai_mai_n378_), .Y(mai_mai_n720_));
  NOi31      m0692(.An(g), .B(h), .C(f), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n623_), .B(mai_mai_n721_), .Y(mai_mai_n722_));
  AO210      m0694(.A0(mai_mai_n722_), .A1(mai_mai_n579_), .B0(mai_mai_n530_), .Y(mai_mai_n723_));
  NO3        m0695(.A(mai_mai_n382_), .B(mai_mai_n517_), .C(h), .Y(mai_mai_n724_));
  AOI210     m0696(.A0(mai_mai_n724_), .A1(mai_mai_n106_), .B0(mai_mai_n491_), .Y(mai_mai_n725_));
  NA4        m0697(.A(mai_mai_n725_), .B(mai_mai_n723_), .C(mai_mai_n720_), .D(mai_mai_n237_), .Y(mai_mai_n726_));
  NA2        m0698(.A(mai_mai_n692_), .B(mai_mai_n74_), .Y(mai_mai_n727_));
  NO4        m0699(.A(mai_mai_n670_), .B(mai_mai_n160_), .C(n), .D(i), .Y(mai_mai_n728_));
  NOi21      m0700(.An(h), .B(j), .Y(mai_mai_n729_));
  NA2        m0701(.A(mai_mai_n729_), .B(f), .Y(mai_mai_n730_));
  INV        m0702(.A(mai_mai_n728_), .Y(mai_mai_n731_));
  OAI220     m0703(.A0(mai_mai_n731_), .A1(mai_mai_n727_), .B0(mai_mai_n581_), .B1(mai_mai_n62_), .Y(mai_mai_n732_));
  AOI210     m0704(.A0(mai_mai_n726_), .A1(l), .B0(mai_mai_n732_), .Y(mai_mai_n733_));
  NO2        m0705(.A(j), .B(i), .Y(mai_mai_n734_));
  NA2        m0706(.A(mai_mai_n734_), .B(mai_mai_n33_), .Y(mai_mai_n735_));
  NA2        m0707(.A(mai_mai_n406_), .B(mai_mai_n114_), .Y(mai_mai_n736_));
  OR2        m0708(.A(mai_mai_n736_), .B(mai_mai_n735_), .Y(mai_mai_n737_));
  NO3        m0709(.A(mai_mai_n138_), .B(mai_mai_n49_), .C(mai_mai_n103_), .Y(mai_mai_n738_));
  NO3        m0710(.A(mai_mai_n534_), .B(mai_mai_n136_), .C(mai_mai_n74_), .Y(mai_mai_n739_));
  NO3        m0711(.A(mai_mai_n477_), .B(mai_mai_n425_), .C(j), .Y(mai_mai_n740_));
  OAI210     m0712(.A0(mai_mai_n739_), .A1(mai_mai_n738_), .B0(mai_mai_n740_), .Y(mai_mai_n741_));
  OAI210     m0713(.A0(mai_mai_n722_), .A1(mai_mai_n62_), .B0(mai_mai_n741_), .Y(mai_mai_n742_));
  NA2        m0714(.A(k), .B(j), .Y(mai_mai_n743_));
  NO3        m0715(.A(mai_mai_n284_), .B(mai_mai_n743_), .C(mai_mai_n40_), .Y(mai_mai_n744_));
  AOI210     m0716(.A0(mai_mai_n522_), .A1(n), .B0(mai_mai_n544_), .Y(mai_mai_n745_));
  NA2        m0717(.A(mai_mai_n745_), .B(mai_mai_n547_), .Y(mai_mai_n746_));
  AN3        m0718(.A(mai_mai_n746_), .B(mai_mai_n744_), .C(mai_mai_n93_), .Y(mai_mai_n747_));
  NA2        m0719(.A(mai_mai_n605_), .B(mai_mai_n293_), .Y(mai_mai_n748_));
  INV        m0720(.A(mai_mai_n748_), .Y(mai_mai_n749_));
  NO2        m0721(.A(mai_mai_n284_), .B(mai_mai_n126_), .Y(mai_mai_n750_));
  AOI220     m0722(.A0(mai_mai_n750_), .A1(mai_mai_n613_), .B0(mai_mai_n700_), .B1(mai_mai_n690_), .Y(mai_mai_n751_));
  NO2        m0723(.A(mai_mai_n710_), .B(mai_mai_n87_), .Y(mai_mai_n752_));
  NA2        m0724(.A(mai_mai_n752_), .B(mai_mai_n576_), .Y(mai_mai_n753_));
  NO2        m0725(.A(mai_mai_n578_), .B(mai_mai_n110_), .Y(mai_mai_n754_));
  OAI210     m0726(.A0(mai_mai_n754_), .A1(mai_mai_n740_), .B0(mai_mai_n658_), .Y(mai_mai_n755_));
  NA3        m0727(.A(mai_mai_n755_), .B(mai_mai_n753_), .C(mai_mai_n751_), .Y(mai_mai_n756_));
  OR4        m0728(.A(mai_mai_n756_), .B(mai_mai_n749_), .C(mai_mai_n747_), .D(mai_mai_n742_), .Y(mai_mai_n757_));
  NA3        m0729(.A(mai_mai_n745_), .B(mai_mai_n547_), .C(mai_mai_n546_), .Y(mai_mai_n758_));
  NA4        m0730(.A(mai_mai_n758_), .B(mai_mai_n205_), .C(mai_mai_n438_), .D(mai_mai_n34_), .Y(mai_mai_n759_));
  OAI220     m0731(.A0(mai_mai_n691_), .A1(mai_mai_n682_), .B0(mai_mai_n318_), .B1(mai_mai_n38_), .Y(mai_mai_n760_));
  INV        m0732(.A(mai_mai_n760_), .Y(mai_mai_n761_));
  NA3        m0733(.A(mai_mai_n537_), .B(mai_mai_n277_), .C(h), .Y(mai_mai_n762_));
  NOi21      m0734(.An(mai_mai_n658_), .B(mai_mai_n762_), .Y(mai_mai_n763_));
  NO2        m0735(.A(mai_mai_n88_), .B(mai_mai_n47_), .Y(mai_mai_n764_));
  NO2        m0736(.A(mai_mai_n762_), .B(mai_mai_n594_), .Y(mai_mai_n765_));
  AOI210     m0737(.A0(mai_mai_n764_), .A1(mai_mai_n627_), .B0(mai_mai_n765_), .Y(mai_mai_n766_));
  NAi41      m0738(.An(mai_mai_n763_), .B(mai_mai_n766_), .C(mai_mai_n761_), .D(mai_mai_n759_), .Y(mai_mai_n767_));
  NA2        m0739(.A(mai_mai_n752_), .B(mai_mai_n226_), .Y(mai_mai_n768_));
  INV        m0740(.A(mai_mai_n322_), .Y(mai_mai_n769_));
  OAI210     m0741(.A0(mai_mai_n710_), .A1(mai_mai_n643_), .B0(mai_mai_n510_), .Y(mai_mai_n770_));
  NA3        m0742(.A(mai_mai_n236_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n771_));
  AOI220     m0743(.A0(mai_mai_n593_), .A1(mai_mai_n29_), .B0(mai_mai_n454_), .B1(mai_mai_n81_), .Y(mai_mai_n772_));
  NA2        m0744(.A(mai_mai_n772_), .B(mai_mai_n771_), .Y(mai_mai_n773_));
  NO2        m0745(.A(mai_mai_n762_), .B(mai_mai_n480_), .Y(mai_mai_n774_));
  AOI210     m0746(.A0(mai_mai_n773_), .A1(mai_mai_n770_), .B0(mai_mai_n774_), .Y(mai_mai_n775_));
  NA3        m0747(.A(mai_mai_n775_), .B(mai_mai_n769_), .C(mai_mai_n768_), .Y(mai_mai_n776_));
  NOi41      m0748(.An(mai_mai_n737_), .B(mai_mai_n776_), .C(mai_mai_n767_), .D(mai_mai_n757_), .Y(mai_mai_n777_));
  OR3        m0749(.A(mai_mai_n691_), .B(mai_mai_n220_), .C(g), .Y(mai_mai_n778_));
  NO3        m0750(.A(mai_mai_n328_), .B(mai_mai_n286_), .C(mai_mai_n105_), .Y(mai_mai_n779_));
  NA2        m0751(.A(mai_mai_n779_), .B(mai_mai_n746_), .Y(mai_mai_n780_));
  NA2        m0752(.A(mai_mai_n46_), .B(mai_mai_n56_), .Y(mai_mai_n781_));
  NO3        m0753(.A(mai_mai_n781_), .B(mai_mai_n735_), .C(mai_mai_n261_), .Y(mai_mai_n782_));
  INV        m0754(.A(mai_mai_n782_), .Y(mai_mai_n783_));
  NA4        m0755(.A(mai_mai_n783_), .B(mai_mai_n780_), .C(mai_mai_n778_), .D(mai_mai_n390_), .Y(mai_mai_n784_));
  OR2        m0756(.A(mai_mai_n643_), .B(mai_mai_n88_), .Y(mai_mai_n785_));
  NOi31      m0757(.An(b), .B(d), .C(a), .Y(mai_mai_n786_));
  NO2        m0758(.A(mai_mai_n786_), .B(mai_mai_n592_), .Y(mai_mai_n787_));
  NO2        m0759(.A(mai_mai_n787_), .B(n), .Y(mai_mai_n788_));
  NO2        m0760(.A(mai_mai_n545_), .B(mai_mai_n81_), .Y(mai_mai_n789_));
  NA2        m0761(.A(mai_mai_n779_), .B(mai_mai_n789_), .Y(mai_mai_n790_));
  OAI210     m0762(.A0(mai_mai_n691_), .A1(mai_mai_n379_), .B0(mai_mai_n790_), .Y(mai_mai_n791_));
  NO2        m0763(.A(mai_mai_n670_), .B(n), .Y(mai_mai_n792_));
  AOI220     m0764(.A0(mai_mai_n750_), .A1(mai_mai_n650_), .B0(mai_mai_n792_), .B1(mai_mai_n681_), .Y(mai_mai_n793_));
  NA2        m0765(.A(mai_mai_n114_), .B(mai_mai_n81_), .Y(mai_mai_n794_));
  AOI210     m0766(.A0(mai_mai_n410_), .A1(mai_mai_n402_), .B0(mai_mai_n794_), .Y(mai_mai_n795_));
  NA2        m0767(.A(mai_mai_n708_), .B(mai_mai_n34_), .Y(mai_mai_n796_));
  NAi21      m0768(.An(mai_mai_n714_), .B(mai_mai_n421_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n257_), .B(i), .Y(mai_mai_n798_));
  NA2        m0770(.A(mai_mai_n697_), .B(mai_mai_n335_), .Y(mai_mai_n799_));
  OAI210     m0771(.A0(mai_mai_n584_), .A1(mai_mai_n583_), .B0(mai_mai_n349_), .Y(mai_mai_n800_));
  AN3        m0772(.A(mai_mai_n800_), .B(mai_mai_n799_), .C(mai_mai_n797_), .Y(mai_mai_n801_));
  NAi41      m0773(.An(mai_mai_n795_), .B(mai_mai_n801_), .C(mai_mai_n796_), .D(mai_mai_n793_), .Y(mai_mai_n802_));
  NO3        m0774(.A(mai_mai_n802_), .B(mai_mai_n791_), .C(mai_mai_n784_), .Y(mai_mai_n803_));
  NA4        m0775(.A(mai_mai_n803_), .B(mai_mai_n777_), .C(mai_mai_n733_), .D(mai_mai_n719_), .Y(mai09));
  INV        m0776(.A(mai_mai_n115_), .Y(mai_mai_n805_));
  NA2        m0777(.A(f), .B(e), .Y(mai_mai_n806_));
  NO2        m0778(.A(mai_mai_n213_), .B(mai_mai_n105_), .Y(mai_mai_n807_));
  NA2        m0779(.A(mai_mai_n807_), .B(g), .Y(mai_mai_n808_));
  NA4        m0780(.A(mai_mai_n296_), .B(mai_mai_n463_), .C(mai_mai_n247_), .D(mai_mai_n112_), .Y(mai_mai_n809_));
  AOI210     m0781(.A0(mai_mai_n809_), .A1(g), .B0(mai_mai_n460_), .Y(mai_mai_n810_));
  AOI210     m0782(.A0(mai_mai_n810_), .A1(mai_mai_n808_), .B0(mai_mai_n806_), .Y(mai_mai_n811_));
  NA2        m0783(.A(mai_mai_n811_), .B(mai_mai_n805_), .Y(mai_mai_n812_));
  NO2        m0784(.A(mai_mai_n192_), .B(mai_mai_n202_), .Y(mai_mai_n813_));
  NA3        m0785(.A(m), .B(l), .C(i), .Y(mai_mai_n814_));
  OAI220     m0786(.A0(mai_mai_n578_), .A1(mai_mai_n814_), .B0(mai_mai_n339_), .B1(mai_mai_n518_), .Y(mai_mai_n815_));
  NA4        m0787(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(g), .D(f), .Y(mai_mai_n816_));
  NAi31      m0788(.An(mai_mai_n815_), .B(mai_mai_n816_), .C(mai_mai_n426_), .Y(mai_mai_n817_));
  OR2        m0789(.A(mai_mai_n817_), .B(mai_mai_n813_), .Y(mai_mai_n818_));
  NA3        m0790(.A(mai_mai_n785_), .B(mai_mai_n559_), .C(mai_mai_n510_), .Y(mai_mai_n819_));
  OA210      m0791(.A0(mai_mai_n819_), .A1(mai_mai_n818_), .B0(mai_mai_n788_), .Y(mai_mai_n820_));
  INV        m0792(.A(mai_mai_n325_), .Y(mai_mai_n821_));
  NO2        m0793(.A(mai_mai_n120_), .B(mai_mai_n119_), .Y(mai_mai_n822_));
  NOi31      m0794(.An(k), .B(m), .C(l), .Y(mai_mai_n823_));
  NO2        m0795(.A(mai_mai_n327_), .B(mai_mai_n823_), .Y(mai_mai_n824_));
  AOI210     m0796(.A0(mai_mai_n824_), .A1(mai_mai_n822_), .B0(mai_mai_n587_), .Y(mai_mai_n825_));
  NA2        m0797(.A(mai_mai_n771_), .B(mai_mai_n318_), .Y(mai_mai_n826_));
  NA2        m0798(.A(mai_mai_n329_), .B(mai_mai_n331_), .Y(mai_mai_n827_));
  OAI210     m0799(.A0(mai_mai_n192_), .A1(mai_mai_n202_), .B0(mai_mai_n827_), .Y(mai_mai_n828_));
  AOI220     m0800(.A0(mai_mai_n828_), .A1(mai_mai_n826_), .B0(mai_mai_n825_), .B1(mai_mai_n821_), .Y(mai_mai_n829_));
  NA2        m0801(.A(mai_mai_n154_), .B(mai_mai_n107_), .Y(mai_mai_n830_));
  NA3        m0802(.A(mai_mai_n830_), .B(mai_mai_n680_), .C(mai_mai_n126_), .Y(mai_mai_n831_));
  NA3        m0803(.A(mai_mai_n831_), .B(mai_mai_n177_), .C(mai_mai_n31_), .Y(mai_mai_n832_));
  NA3        m0804(.A(mai_mai_n832_), .B(mai_mai_n829_), .C(mai_mai_n614_), .Y(mai_mai_n833_));
  NO2        m0805(.A(mai_mai_n574_), .B(mai_mai_n488_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n834_), .B(mai_mai_n177_), .Y(mai_mai_n835_));
  NOi21      m0807(.An(f), .B(d), .Y(mai_mai_n836_));
  NA2        m0808(.A(mai_mai_n836_), .B(m), .Y(mai_mai_n837_));
  NO2        m0809(.A(mai_mai_n837_), .B(mai_mai_n52_), .Y(mai_mai_n838_));
  NOi32      m0810(.An(g), .Bn(f), .C(d), .Y(mai_mai_n839_));
  NA4        m0811(.A(mai_mai_n839_), .B(mai_mai_n593_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n840_));
  NOi21      m0812(.An(mai_mai_n297_), .B(mai_mai_n840_), .Y(mai_mai_n841_));
  AOI210     m0813(.A0(mai_mai_n838_), .A1(mai_mai_n535_), .B0(mai_mai_n841_), .Y(mai_mai_n842_));
  NA2        m0814(.A(mai_mai_n247_), .B(mai_mai_n112_), .Y(mai_mai_n843_));
  AN2        m0815(.A(f), .B(d), .Y(mai_mai_n844_));
  NA3        m0816(.A(mai_mai_n468_), .B(mai_mai_n844_), .C(mai_mai_n81_), .Y(mai_mai_n845_));
  NO3        m0817(.A(mai_mai_n845_), .B(mai_mai_n74_), .C(mai_mai_n203_), .Y(mai_mai_n846_));
  NO2        m0818(.A(mai_mai_n270_), .B(mai_mai_n56_), .Y(mai_mai_n847_));
  NA2        m0819(.A(mai_mai_n843_), .B(mai_mai_n846_), .Y(mai_mai_n848_));
  NAi41      m0820(.An(mai_mai_n479_), .B(mai_mai_n848_), .C(mai_mai_n842_), .D(mai_mai_n835_), .Y(mai_mai_n849_));
  NO4        m0821(.A(mai_mai_n612_), .B(mai_mai_n123_), .C(mai_mai_n314_), .D(mai_mai_n139_), .Y(mai_mai_n850_));
  NO2        m0822(.A(mai_mai_n637_), .B(mai_mai_n314_), .Y(mai_mai_n851_));
  AN2        m0823(.A(mai_mai_n851_), .B(mai_mai_n662_), .Y(mai_mai_n852_));
  NO3        m0824(.A(mai_mai_n852_), .B(mai_mai_n850_), .C(mai_mai_n222_), .Y(mai_mai_n853_));
  NA2        m0825(.A(mai_mai_n592_), .B(mai_mai_n81_), .Y(mai_mai_n854_));
  NA3        m0826(.A(mai_mai_n146_), .B(mai_mai_n101_), .C(mai_mai_n100_), .Y(mai_mai_n855_));
  OAI220     m0827(.A0(mai_mai_n845_), .A1(mai_mai_n415_), .B0(mai_mai_n325_), .B1(mai_mai_n855_), .Y(mai_mai_n856_));
  NOi31      m0828(.An(mai_mai_n211_), .B(mai_mai_n856_), .C(mai_mai_n291_), .Y(mai_mai_n857_));
  NA2        m0829(.A(c), .B(mai_mai_n109_), .Y(mai_mai_n858_));
  NO2        m0830(.A(mai_mai_n858_), .B(mai_mai_n394_), .Y(mai_mai_n859_));
  NA3        m0831(.A(mai_mai_n859_), .B(mai_mai_n499_), .C(f), .Y(mai_mai_n860_));
  OR2        m0832(.A(mai_mai_n643_), .B(mai_mai_n531_), .Y(mai_mai_n861_));
  INV        m0833(.A(mai_mai_n861_), .Y(mai_mai_n862_));
  NA2        m0834(.A(mai_mai_n787_), .B(mai_mai_n104_), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n863_), .B(mai_mai_n862_), .Y(mai_mai_n864_));
  NA4        m0836(.A(mai_mai_n864_), .B(mai_mai_n860_), .C(mai_mai_n857_), .D(mai_mai_n853_), .Y(mai_mai_n865_));
  NO4        m0837(.A(mai_mai_n865_), .B(mai_mai_n849_), .C(mai_mai_n833_), .D(mai_mai_n820_), .Y(mai_mai_n866_));
  OR2        m0838(.A(mai_mai_n845_), .B(mai_mai_n74_), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n105_), .B(j), .Y(mai_mai_n868_));
  NA2        m0840(.A(mai_mai_n807_), .B(g), .Y(mai_mai_n869_));
  AOI210     m0841(.A0(mai_mai_n869_), .A1(mai_mai_n278_), .B0(mai_mai_n867_), .Y(mai_mai_n870_));
  NO2        m0842(.A(mai_mai_n318_), .B(mai_mai_n816_), .Y(mai_mai_n871_));
  NO2        m0843(.A(mai_mai_n218_), .B(mai_mai_n212_), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n872_), .B(mai_mai_n215_), .Y(mai_mai_n873_));
  NO2        m0845(.A(mai_mai_n415_), .B(mai_mai_n806_), .Y(mai_mai_n874_));
  NA2        m0846(.A(mai_mai_n874_), .B(mai_mai_n552_), .Y(mai_mai_n875_));
  NA2        m0847(.A(mai_mai_n875_), .B(mai_mai_n873_), .Y(mai_mai_n876_));
  NA2        m0848(.A(e), .B(d), .Y(mai_mai_n877_));
  OAI220     m0849(.A0(mai_mai_n877_), .A1(c), .B0(mai_mai_n309_), .B1(d), .Y(mai_mai_n878_));
  NA3        m0850(.A(mai_mai_n878_), .B(mai_mai_n443_), .C(mai_mai_n497_), .Y(mai_mai_n879_));
  AOI210     m0851(.A0(mai_mai_n505_), .A1(mai_mai_n167_), .B0(mai_mai_n218_), .Y(mai_mai_n880_));
  INV        m0852(.A(mai_mai_n880_), .Y(mai_mai_n881_));
  NA2        m0853(.A(mai_mai_n270_), .B(mai_mai_n152_), .Y(mai_mai_n882_));
  NA2        m0854(.A(mai_mai_n846_), .B(mai_mai_n882_), .Y(mai_mai_n883_));
  NA3        m0855(.A(mai_mai_n153_), .B(mai_mai_n82_), .C(mai_mai_n34_), .Y(mai_mai_n884_));
  NA4        m0856(.A(mai_mai_n884_), .B(mai_mai_n883_), .C(mai_mai_n881_), .D(mai_mai_n879_), .Y(mai_mai_n885_));
  NO4        m0857(.A(mai_mai_n885_), .B(mai_mai_n876_), .C(mai_mai_n871_), .D(mai_mai_n870_), .Y(mai_mai_n886_));
  NA2        m0858(.A(mai_mai_n821_), .B(mai_mai_n31_), .Y(mai_mai_n887_));
  AO210      m0859(.A0(mai_mai_n887_), .A1(mai_mai_n682_), .B0(mai_mai_n206_), .Y(mai_mai_n888_));
  OAI220     m0860(.A0(mai_mai_n612_), .A1(mai_mai_n61_), .B0(mai_mai_n286_), .B1(j), .Y(mai_mai_n889_));
  AOI220     m0861(.A0(mai_mai_n889_), .A1(mai_mai_n851_), .B0(mai_mai_n603_), .B1(mai_mai_n611_), .Y(mai_mai_n890_));
  INV        m0862(.A(mai_mai_n890_), .Y(mai_mai_n891_));
  OAI210     m0863(.A0(mai_mai_n807_), .A1(mai_mai_n882_), .B0(mai_mai_n839_), .Y(mai_mai_n892_));
  NO2        m0864(.A(mai_mai_n892_), .B(mai_mai_n594_), .Y(mai_mai_n893_));
  AOI210     m0865(.A0(mai_mai_n111_), .A1(mai_mai_n110_), .B0(mai_mai_n246_), .Y(mai_mai_n894_));
  NO2        m0866(.A(mai_mai_n894_), .B(mai_mai_n840_), .Y(mai_mai_n895_));
  BUFFER     m0867(.A(mai_mai_n895_), .Y(mai_mai_n896_));
  NOi31      m0868(.An(mai_mai_n535_), .B(mai_mai_n837_), .C(mai_mai_n278_), .Y(mai_mai_n897_));
  NO4        m0869(.A(mai_mai_n897_), .B(mai_mai_n896_), .C(mai_mai_n893_), .D(mai_mai_n891_), .Y(mai_mai_n898_));
  AO220      m0870(.A0(mai_mai_n443_), .A1(mai_mai_n729_), .B0(mai_mai_n162_), .B1(f), .Y(mai_mai_n899_));
  OAI210     m0871(.A0(mai_mai_n899_), .A1(mai_mai_n446_), .B0(mai_mai_n878_), .Y(mai_mai_n900_));
  NO2        m0872(.A(mai_mai_n425_), .B(mai_mai_n71_), .Y(mai_mai_n901_));
  OAI210     m0873(.A0(mai_mai_n819_), .A1(mai_mai_n901_), .B0(mai_mai_n686_), .Y(mai_mai_n902_));
  AN4        m0874(.A(mai_mai_n902_), .B(mai_mai_n900_), .C(mai_mai_n898_), .D(mai_mai_n888_), .Y(mai_mai_n903_));
  NA4        m0875(.A(mai_mai_n903_), .B(mai_mai_n886_), .C(mai_mai_n866_), .D(mai_mai_n812_), .Y(mai12));
  NO2        m0876(.A(mai_mai_n441_), .B(c), .Y(mai_mai_n905_));
  NO4        m0877(.A(mai_mai_n430_), .B(mai_mai_n238_), .C(mai_mai_n570_), .D(mai_mai_n203_), .Y(mai_mai_n906_));
  NA2        m0878(.A(mai_mai_n906_), .B(mai_mai_n905_), .Y(mai_mai_n907_));
  NA2        m0879(.A(mai_mai_n535_), .B(mai_mai_n901_), .Y(mai_mai_n908_));
  NO2        m0880(.A(mai_mai_n441_), .B(mai_mai_n109_), .Y(mai_mai_n909_));
  NO2        m0881(.A(mai_mai_n822_), .B(mai_mai_n339_), .Y(mai_mai_n910_));
  NO2        m0882(.A(mai_mai_n643_), .B(mai_mai_n363_), .Y(mai_mai_n911_));
  AOI220     m0883(.A0(mai_mai_n911_), .A1(mai_mai_n533_), .B0(mai_mai_n910_), .B1(mai_mai_n909_), .Y(mai_mai_n912_));
  NA4        m0884(.A(mai_mai_n912_), .B(mai_mai_n908_), .C(mai_mai_n907_), .D(mai_mai_n429_), .Y(mai_mai_n913_));
  AOI210     m0885(.A0(mai_mai_n221_), .A1(mai_mai_n324_), .B0(mai_mai_n189_), .Y(mai_mai_n914_));
  OR2        m0886(.A(mai_mai_n914_), .B(mai_mai_n906_), .Y(mai_mai_n915_));
  AOI210     m0887(.A0(mai_mai_n321_), .A1(mai_mai_n375_), .B0(mai_mai_n203_), .Y(mai_mai_n916_));
  OAI210     m0888(.A0(mai_mai_n916_), .A1(mai_mai_n915_), .B0(mai_mai_n389_), .Y(mai_mai_n917_));
  NO2        m0889(.A(mai_mai_n625_), .B(mai_mai_n248_), .Y(mai_mai_n918_));
  NO2        m0890(.A(mai_mai_n578_), .B(mai_mai_n814_), .Y(mai_mai_n919_));
  NO2        m0891(.A(mai_mai_n138_), .B(mai_mai_n225_), .Y(mai_mai_n920_));
  NA3        m0892(.A(mai_mai_n920_), .B(mai_mai_n228_), .C(i), .Y(mai_mai_n921_));
  NA2        m0893(.A(mai_mai_n921_), .B(mai_mai_n917_), .Y(mai_mai_n922_));
  NO3        m0894(.A(mai_mai_n123_), .B(mai_mai_n139_), .C(mai_mai_n203_), .Y(mai_mai_n923_));
  NA2        m0895(.A(mai_mai_n923_), .B(mai_mai_n522_), .Y(mai_mai_n924_));
  INV        m0896(.A(mai_mai_n924_), .Y(mai_mai_n925_));
  NO3        m0897(.A(mai_mai_n648_), .B(mai_mai_n88_), .C(mai_mai_n45_), .Y(mai_mai_n926_));
  NO4        m0898(.A(mai_mai_n926_), .B(mai_mai_n925_), .C(mai_mai_n922_), .D(mai_mai_n913_), .Y(mai_mai_n927_));
  NO2        m0899(.A(mai_mai_n354_), .B(mai_mai_n353_), .Y(mai_mai_n928_));
  NA2        m0900(.A(mai_mai_n575_), .B(mai_mai_n72_), .Y(mai_mai_n929_));
  NA2        m0901(.A(mai_mai_n545_), .B(mai_mai_n132_), .Y(mai_mai_n930_));
  NOi21      m0902(.An(mai_mai_n34_), .B(mai_mai_n637_), .Y(mai_mai_n931_));
  AOI220     m0903(.A0(mai_mai_n931_), .A1(mai_mai_n930_), .B0(mai_mai_n929_), .B1(mai_mai_n928_), .Y(mai_mai_n932_));
  OAI210     m0904(.A0(mai_mai_n237_), .A1(mai_mai_n45_), .B0(mai_mai_n932_), .Y(mai_mai_n933_));
  NA2        m0905(.A(mai_mai_n421_), .B(mai_mai_n250_), .Y(mai_mai_n934_));
  NO3        m0906(.A(mai_mai_n794_), .B(mai_mai_n86_), .C(mai_mai_n394_), .Y(mai_mai_n935_));
  NAi31      m0907(.An(mai_mai_n935_), .B(mai_mai_n934_), .C(mai_mai_n307_), .Y(mai_mai_n936_));
  NO2        m0908(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n937_));
  NO2        m0909(.A(mai_mai_n494_), .B(mai_mai_n286_), .Y(mai_mai_n938_));
  INV        m0910(.A(mai_mai_n938_), .Y(mai_mai_n939_));
  NO2        m0911(.A(mai_mai_n939_), .B(mai_mai_n132_), .Y(mai_mai_n940_));
  NA2        m0912(.A(mai_mai_n619_), .B(mai_mai_n349_), .Y(mai_mai_n941_));
  OAI210     m0913(.A0(mai_mai_n715_), .A1(mai_mai_n941_), .B0(mai_mai_n351_), .Y(mai_mai_n942_));
  NO4        m0914(.A(mai_mai_n942_), .B(mai_mai_n940_), .C(mai_mai_n936_), .D(mai_mai_n933_), .Y(mai_mai_n943_));
  NA2        m0915(.A(mai_mai_n333_), .B(g), .Y(mai_mai_n944_));
  NA2        m0916(.A(mai_mai_n149_), .B(i), .Y(mai_mai_n945_));
  NA2        m0917(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n946_));
  OAI220     m0918(.A0(mai_mai_n946_), .A1(mai_mai_n188_), .B0(mai_mai_n945_), .B1(mai_mai_n88_), .Y(mai_mai_n947_));
  AOI210     m0919(.A0(mai_mai_n404_), .A1(mai_mai_n37_), .B0(mai_mai_n947_), .Y(mai_mai_n948_));
  NO2        m0920(.A(mai_mai_n132_), .B(mai_mai_n81_), .Y(mai_mai_n949_));
  OR2        m0921(.A(mai_mai_n949_), .B(mai_mai_n544_), .Y(mai_mai_n950_));
  NA2        m0922(.A(mai_mai_n545_), .B(mai_mai_n367_), .Y(mai_mai_n951_));
  AOI210     m0923(.A0(mai_mai_n951_), .A1(n), .B0(mai_mai_n950_), .Y(mai_mai_n952_));
  OAI220     m0924(.A0(mai_mai_n952_), .A1(mai_mai_n944_), .B0(mai_mai_n948_), .B1(mai_mai_n318_), .Y(mai_mai_n953_));
  NA3        m0925(.A(mai_mai_n311_), .B(mai_mai_n111_), .C(g), .Y(mai_mai_n954_));
  AOI210     m0926(.A0(mai_mai_n655_), .A1(mai_mai_n954_), .B0(m), .Y(mai_mai_n955_));
  OAI210     m0927(.A0(mai_mai_n955_), .A1(mai_mai_n910_), .B0(mai_mai_n310_), .Y(mai_mai_n956_));
  NA2        m0928(.A(mai_mai_n673_), .B(mai_mai_n854_), .Y(mai_mai_n957_));
  NA2        m0929(.A(mai_mai_n816_), .B(mai_mai_n426_), .Y(mai_mai_n958_));
  NA2        m0930(.A(mai_mai_n958_), .B(mai_mai_n957_), .Y(mai_mai_n959_));
  NA2        m0931(.A(mai_mai_n959_), .B(mai_mai_n956_), .Y(mai_mai_n960_));
  NO2        m0932(.A(mai_mai_n363_), .B(mai_mai_n87_), .Y(mai_mai_n961_));
  OAI210     m0933(.A0(mai_mai_n961_), .A1(mai_mai_n918_), .B0(mai_mai_n226_), .Y(mai_mai_n962_));
  NA2        m0934(.A(mai_mai_n647_), .B(mai_mai_n85_), .Y(mai_mai_n963_));
  NO2        m0935(.A(mai_mai_n449_), .B(mai_mai_n203_), .Y(mai_mai_n964_));
  NA2        m0936(.A(mai_mai_n964_), .B(mai_mai_n368_), .Y(mai_mai_n965_));
  NA2        m0937(.A(mai_mai_n911_), .B(mai_mai_n920_), .Y(mai_mai_n966_));
  NA4        m0938(.A(mai_mai_n966_), .B(mai_mai_n965_), .C(mai_mai_n963_), .D(mai_mai_n962_), .Y(mai_mai_n967_));
  OAI210     m0939(.A0(mai_mai_n958_), .A1(mai_mai_n919_), .B0(mai_mai_n533_), .Y(mai_mai_n968_));
  AOI210     m0940(.A0(mai_mai_n405_), .A1(mai_mai_n398_), .B0(mai_mai_n794_), .Y(mai_mai_n969_));
  OAI210     m0941(.A0(mai_mai_n354_), .A1(mai_mai_n353_), .B0(mai_mai_n102_), .Y(mai_mai_n970_));
  AOI210     m0942(.A0(mai_mai_n970_), .A1(mai_mai_n526_), .B0(mai_mai_n969_), .Y(mai_mai_n971_));
  NA2        m0943(.A(mai_mai_n955_), .B(mai_mai_n909_), .Y(mai_mai_n972_));
  NO3        m0944(.A(mai_mai_n868_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n973_));
  NA2        m0945(.A(mai_mai_n973_), .B(mai_mai_n616_), .Y(mai_mai_n974_));
  NA4        m0946(.A(mai_mai_n974_), .B(mai_mai_n972_), .C(mai_mai_n971_), .D(mai_mai_n968_), .Y(mai_mai_n975_));
  NO4        m0947(.A(mai_mai_n975_), .B(mai_mai_n967_), .C(mai_mai_n960_), .D(mai_mai_n953_), .Y(mai_mai_n976_));
  NAi31      m0948(.An(mai_mai_n130_), .B(mai_mai_n406_), .C(n), .Y(mai_mai_n977_));
  NO3        m0949(.A(mai_mai_n119_), .B(mai_mai_n327_), .C(mai_mai_n823_), .Y(mai_mai_n978_));
  NO2        m0950(.A(mai_mai_n978_), .B(mai_mai_n977_), .Y(mai_mai_n979_));
  NO3        m0951(.A(mai_mai_n257_), .B(mai_mai_n130_), .C(mai_mai_n394_), .Y(mai_mai_n980_));
  AOI210     m0952(.A0(mai_mai_n980_), .A1(mai_mai_n489_), .B0(mai_mai_n979_), .Y(mai_mai_n981_));
  NA2        m0953(.A(mai_mai_n482_), .B(i), .Y(mai_mai_n982_));
  NA2        m0954(.A(mai_mai_n982_), .B(mai_mai_n981_), .Y(mai_mai_n983_));
  NA2        m0955(.A(mai_mai_n218_), .B(mai_mai_n158_), .Y(mai_mai_n984_));
  NO3        m0956(.A(mai_mai_n293_), .B(mai_mai_n431_), .C(mai_mai_n162_), .Y(mai_mai_n985_));
  NOi31      m0957(.An(mai_mai_n984_), .B(mai_mai_n985_), .C(mai_mai_n203_), .Y(mai_mai_n986_));
  NAi21      m0958(.An(mai_mai_n545_), .B(mai_mai_n964_), .Y(mai_mai_n987_));
  NA2        m0959(.A(mai_mai_n424_), .B(mai_mai_n854_), .Y(mai_mai_n988_));
  NO3        m0960(.A(mai_mai_n425_), .B(mai_mai_n296_), .C(mai_mai_n74_), .Y(mai_mai_n989_));
  AOI220     m0961(.A0(mai_mai_n989_), .A1(mai_mai_n988_), .B0(mai_mai_n474_), .B1(g), .Y(mai_mai_n990_));
  NA2        m0962(.A(mai_mai_n990_), .B(mai_mai_n987_), .Y(mai_mai_n991_));
  NO2        m0963(.A(mai_mai_n644_), .B(mai_mai_n363_), .Y(mai_mai_n992_));
  NA2        m0964(.A(mai_mai_n914_), .B(mai_mai_n905_), .Y(mai_mai_n993_));
  NO3        m0965(.A(mai_mai_n534_), .B(mai_mai_n136_), .C(mai_mai_n202_), .Y(mai_mai_n994_));
  OAI210     m0966(.A0(mai_mai_n994_), .A1(mai_mai_n516_), .B0(mai_mai_n364_), .Y(mai_mai_n995_));
  OAI220     m0967(.A0(mai_mai_n911_), .A1(mai_mai_n919_), .B0(mai_mai_n535_), .B1(mai_mai_n414_), .Y(mai_mai_n996_));
  NA3        m0968(.A(mai_mai_n996_), .B(mai_mai_n995_), .C(mai_mai_n993_), .Y(mai_mai_n997_));
  OAI210     m0969(.A0(mai_mai_n914_), .A1(mai_mai_n906_), .B0(mai_mai_n984_), .Y(mai_mai_n998_));
  NA3        m0970(.A(mai_mai_n951_), .B(mai_mai_n478_), .C(mai_mai_n46_), .Y(mai_mai_n999_));
  NA2        m0971(.A(mai_mai_n366_), .B(mai_mai_n364_), .Y(mai_mai_n1000_));
  NA3        m0972(.A(mai_mai_n1000_), .B(mai_mai_n999_), .C(mai_mai_n998_), .Y(mai_mai_n1001_));
  OR3        m0973(.A(mai_mai_n1001_), .B(mai_mai_n997_), .C(mai_mai_n992_), .Y(mai_mai_n1002_));
  NO4        m0974(.A(mai_mai_n1002_), .B(mai_mai_n991_), .C(mai_mai_n986_), .D(mai_mai_n983_), .Y(mai_mai_n1003_));
  NA4        m0975(.A(mai_mai_n1003_), .B(mai_mai_n976_), .C(mai_mai_n943_), .D(mai_mai_n927_), .Y(mai13));
  NA2        m0976(.A(mai_mai_n46_), .B(mai_mai_n84_), .Y(mai_mai_n1005_));
  AN2        m0977(.A(c), .B(b), .Y(mai_mai_n1006_));
  NA3        m0978(.A(mai_mai_n236_), .B(mai_mai_n1006_), .C(m), .Y(mai_mai_n1007_));
  NA2        m0979(.A(mai_mai_n487_), .B(f), .Y(mai_mai_n1008_));
  NO4        m0980(.A(mai_mai_n1008_), .B(mai_mai_n1007_), .C(mai_mai_n1005_), .D(mai_mai_n571_), .Y(mai_mai_n1009_));
  NA2        m0981(.A(mai_mai_n250_), .B(mai_mai_n1006_), .Y(mai_mai_n1010_));
  NO3        m0982(.A(mai_mai_n1010_), .B(mai_mai_n1008_), .C(mai_mai_n945_), .Y(mai_mai_n1011_));
  NAi32      m0983(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1012_));
  NA2        m0984(.A(mai_mai_n129_), .B(mai_mai_n45_), .Y(mai_mai_n1013_));
  NO4        m0985(.A(mai_mai_n1013_), .B(mai_mai_n1012_), .C(mai_mai_n578_), .D(mai_mai_n292_), .Y(mai_mai_n1014_));
  NA2        m0986(.A(mai_mai_n651_), .B(mai_mai_n212_), .Y(mai_mai_n1015_));
  NA2        m0987(.A(mai_mai_n397_), .B(mai_mai_n202_), .Y(mai_mai_n1016_));
  AN2        m0988(.A(d), .B(c), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n1017_), .B(mai_mai_n109_), .Y(mai_mai_n1018_));
  NO4        m0990(.A(mai_mai_n1018_), .B(mai_mai_n1016_), .C(mai_mai_n163_), .D(mai_mai_n154_), .Y(mai_mai_n1019_));
  NA2        m0991(.A(mai_mai_n487_), .B(c), .Y(mai_mai_n1020_));
  NO4        m0992(.A(mai_mai_n1013_), .B(mai_mai_n574_), .C(mai_mai_n1020_), .D(mai_mai_n292_), .Y(mai_mai_n1021_));
  AO210      m0993(.A0(mai_mai_n1019_), .A1(mai_mai_n1015_), .B0(mai_mai_n1021_), .Y(mai_mai_n1022_));
  OR4        m0994(.A(mai_mai_n1022_), .B(mai_mai_n1014_), .C(mai_mai_n1011_), .D(mai_mai_n1009_), .Y(mai_mai_n1023_));
  NAi32      m0995(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1024_));
  NO2        m0996(.A(mai_mai_n1024_), .B(mai_mai_n133_), .Y(mai_mai_n1025_));
  NA2        m0997(.A(mai_mai_n1025_), .B(g), .Y(mai_mai_n1026_));
  OR3        m0998(.A(mai_mai_n212_), .B(mai_mai_n163_), .C(mai_mai_n154_), .Y(mai_mai_n1027_));
  NO2        m0999(.A(mai_mai_n1027_), .B(mai_mai_n1026_), .Y(mai_mai_n1028_));
  NO2        m1000(.A(mai_mai_n1020_), .B(mai_mai_n292_), .Y(mai_mai_n1029_));
  NO2        m1001(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1030_));
  NA2        m1002(.A(mai_mai_n618_), .B(mai_mai_n1030_), .Y(mai_mai_n1031_));
  NOi21      m1003(.An(mai_mai_n1029_), .B(mai_mai_n1031_), .Y(mai_mai_n1032_));
  NO2        m1004(.A(mai_mai_n743_), .B(mai_mai_n105_), .Y(mai_mai_n1033_));
  NOi41      m1005(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1034_));
  NA2        m1006(.A(mai_mai_n1034_), .B(mai_mai_n1033_), .Y(mai_mai_n1035_));
  NO2        m1007(.A(mai_mai_n1035_), .B(mai_mai_n1026_), .Y(mai_mai_n1036_));
  OR3        m1008(.A(e), .B(d), .C(c), .Y(mai_mai_n1037_));
  NA3        m1009(.A(k), .B(j), .C(i), .Y(mai_mai_n1038_));
  NO3        m1010(.A(mai_mai_n1038_), .B(mai_mai_n292_), .C(mai_mai_n87_), .Y(mai_mai_n1039_));
  NOi21      m1011(.An(mai_mai_n1039_), .B(mai_mai_n1037_), .Y(mai_mai_n1040_));
  OR4        m1012(.A(mai_mai_n1040_), .B(mai_mai_n1036_), .C(mai_mai_n1032_), .D(mai_mai_n1028_), .Y(mai_mai_n1041_));
  NA3        m1013(.A(mai_mai_n457_), .B(mai_mai_n320_), .C(mai_mai_n56_), .Y(mai_mai_n1042_));
  NO2        m1014(.A(mai_mai_n1042_), .B(mai_mai_n1031_), .Y(mai_mai_n1043_));
  NO3        m1015(.A(mai_mai_n1042_), .B(mai_mai_n574_), .C(mai_mai_n438_), .Y(mai_mai_n1044_));
  NO2        m1016(.A(f), .B(c), .Y(mai_mai_n1045_));
  NOi21      m1017(.An(mai_mai_n1045_), .B(mai_mai_n430_), .Y(mai_mai_n1046_));
  NA2        m1018(.A(mai_mai_n1046_), .B(mai_mai_n59_), .Y(mai_mai_n1047_));
  OR2        m1019(.A(k), .B(i), .Y(mai_mai_n1048_));
  NO3        m1020(.A(mai_mai_n1048_), .B(mai_mai_n232_), .C(l), .Y(mai_mai_n1049_));
  NOi31      m1021(.An(mai_mai_n1049_), .B(mai_mai_n1047_), .C(j), .Y(mai_mai_n1050_));
  OR3        m1022(.A(mai_mai_n1050_), .B(mai_mai_n1044_), .C(mai_mai_n1043_), .Y(mai_mai_n1051_));
  OR3        m1023(.A(mai_mai_n1051_), .B(mai_mai_n1041_), .C(mai_mai_n1023_), .Y(mai02));
  OR2        m1024(.A(l), .B(k), .Y(mai_mai_n1053_));
  OR3        m1025(.A(h), .B(g), .C(f), .Y(mai_mai_n1054_));
  OR3        m1026(.A(n), .B(m), .C(i), .Y(mai_mai_n1055_));
  NO4        m1027(.A(mai_mai_n1055_), .B(mai_mai_n1054_), .C(mai_mai_n1053_), .D(mai_mai_n1037_), .Y(mai_mai_n1056_));
  NOi31      m1028(.An(e), .B(d), .C(c), .Y(mai_mai_n1057_));
  AOI210     m1029(.A0(mai_mai_n1039_), .A1(mai_mai_n1057_), .B0(mai_mai_n1014_), .Y(mai_mai_n1058_));
  AN3        m1030(.A(g), .B(f), .C(c), .Y(mai_mai_n1059_));
  NA3        m1031(.A(mai_mai_n1059_), .B(mai_mai_n457_), .C(h), .Y(mai_mai_n1060_));
  OR2        m1032(.A(mai_mai_n1038_), .B(mai_mai_n292_), .Y(mai_mai_n1061_));
  OR2        m1033(.A(mai_mai_n1061_), .B(mai_mai_n1060_), .Y(mai_mai_n1062_));
  NO3        m1034(.A(mai_mai_n1042_), .B(mai_mai_n1013_), .C(mai_mai_n574_), .Y(mai_mai_n1063_));
  NO2        m1035(.A(mai_mai_n1063_), .B(mai_mai_n1028_), .Y(mai_mai_n1064_));
  NA3        m1036(.A(l), .B(k), .C(j), .Y(mai_mai_n1065_));
  NA2        m1037(.A(i), .B(h), .Y(mai_mai_n1066_));
  NO3        m1038(.A(mai_mai_n1066_), .B(mai_mai_n1065_), .C(mai_mai_n123_), .Y(mai_mai_n1067_));
  NO3        m1039(.A(mai_mai_n131_), .B(mai_mai_n268_), .C(mai_mai_n203_), .Y(mai_mai_n1068_));
  AOI210     m1040(.A0(mai_mai_n1068_), .A1(mai_mai_n1067_), .B0(mai_mai_n1032_), .Y(mai_mai_n1069_));
  NA3        m1041(.A(c), .B(b), .C(a), .Y(mai_mai_n1070_));
  NO3        m1042(.A(mai_mai_n1070_), .B(mai_mai_n877_), .C(mai_mai_n202_), .Y(mai_mai_n1071_));
  NO4        m1043(.A(mai_mai_n1038_), .B(mai_mai_n286_), .C(mai_mai_n49_), .D(mai_mai_n105_), .Y(mai_mai_n1072_));
  AOI210     m1044(.A0(mai_mai_n1072_), .A1(mai_mai_n1071_), .B0(mai_mai_n1043_), .Y(mai_mai_n1073_));
  AN4        m1045(.A(mai_mai_n1073_), .B(mai_mai_n1069_), .C(mai_mai_n1064_), .D(mai_mai_n1062_), .Y(mai_mai_n1074_));
  NO2        m1046(.A(mai_mai_n1018_), .B(mai_mai_n1016_), .Y(mai_mai_n1075_));
  NA2        m1047(.A(mai_mai_n1035_), .B(mai_mai_n1027_), .Y(mai_mai_n1076_));
  AOI210     m1048(.A0(mai_mai_n1076_), .A1(mai_mai_n1075_), .B0(mai_mai_n1009_), .Y(mai_mai_n1077_));
  NAi41      m1049(.An(mai_mai_n1056_), .B(mai_mai_n1077_), .C(mai_mai_n1074_), .D(mai_mai_n1058_), .Y(mai03));
  INV        m1050(.A(mai_mai_n355_), .Y(mai_mai_n1079_));
  NO2        m1051(.A(mai_mai_n1079_), .B(mai_mai_n970_), .Y(mai_mai_n1080_));
  NO2        m1052(.A(mai_mai_n828_), .B(mai_mai_n817_), .Y(mai_mai_n1081_));
  OAI220     m1053(.A0(mai_mai_n1081_), .A1(mai_mai_n673_), .B0(mai_mai_n1080_), .B1(mai_mai_n575_), .Y(mai_mai_n1082_));
  NOi31      m1054(.An(i), .B(k), .C(j), .Y(mai_mai_n1083_));
  NA4        m1055(.A(mai_mai_n1083_), .B(mai_mai_n1057_), .C(mai_mai_n329_), .D(mai_mai_n320_), .Y(mai_mai_n1084_));
  OAI210     m1056(.A0(mai_mai_n794_), .A1(mai_mai_n407_), .B0(mai_mai_n1084_), .Y(mai_mai_n1085_));
  NOi31      m1057(.An(m), .B(n), .C(f), .Y(mai_mai_n1086_));
  NA2        m1058(.A(mai_mai_n1086_), .B(mai_mai_n51_), .Y(mai_mai_n1087_));
  AN2        m1059(.A(e), .B(c), .Y(mai_mai_n1088_));
  NA2        m1060(.A(mai_mai_n1088_), .B(a), .Y(mai_mai_n1089_));
  OAI220     m1061(.A0(mai_mai_n1089_), .A1(mai_mai_n1087_), .B0(mai_mai_n861_), .B1(mai_mai_n413_), .Y(mai_mai_n1090_));
  NA2        m1062(.A(mai_mai_n497_), .B(l), .Y(mai_mai_n1091_));
  NOi31      m1063(.An(mai_mai_n839_), .B(mai_mai_n1007_), .C(mai_mai_n1091_), .Y(mai_mai_n1092_));
  NO4        m1064(.A(mai_mai_n1092_), .B(mai_mai_n1090_), .C(mai_mai_n1085_), .D(mai_mai_n969_), .Y(mai_mai_n1093_));
  NO2        m1065(.A(mai_mai_n268_), .B(a), .Y(mai_mai_n1094_));
  INV        m1066(.A(mai_mai_n1014_), .Y(mai_mai_n1095_));
  NO2        m1067(.A(mai_mai_n1066_), .B(mai_mai_n477_), .Y(mai_mai_n1096_));
  NO2        m1068(.A(mai_mai_n84_), .B(g), .Y(mai_mai_n1097_));
  AOI210     m1069(.A0(mai_mai_n1097_), .A1(mai_mai_n1096_), .B0(mai_mai_n1049_), .Y(mai_mai_n1098_));
  OR2        m1070(.A(mai_mai_n1098_), .B(mai_mai_n1047_), .Y(mai_mai_n1099_));
  NA3        m1071(.A(mai_mai_n1099_), .B(mai_mai_n1095_), .C(mai_mai_n1093_), .Y(mai_mai_n1100_));
  NO4        m1072(.A(mai_mai_n1100_), .B(mai_mai_n1082_), .C(mai_mai_n795_), .D(mai_mai_n557_), .Y(mai_mai_n1101_));
  NA2        m1073(.A(c), .B(b), .Y(mai_mai_n1102_));
  NO2        m1074(.A(mai_mai_n685_), .B(mai_mai_n1102_), .Y(mai_mai_n1103_));
  OAI210     m1075(.A0(mai_mai_n837_), .A1(mai_mai_n810_), .B0(mai_mai_n400_), .Y(mai_mai_n1104_));
  OAI210     m1076(.A0(mai_mai_n1104_), .A1(mai_mai_n838_), .B0(mai_mai_n1103_), .Y(mai_mai_n1105_));
  NAi21      m1077(.An(mai_mai_n408_), .B(mai_mai_n1103_), .Y(mai_mai_n1106_));
  NA3        m1078(.A(mai_mai_n414_), .B(mai_mai_n550_), .C(f), .Y(mai_mai_n1107_));
  OAI210     m1079(.A0(mai_mai_n539_), .A1(mai_mai_n39_), .B0(mai_mai_n1094_), .Y(mai_mai_n1108_));
  NA3        m1080(.A(mai_mai_n1108_), .B(mai_mai_n1107_), .C(mai_mai_n1106_), .Y(mai_mai_n1109_));
  INV        m1081(.A(mai_mai_n247_), .Y(mai_mai_n1110_));
  OAI210     m1082(.A0(mai_mai_n1110_), .A1(mai_mai_n272_), .B0(g), .Y(mai_mai_n1111_));
  NAi21      m1083(.An(f), .B(d), .Y(mai_mai_n1112_));
  NO2        m1084(.A(mai_mai_n1112_), .B(mai_mai_n1070_), .Y(mai_mai_n1113_));
  INV        m1085(.A(mai_mai_n1113_), .Y(mai_mai_n1114_));
  AOI210     m1086(.A0(mai_mai_n1111_), .A1(mai_mai_n278_), .B0(mai_mai_n1114_), .Y(mai_mai_n1115_));
  AOI210     m1087(.A0(mai_mai_n1115_), .A1(mai_mai_n106_), .B0(mai_mai_n1109_), .Y(mai_mai_n1116_));
  NA2        m1088(.A(mai_mai_n460_), .B(mai_mai_n459_), .Y(mai_mai_n1117_));
  NO2        m1089(.A(mai_mai_n169_), .B(mai_mai_n225_), .Y(mai_mai_n1118_));
  NA2        m1090(.A(mai_mai_n1118_), .B(m), .Y(mai_mai_n1119_));
  NA3        m1091(.A(mai_mai_n894_), .B(mai_mai_n1091_), .C(mai_mai_n463_), .Y(mai_mai_n1120_));
  OAI210     m1092(.A0(mai_mai_n1120_), .A1(mai_mai_n297_), .B0(mai_mai_n461_), .Y(mai_mai_n1121_));
  AOI210     m1093(.A0(mai_mai_n1121_), .A1(mai_mai_n1117_), .B0(mai_mai_n1119_), .Y(mai_mai_n1122_));
  NA2        m1094(.A(mai_mai_n552_), .B(mai_mai_n396_), .Y(mai_mai_n1123_));
  NA2        m1095(.A(mai_mai_n145_), .B(mai_mai_n33_), .Y(mai_mai_n1124_));
  AOI210     m1096(.A0(mai_mai_n941_), .A1(mai_mai_n1124_), .B0(mai_mai_n203_), .Y(mai_mai_n1125_));
  OAI210     m1097(.A0(mai_mai_n1125_), .A1(mai_mai_n434_), .B0(mai_mai_n1113_), .Y(mai_mai_n1126_));
  AOI210     m1098(.A0(mai_mai_n1118_), .A1(mai_mai_n416_), .B0(mai_mai_n935_), .Y(mai_mai_n1127_));
  NA3        m1099(.A(mai_mai_n1127_), .B(mai_mai_n1126_), .C(mai_mai_n1123_), .Y(mai_mai_n1128_));
  NO2        m1100(.A(mai_mai_n1128_), .B(mai_mai_n1122_), .Y(mai_mai_n1129_));
  NA4        m1101(.A(mai_mai_n1129_), .B(mai_mai_n1116_), .C(mai_mai_n1105_), .D(mai_mai_n1101_), .Y(mai00));
  AOI210     m1102(.A0(mai_mai_n285_), .A1(mai_mai_n203_), .B0(mai_mai_n260_), .Y(mai_mai_n1131_));
  NO2        m1103(.A(mai_mai_n1131_), .B(mai_mai_n565_), .Y(mai_mai_n1132_));
  AOI210     m1104(.A0(mai_mai_n874_), .A1(mai_mai_n920_), .B0(mai_mai_n1085_), .Y(mai_mai_n1133_));
  NO2        m1105(.A(mai_mai_n1063_), .B(mai_mai_n935_), .Y(mai_mai_n1134_));
  NA3        m1106(.A(mai_mai_n1134_), .B(mai_mai_n1133_), .C(mai_mai_n971_), .Y(mai_mai_n1135_));
  NA2        m1107(.A(mai_mai_n499_), .B(f), .Y(mai_mai_n1136_));
  OAI210     m1108(.A0(mai_mai_n978_), .A1(mai_mai_n40_), .B0(mai_mai_n630_), .Y(mai_mai_n1137_));
  NA3        m1109(.A(mai_mai_n1137_), .B(mai_mai_n243_), .C(n), .Y(mai_mai_n1138_));
  AOI210     m1110(.A0(mai_mai_n1138_), .A1(mai_mai_n1136_), .B0(mai_mai_n1018_), .Y(mai_mai_n1139_));
  NO4        m1111(.A(mai_mai_n1139_), .B(mai_mai_n1135_), .C(mai_mai_n1132_), .D(mai_mai_n1041_), .Y(mai_mai_n1140_));
  NA3        m1112(.A(mai_mai_n153_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1141_));
  NA3        m1113(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1142_));
  NOi31      m1114(.An(n), .B(m), .C(i), .Y(mai_mai_n1143_));
  NA3        m1115(.A(mai_mai_n1143_), .B(mai_mai_n633_), .C(mai_mai_n51_), .Y(mai_mai_n1144_));
  OAI210     m1116(.A0(mai_mai_n1142_), .A1(mai_mai_n1141_), .B0(mai_mai_n1144_), .Y(mai_mai_n1145_));
  INV        m1117(.A(mai_mai_n564_), .Y(mai_mai_n1146_));
  NO3        m1118(.A(mai_mai_n1146_), .B(mai_mai_n1145_), .C(mai_mai_n897_), .Y(mai_mai_n1147_));
  NA3        m1119(.A(mai_mai_n369_), .B(mai_mai_n208_), .C(g), .Y(mai_mai_n1148_));
  OR2        m1120(.A(mai_mai_n1148_), .B(mai_mai_n1142_), .Y(mai_mai_n1149_));
  NO2        m1121(.A(h), .B(g), .Y(mai_mai_n1150_));
  NA4        m1122(.A(mai_mai_n489_), .B(mai_mai_n457_), .C(mai_mai_n1150_), .D(mai_mai_n1006_), .Y(mai_mai_n1151_));
  NA2        m1123(.A(mai_mai_n923_), .B(mai_mai_n563_), .Y(mai_mai_n1152_));
  NA3        m1124(.A(mai_mai_n1152_), .B(mai_mai_n1151_), .C(mai_mai_n1149_), .Y(mai_mai_n1153_));
  NO2        m1125(.A(mai_mai_n1153_), .B(mai_mai_n251_), .Y(mai_mai_n1154_));
  NO2        m1126(.A(mai_mai_n227_), .B(mai_mai_n168_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n1155_), .B(mai_mai_n414_), .Y(mai_mai_n1156_));
  NA3        m1128(.A(mai_mai_n166_), .B(mai_mai_n105_), .C(g), .Y(mai_mai_n1157_));
  NA3        m1129(.A(mai_mai_n457_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1158_));
  NOi31      m1130(.An(mai_mai_n847_), .B(mai_mai_n1158_), .C(mai_mai_n1157_), .Y(mai_mai_n1159_));
  NAi31      m1131(.An(mai_mai_n173_), .B(mai_mai_n834_), .C(mai_mai_n457_), .Y(mai_mai_n1160_));
  NAi31      m1132(.An(mai_mai_n1159_), .B(mai_mai_n1160_), .C(mai_mai_n1156_), .Y(mai_mai_n1161_));
  NO2        m1133(.A(mai_mai_n259_), .B(mai_mai_n74_), .Y(mai_mai_n1162_));
  NO3        m1134(.A(mai_mai_n413_), .B(mai_mai_n806_), .C(n), .Y(mai_mai_n1163_));
  AOI210     m1135(.A0(mai_mai_n1163_), .A1(mai_mai_n1162_), .B0(mai_mai_n1056_), .Y(mai_mai_n1164_));
  NAi31      m1136(.An(mai_mai_n1021_), .B(mai_mai_n1164_), .C(mai_mai_n73_), .Y(mai_mai_n1165_));
  NO4        m1137(.A(mai_mai_n1165_), .B(mai_mai_n1161_), .C(mai_mai_n566_), .D(mai_mai_n509_), .Y(mai_mai_n1166_));
  AN3        m1138(.A(mai_mai_n1166_), .B(mai_mai_n1154_), .C(mai_mai_n1147_), .Y(mai_mai_n1167_));
  NA3        m1139(.A(mai_mai_n1086_), .B(mai_mai_n597_), .C(mai_mai_n456_), .Y(mai_mai_n1168_));
  NA3        m1140(.A(mai_mai_n1168_), .B(mai_mai_n553_), .C(mai_mai_n230_), .Y(mai_mai_n1169_));
  NA2        m1141(.A(mai_mai_n1079_), .B(mai_mai_n526_), .Y(mai_mai_n1170_));
  NA4        m1142(.A(mai_mai_n633_), .B(mai_mai_n194_), .C(mai_mai_n208_), .D(mai_mai_n149_), .Y(mai_mai_n1171_));
  NA3        m1143(.A(mai_mai_n1171_), .B(mai_mai_n1170_), .C(mai_mai_n282_), .Y(mai_mai_n1172_));
  OAI210     m1144(.A0(mai_mai_n455_), .A1(mai_mai_n113_), .B0(mai_mai_n840_), .Y(mai_mai_n1173_));
  AOI220     m1145(.A0(mai_mai_n1173_), .A1(mai_mai_n1120_), .B0(mai_mai_n552_), .B1(mai_mai_n396_), .Y(mai_mai_n1174_));
  OR4        m1146(.A(mai_mai_n1018_), .B(mai_mai_n257_), .C(mai_mai_n210_), .D(e), .Y(mai_mai_n1175_));
  NO2        m1147(.A(mai_mai_n206_), .B(mai_mai_n203_), .Y(mai_mai_n1176_));
  NA2        m1148(.A(n), .B(e), .Y(mai_mai_n1177_));
  NO2        m1149(.A(mai_mai_n1177_), .B(mai_mai_n133_), .Y(mai_mai_n1178_));
  AOI220     m1150(.A0(mai_mai_n1178_), .A1(mai_mai_n258_), .B0(mai_mai_n821_), .B1(mai_mai_n1176_), .Y(mai_mai_n1179_));
  NA3        m1151(.A(mai_mai_n1179_), .B(mai_mai_n1175_), .C(mai_mai_n1174_), .Y(mai_mai_n1180_));
  AOI210     m1152(.A0(mai_mai_n1178_), .A1(mai_mai_n825_), .B0(mai_mai_n795_), .Y(mai_mai_n1181_));
  AOI220     m1153(.A0(mai_mai_n931_), .A1(mai_mai_n563_), .B0(mai_mai_n633_), .B1(mai_mai_n233_), .Y(mai_mai_n1182_));
  NO2        m1154(.A(mai_mai_n68_), .B(h), .Y(mai_mai_n1183_));
  NO3        m1155(.A(mai_mai_n1018_), .B(mai_mai_n1016_), .C(mai_mai_n707_), .Y(mai_mai_n1184_));
  NO2        m1156(.A(mai_mai_n1053_), .B(mai_mai_n123_), .Y(mai_mai_n1185_));
  AN2        m1157(.A(mai_mai_n1185_), .B(mai_mai_n1068_), .Y(mai_mai_n1186_));
  OAI210     m1158(.A0(mai_mai_n1186_), .A1(mai_mai_n1184_), .B0(mai_mai_n1183_), .Y(mai_mai_n1187_));
  NA4        m1159(.A(mai_mai_n1187_), .B(mai_mai_n1182_), .C(mai_mai_n1181_), .D(mai_mai_n842_), .Y(mai_mai_n1188_));
  NO4        m1160(.A(mai_mai_n1188_), .B(mai_mai_n1180_), .C(mai_mai_n1172_), .D(mai_mai_n1169_), .Y(mai_mai_n1189_));
  NA2        m1161(.A(mai_mai_n811_), .B(mai_mai_n738_), .Y(mai_mai_n1190_));
  NA4        m1162(.A(mai_mai_n1190_), .B(mai_mai_n1189_), .C(mai_mai_n1167_), .D(mai_mai_n1140_), .Y(mai01));
  AN2        m1163(.A(mai_mai_n995_), .B(mai_mai_n993_), .Y(mai_mai_n1192_));
  NO4        m1164(.A(mai_mai_n782_), .B(mai_mai_n774_), .C(mai_mai_n471_), .D(mai_mai_n266_), .Y(mai_mai_n1193_));
  NA2        m1165(.A(mai_mai_n380_), .B(i), .Y(mai_mai_n1194_));
  NA3        m1166(.A(mai_mai_n1194_), .B(mai_mai_n1193_), .C(mai_mai_n1192_), .Y(mai_mai_n1195_));
  NA2        m1167(.A(mai_mai_n545_), .B(mai_mai_n256_), .Y(mai_mai_n1196_));
  NA2        m1168(.A(mai_mai_n938_), .B(mai_mai_n1196_), .Y(mai_mai_n1197_));
  NA3        m1169(.A(mai_mai_n1197_), .B(mai_mai_n890_), .C(mai_mai_n319_), .Y(mai_mai_n1198_));
  NA2        m1170(.A(mai_mai_n45_), .B(f), .Y(mai_mai_n1199_));
  NA2        m1171(.A(mai_mai_n692_), .B(mai_mai_n91_), .Y(mai_mai_n1200_));
  NO2        m1172(.A(mai_mai_n1200_), .B(mai_mai_n1199_), .Y(mai_mai_n1201_));
  INV        m1173(.A(mai_mai_n111_), .Y(mai_mai_n1202_));
  OA220      m1174(.A0(mai_mai_n1202_), .A1(mai_mai_n573_), .B0(mai_mai_n645_), .B1(mai_mai_n355_), .Y(mai_mai_n1203_));
  NAi41      m1175(.An(mai_mai_n148_), .B(mai_mai_n1203_), .C(mai_mai_n1171_), .D(mai_mai_n873_), .Y(mai_mai_n1204_));
  NO3        m1176(.A(mai_mai_n763_), .B(mai_mai_n657_), .C(mai_mai_n502_), .Y(mai_mai_n1205_));
  OR2        m1177(.A(mai_mai_n183_), .B(mai_mai_n181_), .Y(mai_mai_n1206_));
  NA3        m1178(.A(mai_mai_n1206_), .B(mai_mai_n1205_), .C(mai_mai_n127_), .Y(mai_mai_n1207_));
  NO4        m1179(.A(mai_mai_n1207_), .B(mai_mai_n1204_), .C(mai_mai_n1198_), .D(mai_mai_n1195_), .Y(mai_mai_n1208_));
  INV        m1180(.A(mai_mai_n1148_), .Y(mai_mai_n1209_));
  NA2        m1181(.A(mai_mai_n1209_), .B(mai_mai_n522_), .Y(mai_mai_n1210_));
  NA2        m1182(.A(mai_mai_n528_), .B(mai_mai_n382_), .Y(mai_mai_n1211_));
  NOi21      m1183(.An(mai_mai_n554_), .B(mai_mai_n570_), .Y(mai_mai_n1212_));
  NA2        m1184(.A(mai_mai_n1212_), .B(mai_mai_n1211_), .Y(mai_mai_n1213_));
  AOI210     m1185(.A0(mai_mai_n192_), .A1(mai_mai_n86_), .B0(mai_mai_n202_), .Y(mai_mai_n1214_));
  OAI210     m1186(.A0(mai_mai_n788_), .A1(mai_mai_n414_), .B0(mai_mai_n1214_), .Y(mai_mai_n1215_));
  NA2        m1187(.A(mai_mai_n191_), .B(mai_mai_n34_), .Y(mai_mai_n1216_));
  OR2        m1188(.A(mai_mai_n1216_), .B(mai_mai_n318_), .Y(mai_mai_n1217_));
  NA4        m1189(.A(mai_mai_n1217_), .B(mai_mai_n1215_), .C(mai_mai_n1213_), .D(mai_mai_n1210_), .Y(mai_mai_n1218_));
  AOI210     m1190(.A0(mai_mai_n585_), .A1(mai_mai_n111_), .B0(mai_mai_n591_), .Y(mai_mai_n1219_));
  OAI210     m1191(.A0(mai_mai_n1202_), .A1(mai_mai_n582_), .B0(mai_mai_n1219_), .Y(mai_mai_n1220_));
  NA2        m1192(.A(mai_mai_n265_), .B(mai_mai_n183_), .Y(mai_mai_n1221_));
  NA2        m1193(.A(mai_mai_n1221_), .B(mai_mai_n650_), .Y(mai_mai_n1222_));
  NO3        m1194(.A(mai_mai_n794_), .B(mai_mai_n192_), .C(mai_mai_n394_), .Y(mai_mai_n1223_));
  NO2        m1195(.A(mai_mai_n1223_), .B(mai_mai_n935_), .Y(mai_mai_n1224_));
  OAI210     m1196(.A0(mai_mai_n1201_), .A1(mai_mai_n313_), .B0(mai_mai_n658_), .Y(mai_mai_n1225_));
  NA4        m1197(.A(mai_mai_n1225_), .B(mai_mai_n1224_), .C(mai_mai_n1222_), .D(mai_mai_n766_), .Y(mai_mai_n1226_));
  NO3        m1198(.A(mai_mai_n1226_), .B(mai_mai_n1220_), .C(mai_mai_n1218_), .Y(mai_mai_n1227_));
  NA3        m1199(.A(mai_mai_n593_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1228_));
  NO2        m1200(.A(mai_mai_n1228_), .B(mai_mai_n192_), .Y(mai_mai_n1229_));
  AOI210     m1201(.A0(mai_mai_n495_), .A1(mai_mai_n58_), .B0(mai_mai_n1229_), .Y(mai_mai_n1230_));
  OR3        m1202(.A(mai_mai_n1200_), .B(mai_mai_n594_), .C(mai_mai_n1199_), .Y(mai_mai_n1231_));
  NO2        m1203(.A(mai_mai_n195_), .B(mai_mai_n104_), .Y(mai_mai_n1232_));
  NO2        m1204(.A(mai_mai_n1232_), .B(mai_mai_n1145_), .Y(mai_mai_n1233_));
  NA4        m1205(.A(mai_mai_n1233_), .B(mai_mai_n1231_), .C(mai_mai_n1230_), .D(mai_mai_n737_), .Y(mai_mai_n1234_));
  NO2        m1206(.A(mai_mai_n945_), .B(mai_mai_n220_), .Y(mai_mai_n1235_));
  NO2        m1207(.A(mai_mai_n946_), .B(mai_mai_n547_), .Y(mai_mai_n1236_));
  OAI210     m1208(.A0(mai_mai_n1236_), .A1(mai_mai_n1235_), .B0(mai_mai_n327_), .Y(mai_mai_n1237_));
  NO3        m1209(.A(mai_mai_n78_), .B(mai_mai_n286_), .C(mai_mai_n45_), .Y(mai_mai_n1238_));
  OR2        m1210(.A(mai_mai_n1148_), .B(mai_mai_n1142_), .Y(mai_mai_n1239_));
  NO2        m1211(.A(mai_mai_n355_), .B(mai_mai_n72_), .Y(mai_mai_n1240_));
  INV        m1212(.A(mai_mai_n1240_), .Y(mai_mai_n1241_));
  NA2        m1213(.A(mai_mai_n1238_), .B(mai_mai_n789_), .Y(mai_mai_n1242_));
  NA4        m1214(.A(mai_mai_n1242_), .B(mai_mai_n1241_), .C(mai_mai_n1239_), .D(mai_mai_n372_), .Y(mai_mai_n1243_));
  NOi31      m1215(.An(mai_mai_n1237_), .B(mai_mai_n1243_), .C(mai_mai_n1234_), .Y(mai_mai_n1244_));
  NO2        m1216(.A(mai_mai_n122_), .B(mai_mai_n45_), .Y(mai_mai_n1245_));
  NO2        m1217(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1246_));
  AO220      m1218(.A0(mai_mai_n1246_), .A1(mai_mai_n613_), .B0(mai_mai_n1245_), .B1(mai_mai_n690_), .Y(mai_mai_n1247_));
  NA2        m1219(.A(mai_mai_n1247_), .B(mai_mai_n327_), .Y(mai_mai_n1248_));
  NO3        m1220(.A(mai_mai_n1066_), .B(mai_mai_n163_), .C(mai_mai_n84_), .Y(mai_mai_n1249_));
  NA2        m1221(.A(mai_mai_n1238_), .B(mai_mai_n949_), .Y(mai_mai_n1250_));
  NA2        m1222(.A(mai_mai_n1250_), .B(mai_mai_n1248_), .Y(mai_mai_n1251_));
  NO2        m1223(.A(mai_mai_n605_), .B(mai_mai_n604_), .Y(mai_mai_n1252_));
  NO4        m1224(.A(mai_mai_n1066_), .B(mai_mai_n1252_), .C(mai_mai_n161_), .D(mai_mai_n84_), .Y(mai_mai_n1253_));
  NO3        m1225(.A(mai_mai_n1253_), .B(mai_mai_n1251_), .C(mai_mai_n624_), .Y(mai_mai_n1254_));
  NA4        m1226(.A(mai_mai_n1254_), .B(mai_mai_n1244_), .C(mai_mai_n1227_), .D(mai_mai_n1208_), .Y(mai06));
  NO2        m1227(.A(mai_mai_n395_), .B(mai_mai_n551_), .Y(mai_mai_n1256_));
  INV        m1228(.A(mai_mai_n714_), .Y(mai_mai_n1257_));
  OAI210     m1229(.A0(mai_mai_n1257_), .A1(mai_mai_n252_), .B0(mai_mai_n1256_), .Y(mai_mai_n1258_));
  NO2        m1230(.A(mai_mai_n212_), .B(mai_mai_n95_), .Y(mai_mai_n1259_));
  OAI210     m1231(.A0(mai_mai_n1259_), .A1(mai_mai_n1249_), .B0(mai_mai_n368_), .Y(mai_mai_n1260_));
  NO3        m1232(.A(mai_mai_n589_), .B(mai_mai_n786_), .C(mai_mai_n592_), .Y(mai_mai_n1261_));
  OR2        m1233(.A(mai_mai_n1261_), .B(mai_mai_n861_), .Y(mai_mai_n1262_));
  NA4        m1234(.A(mai_mai_n1262_), .B(mai_mai_n1260_), .C(mai_mai_n1258_), .D(mai_mai_n1237_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(mai_mai_n1263_), .B(mai_mai_n242_), .Y(mai_mai_n1264_));
  NO2        m1236(.A(mai_mai_n286_), .B(mai_mai_n45_), .Y(mai_mai_n1265_));
  AOI210     m1237(.A0(mai_mai_n1265_), .A1(mai_mai_n950_), .B0(mai_mai_n1235_), .Y(mai_mai_n1266_));
  AOI210     m1238(.A0(mai_mai_n1265_), .A1(mai_mai_n548_), .B0(mai_mai_n1247_), .Y(mai_mai_n1267_));
  AOI210     m1239(.A0(mai_mai_n1267_), .A1(mai_mai_n1266_), .B0(mai_mai_n324_), .Y(mai_mai_n1268_));
  OAI210     m1240(.A0(mai_mai_n86_), .A1(mai_mai_n40_), .B0(mai_mai_n656_), .Y(mai_mai_n1269_));
  NA2        m1241(.A(mai_mai_n1269_), .B(mai_mai_n627_), .Y(mai_mai_n1270_));
  NO2        m1242(.A(mai_mai_n505_), .B(mai_mai_n158_), .Y(mai_mai_n1271_));
  NO2        m1243(.A(mai_mai_n598_), .B(mai_mai_n1087_), .Y(mai_mai_n1272_));
  OAI210     m1244(.A0(mai_mai_n450_), .A1(mai_mai_n235_), .B0(mai_mai_n884_), .Y(mai_mai_n1273_));
  NO3        m1245(.A(mai_mai_n1273_), .B(mai_mai_n1272_), .C(mai_mai_n1271_), .Y(mai_mai_n1274_));
  OR2        m1246(.A(mai_mai_n590_), .B(mai_mai_n588_), .Y(mai_mai_n1275_));
  NO2        m1247(.A(mai_mai_n354_), .B(mai_mai_n126_), .Y(mai_mai_n1276_));
  AOI210     m1248(.A0(mai_mai_n1276_), .A1(mai_mai_n576_), .B0(mai_mai_n1275_), .Y(mai_mai_n1277_));
  NA3        m1249(.A(mai_mai_n1277_), .B(mai_mai_n1274_), .C(mai_mai_n1270_), .Y(mai_mai_n1278_));
  NO2        m1250(.A(mai_mai_n730_), .B(mai_mai_n353_), .Y(mai_mai_n1279_));
  NO2        m1251(.A(mai_mai_n658_), .B(mai_mai_n739_), .Y(mai_mai_n1280_));
  NOi21      m1252(.An(mai_mai_n1279_), .B(mai_mai_n1280_), .Y(mai_mai_n1281_));
  AN2        m1253(.A(mai_mai_n931_), .B(mai_mai_n629_), .Y(mai_mai_n1282_));
  NO4        m1254(.A(mai_mai_n1282_), .B(mai_mai_n1281_), .C(mai_mai_n1278_), .D(mai_mai_n1268_), .Y(mai_mai_n1283_));
  NO2        m1255(.A(mai_mai_n781_), .B(mai_mai_n261_), .Y(mai_mai_n1284_));
  OAI220     m1256(.A0(mai_mai_n714_), .A1(mai_mai_n47_), .B0(mai_mai_n212_), .B1(mai_mai_n607_), .Y(mai_mai_n1285_));
  OAI210     m1257(.A0(mai_mai_n261_), .A1(c), .B0(mai_mai_n626_), .Y(mai_mai_n1286_));
  AOI220     m1258(.A0(mai_mai_n1286_), .A1(mai_mai_n1285_), .B0(mai_mai_n1284_), .B1(mai_mai_n252_), .Y(mai_mai_n1287_));
  NO3        m1259(.A(mai_mai_n232_), .B(mai_mai_n95_), .C(mai_mai_n268_), .Y(mai_mai_n1288_));
  OAI220     m1260(.A0(mai_mai_n682_), .A1(mai_mai_n235_), .B0(mai_mai_n501_), .B1(mai_mai_n505_), .Y(mai_mai_n1289_));
  NO3        m1261(.A(mai_mai_n1289_), .B(mai_mai_n1288_), .C(mai_mai_n1090_), .Y(mai_mai_n1290_));
  NA4        m1262(.A(mai_mai_n772_), .B(mai_mai_n771_), .C(mai_mai_n424_), .D(mai_mai_n854_), .Y(mai_mai_n1291_));
  NAi31      m1263(.An(mai_mai_n730_), .B(mai_mai_n1291_), .C(mai_mai_n191_), .Y(mai_mai_n1292_));
  NA4        m1264(.A(mai_mai_n1292_), .B(mai_mai_n1290_), .C(mai_mai_n1287_), .D(mai_mai_n1182_), .Y(mai_mai_n1293_));
  NOi31      m1265(.An(mai_mai_n1261_), .B(mai_mai_n454_), .C(mai_mai_n381_), .Y(mai_mai_n1294_));
  OR3        m1266(.A(mai_mai_n1294_), .B(mai_mai_n762_), .C(mai_mai_n531_), .Y(mai_mai_n1295_));
  OR3        m1267(.A(mai_mai_n357_), .B(mai_mai_n212_), .C(mai_mai_n607_), .Y(mai_mai_n1296_));
  NA2        m1268(.A(mai_mai_n1296_), .B(mai_mai_n1295_), .Y(mai_mai_n1297_));
  AOI220     m1269(.A0(mai_mai_n1279_), .A1(mai_mai_n738_), .B0(mai_mai_n1276_), .B1(mai_mai_n226_), .Y(mai_mai_n1298_));
  AN2        m1270(.A(mai_mai_n906_), .B(mai_mai_n905_), .Y(mai_mai_n1299_));
  NO4        m1271(.A(mai_mai_n1299_), .B(mai_mai_n852_), .C(mai_mai_n491_), .D(mai_mai_n474_), .Y(mai_mai_n1300_));
  NA3        m1272(.A(mai_mai_n1300_), .B(mai_mai_n1298_), .C(mai_mai_n1242_), .Y(mai_mai_n1301_));
  NAi21      m1273(.An(j), .B(i), .Y(mai_mai_n1302_));
  NO4        m1274(.A(mai_mai_n1252_), .B(mai_mai_n1302_), .C(mai_mai_n430_), .D(mai_mai_n223_), .Y(mai_mai_n1303_));
  NO4        m1275(.A(mai_mai_n1303_), .B(mai_mai_n1301_), .C(mai_mai_n1297_), .D(mai_mai_n1293_), .Y(mai_mai_n1304_));
  NA4        m1276(.A(mai_mai_n1304_), .B(mai_mai_n1283_), .C(mai_mai_n1264_), .D(mai_mai_n1254_), .Y(mai07));
  NOi21      m1277(.An(j), .B(k), .Y(mai_mai_n1306_));
  NA4        m1278(.A(mai_mai_n166_), .B(mai_mai_n101_), .C(mai_mai_n1306_), .D(f), .Y(mai_mai_n1307_));
  NAi32      m1279(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1308_));
  NO3        m1280(.A(mai_mai_n1308_), .B(g), .C(f), .Y(mai_mai_n1309_));
  OAI210     m1281(.A0(mai_mai_n308_), .A1(mai_mai_n476_), .B0(mai_mai_n1309_), .Y(mai_mai_n1310_));
  NAi21      m1282(.An(f), .B(c), .Y(mai_mai_n1311_));
  OR2        m1283(.A(e), .B(d), .Y(mai_mai_n1312_));
  OAI220     m1284(.A0(mai_mai_n1312_), .A1(mai_mai_n1311_), .B0(mai_mai_n617_), .B1(mai_mai_n309_), .Y(mai_mai_n1313_));
  NA3        m1285(.A(mai_mai_n1313_), .B(mai_mai_n1030_), .C(mai_mai_n166_), .Y(mai_mai_n1314_));
  NOi31      m1286(.An(n), .B(m), .C(b), .Y(mai_mai_n1315_));
  NO3        m1287(.A(mai_mai_n123_), .B(mai_mai_n438_), .C(h), .Y(mai_mai_n1316_));
  NA3        m1288(.A(mai_mai_n1314_), .B(mai_mai_n1310_), .C(mai_mai_n1307_), .Y(mai_mai_n1317_));
  NOi41      m1289(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1318_));
  NA3        m1290(.A(mai_mai_n1318_), .B(mai_mai_n844_), .C(mai_mai_n397_), .Y(mai_mai_n1319_));
  NOi21      m1291(.An(h), .B(k), .Y(mai_mai_n1320_));
  NO2        m1292(.A(mai_mai_n1319_), .B(mai_mai_n56_), .Y(mai_mai_n1321_));
  NO2        m1293(.A(k), .B(i), .Y(mai_mai_n1322_));
  NA3        m1294(.A(mai_mai_n1322_), .B(mai_mai_n872_), .C(mai_mai_n166_), .Y(mai_mai_n1323_));
  NA2        m1295(.A(mai_mai_n84_), .B(mai_mai_n45_), .Y(mai_mai_n1324_));
  NO2        m1296(.A(mai_mai_n1024_), .B(mai_mai_n430_), .Y(mai_mai_n1325_));
  NA3        m1297(.A(mai_mai_n1325_), .B(mai_mai_n1324_), .C(mai_mai_n203_), .Y(mai_mai_n1326_));
  NO2        m1298(.A(mai_mai_n1038_), .B(mai_mai_n292_), .Y(mai_mai_n1327_));
  NA2        m1299(.A(mai_mai_n532_), .B(mai_mai_n79_), .Y(mai_mai_n1328_));
  NA2        m1300(.A(mai_mai_n1183_), .B(mai_mai_n276_), .Y(mai_mai_n1329_));
  NA4        m1301(.A(mai_mai_n1329_), .B(mai_mai_n1328_), .C(mai_mai_n1326_), .D(mai_mai_n1323_), .Y(mai_mai_n1330_));
  NO3        m1302(.A(mai_mai_n1330_), .B(mai_mai_n1321_), .C(mai_mai_n1317_), .Y(mai_mai_n1331_));
  NO3        m1303(.A(e), .B(d), .C(c), .Y(mai_mai_n1332_));
  NA2        m1304(.A(mai_mai_n1509_), .B(mai_mai_n1332_), .Y(mai_mai_n1333_));
  NO2        m1305(.A(mai_mai_n1333_), .B(mai_mai_n203_), .Y(mai_mai_n1334_));
  OR2        m1306(.A(h), .B(f), .Y(mai_mai_n1335_));
  NO3        m1307(.A(n), .B(m), .C(i), .Y(mai_mai_n1336_));
  OAI210     m1308(.A0(mai_mai_n1088_), .A1(mai_mai_n143_), .B0(mai_mai_n1336_), .Y(mai_mai_n1337_));
  NO2        m1309(.A(mai_mai_n1337_), .B(mai_mai_n1335_), .Y(mai_mai_n1338_));
  NA3        m1310(.A(mai_mai_n679_), .B(mai_mai_n666_), .C(mai_mai_n105_), .Y(mai_mai_n1339_));
  NO2        m1311(.A(mai_mai_n1339_), .B(mai_mai_n45_), .Y(mai_mai_n1340_));
  NO2        m1312(.A(l), .B(k), .Y(mai_mai_n1341_));
  NOi41      m1313(.An(mai_mai_n537_), .B(mai_mai_n1341_), .C(mai_mai_n469_), .D(mai_mai_n430_), .Y(mai_mai_n1342_));
  NO3        m1314(.A(mai_mai_n430_), .B(d), .C(c), .Y(mai_mai_n1343_));
  NO4        m1315(.A(mai_mai_n1342_), .B(mai_mai_n1340_), .C(mai_mai_n1338_), .D(mai_mai_n1334_), .Y(mai_mai_n1344_));
  NO2        m1316(.A(mai_mai_n134_), .B(h), .Y(mai_mai_n1345_));
  NO2        m1317(.A(mai_mai_n1048_), .B(l), .Y(mai_mai_n1346_));
  NO2        m1318(.A(g), .B(c), .Y(mai_mai_n1347_));
  NA3        m1319(.A(mai_mai_n1347_), .B(mai_mai_n131_), .C(mai_mai_n174_), .Y(mai_mai_n1348_));
  NO2        m1320(.A(mai_mai_n1348_), .B(mai_mai_n1346_), .Y(mai_mai_n1349_));
  NA2        m1321(.A(mai_mai_n1349_), .B(mai_mai_n166_), .Y(mai_mai_n1350_));
  OAI210     m1322(.A0(mai_mai_n1320_), .A1(mai_mai_n202_), .B0(mai_mai_n1048_), .Y(mai_mai_n1351_));
  NO2        m1323(.A(mai_mai_n441_), .B(a), .Y(mai_mai_n1352_));
  NA3        m1324(.A(mai_mai_n1352_), .B(mai_mai_n1351_), .C(mai_mai_n106_), .Y(mai_mai_n1353_));
  NO2        m1325(.A(i), .B(h), .Y(mai_mai_n1354_));
  AOI210     m1326(.A0(mai_mai_n1112_), .A1(h), .B0(mai_mai_n401_), .Y(mai_mai_n1355_));
  NA2        m1327(.A(mai_mai_n128_), .B(mai_mai_n208_), .Y(mai_mai_n1356_));
  NO2        m1328(.A(mai_mai_n1356_), .B(mai_mai_n1355_), .Y(mai_mai_n1357_));
  NO2        m1329(.A(mai_mai_n735_), .B(mai_mai_n175_), .Y(mai_mai_n1358_));
  NOi31      m1330(.An(m), .B(n), .C(b), .Y(mai_mai_n1359_));
  NOi31      m1331(.An(f), .B(d), .C(c), .Y(mai_mai_n1360_));
  NA2        m1332(.A(mai_mai_n1360_), .B(mai_mai_n1359_), .Y(mai_mai_n1361_));
  INV        m1333(.A(mai_mai_n1361_), .Y(mai_mai_n1362_));
  NO3        m1334(.A(mai_mai_n1362_), .B(mai_mai_n1358_), .C(mai_mai_n1357_), .Y(mai_mai_n1363_));
  NA2        m1335(.A(mai_mai_n1059_), .B(mai_mai_n457_), .Y(mai_mai_n1364_));
  NO4        m1336(.A(mai_mai_n1364_), .B(mai_mai_n1033_), .C(mai_mai_n430_), .D(mai_mai_n45_), .Y(mai_mai_n1365_));
  OAI210     m1337(.A0(mai_mai_n169_), .A1(mai_mai_n517_), .B0(mai_mai_n1034_), .Y(mai_mai_n1366_));
  NO3        m1338(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1367_));
  INV        m1339(.A(mai_mai_n1366_), .Y(mai_mai_n1368_));
  NO2        m1340(.A(mai_mai_n1368_), .B(mai_mai_n1365_), .Y(mai_mai_n1369_));
  AN4        m1341(.A(mai_mai_n1369_), .B(mai_mai_n1363_), .C(mai_mai_n1353_), .D(mai_mai_n1350_), .Y(mai_mai_n1370_));
  NA2        m1342(.A(mai_mai_n1315_), .B(mai_mai_n365_), .Y(mai_mai_n1371_));
  NO2        m1343(.A(mai_mai_n1371_), .B(mai_mai_n1015_), .Y(mai_mai_n1372_));
  NO2        m1344(.A(mai_mai_n175_), .B(b), .Y(mai_mai_n1373_));
  AOI220     m1345(.A0(mai_mai_n1143_), .A1(mai_mai_n1373_), .B0(mai_mai_n1067_), .B1(mai_mai_n1364_), .Y(mai_mai_n1374_));
  NAi21      m1346(.An(mai_mai_n1372_), .B(mai_mai_n1374_), .Y(mai_mai_n1375_));
  NO4        m1347(.A(mai_mai_n123_), .B(g), .C(f), .D(e), .Y(mai_mai_n1376_));
  NA3        m1348(.A(mai_mai_n1322_), .B(mai_mai_n277_), .C(h), .Y(mai_mai_n1377_));
  NA2        m1349(.A(mai_mai_n182_), .B(mai_mai_n93_), .Y(mai_mai_n1378_));
  OR2        m1350(.A(e), .B(a), .Y(mai_mai_n1379_));
  NA2        m1351(.A(mai_mai_n30_), .B(h), .Y(mai_mai_n1380_));
  NO2        m1352(.A(mai_mai_n1380_), .B(mai_mai_n1055_), .Y(mai_mai_n1381_));
  NOi41      m1353(.An(h), .B(f), .C(e), .D(a), .Y(mai_mai_n1382_));
  NA2        m1354(.A(mai_mai_n1382_), .B(mai_mai_n106_), .Y(mai_mai_n1383_));
  NA2        m1355(.A(mai_mai_n1318_), .B(mai_mai_n1341_), .Y(mai_mai_n1384_));
  NA2        m1356(.A(mai_mai_n1384_), .B(mai_mai_n1383_), .Y(mai_mai_n1385_));
  OR3        m1357(.A(mai_mai_n531_), .B(mai_mai_n530_), .C(mai_mai_n105_), .Y(mai_mai_n1386_));
  NA2        m1358(.A(mai_mai_n1086_), .B(mai_mai_n394_), .Y(mai_mai_n1387_));
  NO2        m1359(.A(mai_mai_n1387_), .B(mai_mai_n423_), .Y(mai_mai_n1388_));
  AO210      m1360(.A0(mai_mai_n1388_), .A1(mai_mai_n109_), .B0(mai_mai_n1385_), .Y(mai_mai_n1389_));
  NO3        m1361(.A(mai_mai_n1389_), .B(mai_mai_n1381_), .C(mai_mai_n1375_), .Y(mai_mai_n1390_));
  NA4        m1362(.A(mai_mai_n1390_), .B(mai_mai_n1370_), .C(mai_mai_n1344_), .D(mai_mai_n1331_), .Y(mai_mai_n1391_));
  NO2        m1363(.A(mai_mai_n1102_), .B(mai_mai_n103_), .Y(mai_mai_n1392_));
  NA2        m1364(.A(mai_mai_n365_), .B(mai_mai_n56_), .Y(mai_mai_n1393_));
  NA2        m1365(.A(mai_mai_n204_), .B(mai_mai_n166_), .Y(mai_mai_n1394_));
  AOI210     m1366(.A0(mai_mai_n1394_), .A1(mai_mai_n1157_), .B0(mai_mai_n1393_), .Y(mai_mai_n1395_));
  NO2        m1367(.A(mai_mai_n377_), .B(j), .Y(mai_mai_n1396_));
  NA3        m1368(.A(mai_mai_n1367_), .B(mai_mai_n1312_), .C(mai_mai_n1086_), .Y(mai_mai_n1397_));
  NAi41      m1369(.An(mai_mai_n1354_), .B(mai_mai_n1046_), .C(mai_mai_n154_), .D(mai_mai_n137_), .Y(mai_mai_n1398_));
  NA2        m1370(.A(mai_mai_n1398_), .B(mai_mai_n1397_), .Y(mai_mai_n1399_));
  NA3        m1371(.A(g), .B(mai_mai_n1396_), .C(mai_mai_n145_), .Y(mai_mai_n1400_));
  INV        m1372(.A(mai_mai_n1400_), .Y(mai_mai_n1401_));
  NO3        m1373(.A(mai_mai_n730_), .B(mai_mai_n161_), .C(mai_mai_n397_), .Y(mai_mai_n1402_));
  NO3        m1374(.A(mai_mai_n1402_), .B(mai_mai_n1401_), .C(mai_mai_n1399_), .Y(mai_mai_n1403_));
  NO3        m1375(.A(mai_mai_n1055_), .B(mai_mai_n570_), .C(g), .Y(mai_mai_n1404_));
  NOi21      m1376(.An(mai_mai_n1394_), .B(mai_mai_n1404_), .Y(mai_mai_n1405_));
  AOI210     m1377(.A0(mai_mai_n1405_), .A1(mai_mai_n1378_), .B0(mai_mai_n1024_), .Y(mai_mai_n1406_));
  OR2        m1378(.A(n), .B(i), .Y(mai_mai_n1407_));
  OAI210     m1379(.A0(mai_mai_n1407_), .A1(mai_mai_n1045_), .B0(mai_mai_n49_), .Y(mai_mai_n1408_));
  AOI220     m1380(.A0(mai_mai_n1408_), .A1(mai_mai_n1150_), .B0(mai_mai_n798_), .B1(mai_mai_n182_), .Y(mai_mai_n1409_));
  INV        m1381(.A(mai_mai_n1409_), .Y(mai_mai_n1410_));
  OAI220     m1382(.A0(mai_mai_n651_), .A1(g), .B0(mai_mai_n212_), .B1(c), .Y(mai_mai_n1411_));
  INV        m1383(.A(mai_mai_n1411_), .Y(mai_mai_n1412_));
  NO2        m1384(.A(mai_mai_n123_), .B(l), .Y(mai_mai_n1413_));
  NO2        m1385(.A(mai_mai_n212_), .B(k), .Y(mai_mai_n1414_));
  OAI210     m1386(.A0(mai_mai_n1414_), .A1(mai_mai_n1354_), .B0(mai_mai_n1413_), .Y(mai_mai_n1415_));
  OAI220     m1387(.A0(mai_mai_n1415_), .A1(mai_mai_n31_), .B0(mai_mai_n1412_), .B1(mai_mai_n163_), .Y(mai_mai_n1416_));
  NO3        m1388(.A(mai_mai_n1386_), .B(mai_mai_n457_), .C(mai_mai_n339_), .Y(mai_mai_n1417_));
  NO4        m1389(.A(mai_mai_n1417_), .B(mai_mai_n1416_), .C(mai_mai_n1410_), .D(mai_mai_n1406_), .Y(mai_mai_n1418_));
  NO3        m1390(.A(mai_mai_n1070_), .B(mai_mai_n1312_), .C(mai_mai_n49_), .Y(mai_mai_n1419_));
  NO2        m1391(.A(mai_mai_n1055_), .B(h), .Y(mai_mai_n1420_));
  NA3        m1392(.A(mai_mai_n1420_), .B(d), .C(mai_mai_n1016_), .Y(mai_mai_n1421_));
  NO2        m1393(.A(mai_mai_n1421_), .B(c), .Y(mai_mai_n1422_));
  NA3        m1394(.A(mai_mai_n1392_), .B(mai_mai_n457_), .C(f), .Y(mai_mai_n1423_));
  NA2        m1395(.A(mai_mai_n166_), .B(mai_mai_n105_), .Y(mai_mai_n1424_));
  NO2        m1396(.A(mai_mai_n1306_), .B(mai_mai_n42_), .Y(mai_mai_n1425_));
  AOI210     m1397(.A0(mai_mai_n106_), .A1(mai_mai_n40_), .B0(mai_mai_n1425_), .Y(mai_mai_n1426_));
  NO2        m1398(.A(mai_mai_n1426_), .B(mai_mai_n1423_), .Y(mai_mai_n1427_));
  NOi21      m1399(.An(d), .B(f), .Y(mai_mai_n1428_));
  NO2        m1400(.A(mai_mai_n1312_), .B(f), .Y(mai_mai_n1429_));
  NA2        m1401(.A(mai_mai_n1352_), .B(mai_mai_n1425_), .Y(mai_mai_n1430_));
  INV        m1402(.A(mai_mai_n1430_), .Y(mai_mai_n1431_));
  NO3        m1403(.A(mai_mai_n1431_), .B(mai_mai_n1427_), .C(mai_mai_n1422_), .Y(mai_mai_n1432_));
  NA4        m1404(.A(mai_mai_n1432_), .B(mai_mai_n1418_), .C(mai_mai_n1403_), .D(mai_mai_n1510_), .Y(mai_mai_n1433_));
  NO3        m1405(.A(mai_mai_n1059_), .B(mai_mai_n1045_), .C(mai_mai_n40_), .Y(mai_mai_n1434_));
  NO2        m1406(.A(mai_mai_n457_), .B(mai_mai_n286_), .Y(mai_mai_n1435_));
  OAI210     m1407(.A0(mai_mai_n1435_), .A1(mai_mai_n1434_), .B0(mai_mai_n1327_), .Y(mai_mai_n1436_));
  OAI210     m1408(.A0(mai_mai_n1376_), .A1(mai_mai_n1315_), .B0(mai_mai_n858_), .Y(mai_mai_n1437_));
  NO2        m1409(.A(mai_mai_n1012_), .B(mai_mai_n123_), .Y(mai_mai_n1438_));
  NA2        m1410(.A(mai_mai_n1438_), .B(mai_mai_n612_), .Y(mai_mai_n1439_));
  NA3        m1411(.A(mai_mai_n1439_), .B(mai_mai_n1437_), .C(mai_mai_n1436_), .Y(mai_mai_n1440_));
  NA2        m1412(.A(mai_mai_n1347_), .B(mai_mai_n1428_), .Y(mai_mai_n1441_));
  NO2        m1413(.A(mai_mai_n1441_), .B(m), .Y(mai_mai_n1442_));
  NO2        m1414(.A(mai_mai_n138_), .B(mai_mai_n168_), .Y(mai_mai_n1443_));
  OAI210     m1415(.A0(mai_mai_n1443_), .A1(mai_mai_n103_), .B0(mai_mai_n1359_), .Y(mai_mai_n1444_));
  INV        m1416(.A(mai_mai_n1444_), .Y(mai_mai_n1445_));
  NO3        m1417(.A(mai_mai_n1445_), .B(mai_mai_n1442_), .C(mai_mai_n1440_), .Y(mai_mai_n1446_));
  NO2        m1418(.A(mai_mai_n1311_), .B(e), .Y(mai_mai_n1447_));
  NA2        m1419(.A(mai_mai_n1447_), .B(mai_mai_n392_), .Y(mai_mai_n1448_));
  NA2        m1420(.A(mai_mai_n1097_), .B(mai_mai_n619_), .Y(mai_mai_n1449_));
  OR3        m1421(.A(mai_mai_n1414_), .B(mai_mai_n1183_), .C(mai_mai_n123_), .Y(mai_mai_n1450_));
  OAI220     m1422(.A0(mai_mai_n1450_), .A1(mai_mai_n1448_), .B0(mai_mai_n1449_), .B1(mai_mai_n432_), .Y(mai_mai_n1451_));
  INV        m1423(.A(mai_mai_n1451_), .Y(mai_mai_n1452_));
  NO2        m1424(.A(mai_mai_n168_), .B(c), .Y(mai_mai_n1453_));
  OAI210     m1425(.A0(mai_mai_n1453_), .A1(mai_mai_n1447_), .B0(mai_mai_n166_), .Y(mai_mai_n1454_));
  AOI220     m1426(.A0(mai_mai_n1454_), .A1(mai_mai_n1047_), .B0(mai_mai_n524_), .B1(mai_mai_n353_), .Y(mai_mai_n1455_));
  NA2        m1427(.A(mai_mai_n530_), .B(g), .Y(mai_mai_n1456_));
  AOI210     m1428(.A0(mai_mai_n1456_), .A1(mai_mai_n1343_), .B0(mai_mai_n1419_), .Y(mai_mai_n1457_));
  NO2        m1429(.A(mai_mai_n1379_), .B(f), .Y(mai_mai_n1458_));
  NO2        m1430(.A(mai_mai_n1457_), .B(mai_mai_n202_), .Y(mai_mai_n1459_));
  AOI210     m1431(.A0(mai_mai_n877_), .A1(mai_mai_n403_), .B0(mai_mai_n97_), .Y(mai_mai_n1460_));
  OR2        m1432(.A(mai_mai_n1460_), .B(mai_mai_n530_), .Y(mai_mai_n1461_));
  NA2        m1433(.A(mai_mai_n1458_), .B(mai_mai_n1324_), .Y(mai_mai_n1462_));
  OAI220     m1434(.A0(mai_mai_n1462_), .A1(mai_mai_n49_), .B0(mai_mai_n1461_), .B1(mai_mai_n161_), .Y(mai_mai_n1463_));
  NA4        m1435(.A(mai_mai_n1068_), .B(mai_mai_n1065_), .C(mai_mai_n208_), .D(mai_mai_n68_), .Y(mai_mai_n1464_));
  NA2        m1436(.A(mai_mai_n1316_), .B(mai_mai_n169_), .Y(mai_mai_n1465_));
  NO2        m1437(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1466_));
  OAI210     m1438(.A0(mai_mai_n1379_), .A1(mai_mai_n836_), .B0(mai_mai_n476_), .Y(mai_mai_n1467_));
  OAI210     m1439(.A0(mai_mai_n1467_), .A1(mai_mai_n1071_), .B0(mai_mai_n1466_), .Y(mai_mai_n1468_));
  NO2        m1440(.A(mai_mai_n238_), .B(g), .Y(mai_mai_n1469_));
  NO2        m1441(.A(m), .B(i), .Y(mai_mai_n1470_));
  BUFFER     m1442(.A(mai_mai_n1470_), .Y(mai_mai_n1471_));
  AOI220     m1443(.A0(mai_mai_n1471_), .A1(mai_mai_n1345_), .B0(mai_mai_n1046_), .B1(mai_mai_n1469_), .Y(mai_mai_n1472_));
  NA4        m1444(.A(mai_mai_n1472_), .B(mai_mai_n1468_), .C(mai_mai_n1465_), .D(mai_mai_n1464_), .Y(mai_mai_n1473_));
  NO4        m1445(.A(mai_mai_n1473_), .B(mai_mai_n1463_), .C(mai_mai_n1459_), .D(mai_mai_n1455_), .Y(mai_mai_n1474_));
  NA3        m1446(.A(mai_mai_n1474_), .B(mai_mai_n1452_), .C(mai_mai_n1446_), .Y(mai_mai_n1475_));
  NA3        m1447(.A(mai_mai_n937_), .B(mai_mai_n128_), .C(mai_mai_n46_), .Y(mai_mai_n1476_));
  AOI210     m1448(.A0(mai_mai_n135_), .A1(c), .B0(mai_mai_n1476_), .Y(mai_mai_n1477_));
  INV        m1449(.A(mai_mai_n172_), .Y(mai_mai_n1478_));
  NA2        m1450(.A(mai_mai_n1478_), .B(mai_mai_n1420_), .Y(mai_mai_n1479_));
  OR2        m1451(.A(mai_mai_n124_), .B(mai_mai_n1371_), .Y(mai_mai_n1480_));
  NA2        m1452(.A(mai_mai_n1480_), .B(mai_mai_n1479_), .Y(mai_mai_n1481_));
  NO2        m1453(.A(mai_mai_n1481_), .B(mai_mai_n1477_), .Y(mai_mai_n1482_));
  AOI210     m1454(.A0(mai_mai_n143_), .A1(mai_mai_n56_), .B0(mai_mai_n1447_), .Y(mai_mai_n1483_));
  NO2        m1455(.A(mai_mai_n1483_), .B(mai_mai_n1424_), .Y(mai_mai_n1484_));
  NOi21      m1456(.An(mai_mai_n1316_), .B(e), .Y(mai_mai_n1485_));
  NO2        m1457(.A(mai_mai_n1485_), .B(mai_mai_n1484_), .Y(mai_mai_n1486_));
  AN2        m1458(.A(mai_mai_n1068_), .B(mai_mai_n1053_), .Y(mai_mai_n1487_));
  NA2        m1459(.A(mai_mai_n1030_), .B(mai_mai_n146_), .Y(mai_mai_n1488_));
  NOi31      m1460(.An(mai_mai_n30_), .B(mai_mai_n1488_), .C(n), .Y(mai_mai_n1489_));
  AOI210     m1461(.A0(mai_mai_n1487_), .A1(mai_mai_n1143_), .B0(mai_mai_n1489_), .Y(mai_mai_n1490_));
  NO2        m1462(.A(mai_mai_n1423_), .B(mai_mai_n69_), .Y(mai_mai_n1491_));
  NA2        m1463(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1492_));
  NO2        m1464(.A(mai_mai_n1322_), .B(mai_mai_n111_), .Y(mai_mai_n1493_));
  OAI220     m1465(.A0(mai_mai_n1493_), .A1(mai_mai_n1371_), .B0(mai_mai_n1387_), .B1(mai_mai_n1492_), .Y(mai_mai_n1494_));
  NO2        m1466(.A(mai_mai_n1494_), .B(mai_mai_n1491_), .Y(mai_mai_n1495_));
  NA4        m1467(.A(mai_mai_n1495_), .B(mai_mai_n1490_), .C(mai_mai_n1486_), .D(mai_mai_n1482_), .Y(mai_mai_n1496_));
  OR4        m1468(.A(mai_mai_n1496_), .B(mai_mai_n1475_), .C(mai_mai_n1433_), .D(mai_mai_n1391_), .Y(mai04));
  NOi31      m1469(.An(mai_mai_n1376_), .B(mai_mai_n1377_), .C(mai_mai_n1018_), .Y(mai_mai_n1498_));
  NA2        m1470(.A(mai_mai_n1429_), .B(mai_mai_n798_), .Y(mai_mai_n1499_));
  NO3        m1471(.A(mai_mai_n1499_), .B(mai_mai_n1007_), .C(mai_mai_n477_), .Y(mai_mai_n1500_));
  OR3        m1472(.A(mai_mai_n1500_), .B(mai_mai_n1498_), .C(mai_mai_n1036_), .Y(mai_mai_n1501_));
  NO3        m1473(.A(mai_mai_n1324_), .B(mai_mai_n87_), .C(k), .Y(mai_mai_n1502_));
  AOI210     m1474(.A0(mai_mai_n1502_), .A1(mai_mai_n1029_), .B0(mai_mai_n1159_), .Y(mai_mai_n1503_));
  NA2        m1475(.A(mai_mai_n1503_), .B(mai_mai_n1187_), .Y(mai_mai_n1504_));
  NO4        m1476(.A(mai_mai_n1504_), .B(mai_mai_n1501_), .C(mai_mai_n1044_), .D(mai_mai_n1023_), .Y(mai_mai_n1505_));
  NA4        m1477(.A(mai_mai_n1505_), .B(mai_mai_n1099_), .C(mai_mai_n1084_), .D(mai_mai_n1074_), .Y(mai05));
  INV        m1478(.A(m), .Y(mai_mai_n1509_));
  INV        m1479(.A(mai_mai_n1395_), .Y(mai_mai_n1510_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi31      u0013(.An(n), .B(m), .C(l), .Y(men_men_n42_));
  INV        u0014(.A(i), .Y(men_men_n43_));
  AN2        u0015(.A(h), .B(g), .Y(men_men_n44_));
  NA2        u0016(.A(men_men_n44_), .B(men_men_n43_), .Y(men_men_n45_));
  NO2        u0017(.A(men_men_n45_), .B(men_men_n42_), .Y(men_men_n46_));
  NAi21      u0018(.An(n), .B(m), .Y(men_men_n47_));
  NOi32      u0019(.An(k), .Bn(h), .C(l), .Y(men_men_n48_));
  NOi32      u0020(.An(k), .Bn(h), .C(g), .Y(men_men_n49_));
  INV        u0021(.A(men_men_n39_), .Y(men_men_n50_));
  NO2        u0022(.A(men_men_n50_), .B(men_men_n32_), .Y(men_men_n51_));
  INV        u0023(.A(c), .Y(men_men_n52_));
  NA2        u0024(.A(e), .B(b), .Y(men_men_n53_));
  NO2        u0025(.A(men_men_n53_), .B(men_men_n52_), .Y(men_men_n54_));
  INV        u0026(.A(d), .Y(men_men_n55_));
  NA2        u0027(.A(g), .B(men_men_n55_), .Y(men_men_n56_));
  NAi21      u0028(.An(i), .B(h), .Y(men_men_n57_));
  NAi31      u0029(.An(i), .B(l), .C(j), .Y(men_men_n58_));
  OAI220     u0030(.A0(men_men_n58_), .A1(men_men_n47_), .B0(men_men_n57_), .B1(men_men_n42_), .Y(men_men_n59_));
  NAi31      u0031(.An(men_men_n56_), .B(men_men_n59_), .C(men_men_n54_), .Y(men_men_n60_));
  NAi41      u0032(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n61_));
  NA2        u0033(.A(g), .B(f), .Y(men_men_n62_));
  NO2        u0034(.A(men_men_n62_), .B(men_men_n61_), .Y(men_men_n63_));
  NAi21      u0035(.An(i), .B(j), .Y(men_men_n64_));
  NAi32      u0036(.An(n), .Bn(k), .C(m), .Y(men_men_n65_));
  NO2        u0037(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NAi31      u0038(.An(l), .B(m), .C(k), .Y(men_men_n67_));
  NAi21      u0039(.An(e), .B(h), .Y(men_men_n68_));
  NAi41      u0040(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n69_));
  NA2        u0041(.A(men_men_n66_), .B(men_men_n63_), .Y(men_men_n70_));
  INV        u0042(.A(m), .Y(men_men_n71_));
  NOi21      u0043(.An(k), .B(l), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n72_), .B(men_men_n71_), .Y(men_men_n73_));
  AN4        u0045(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n74_));
  NOi31      u0046(.An(h), .B(g), .C(f), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  NAi32      u0048(.An(m), .Bn(k), .C(j), .Y(men_men_n77_));
  NOi32      u0049(.An(h), .Bn(g), .C(f), .Y(men_men_n78_));
  NA2        u0050(.A(men_men_n78_), .B(men_men_n74_), .Y(men_men_n79_));
  OA220      u0051(.A0(men_men_n79_), .A1(men_men_n77_), .B0(men_men_n76_), .B1(men_men_n73_), .Y(men_men_n80_));
  NA3        u0052(.A(men_men_n80_), .B(men_men_n70_), .C(men_men_n60_), .Y(men_men_n81_));
  INV        u0053(.A(n), .Y(men_men_n82_));
  NOi32      u0054(.An(e), .Bn(b), .C(d), .Y(men_men_n83_));
  NA2        u0055(.A(men_men_n83_), .B(men_men_n82_), .Y(men_men_n84_));
  INV        u0056(.A(j), .Y(men_men_n85_));
  AN3        u0057(.A(m), .B(k), .C(i), .Y(men_men_n86_));
  NA3        u0058(.A(men_men_n86_), .B(men_men_n85_), .C(g), .Y(men_men_n87_));
  NO2        u0059(.A(men_men_n87_), .B(f), .Y(men_men_n88_));
  NAi32      u0060(.An(g), .Bn(f), .C(h), .Y(men_men_n89_));
  NAi31      u0061(.An(j), .B(m), .C(l), .Y(men_men_n90_));
  NO2        u0062(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n91_));
  NA2        u0063(.A(m), .B(l), .Y(men_men_n92_));
  NAi31      u0064(.An(k), .B(j), .C(g), .Y(men_men_n93_));
  NO3        u0065(.A(men_men_n93_), .B(men_men_n92_), .C(f), .Y(men_men_n94_));
  AN2        u0066(.A(j), .B(g), .Y(men_men_n95_));
  NOi32      u0067(.An(m), .Bn(l), .C(i), .Y(men_men_n96_));
  NOi21      u0068(.An(g), .B(i), .Y(men_men_n97_));
  NOi32      u0069(.An(m), .Bn(j), .C(k), .Y(men_men_n98_));
  AOI220     u0070(.A0(men_men_n98_), .A1(men_men_n97_), .B0(men_men_n96_), .B1(men_men_n95_), .Y(men_men_n99_));
  NO2        u0071(.A(men_men_n99_), .B(f), .Y(men_men_n100_));
  NO4        u0072(.A(men_men_n100_), .B(men_men_n94_), .C(men_men_n91_), .D(men_men_n88_), .Y(men_men_n101_));
  NAi41      u0073(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n102_));
  AN2        u0074(.A(e), .B(b), .Y(men_men_n103_));
  NOi31      u0075(.An(c), .B(h), .C(f), .Y(men_men_n104_));
  NA2        u0076(.A(men_men_n104_), .B(men_men_n103_), .Y(men_men_n105_));
  NO2        u0077(.A(men_men_n105_), .B(men_men_n102_), .Y(men_men_n106_));
  NOi21      u0078(.An(g), .B(f), .Y(men_men_n107_));
  NOi21      u0079(.An(i), .B(h), .Y(men_men_n108_));
  NA3        u0080(.A(men_men_n108_), .B(men_men_n107_), .C(men_men_n36_), .Y(men_men_n109_));
  INV        u0081(.A(a), .Y(men_men_n110_));
  NA2        u0082(.A(men_men_n103_), .B(men_men_n110_), .Y(men_men_n111_));
  INV        u0083(.A(l), .Y(men_men_n112_));
  NOi21      u0084(.An(m), .B(n), .Y(men_men_n113_));
  AN2        u0085(.A(k), .B(h), .Y(men_men_n114_));
  NO2        u0086(.A(men_men_n109_), .B(men_men_n84_), .Y(men_men_n115_));
  INV        u0087(.A(b), .Y(men_men_n116_));
  NA2        u0088(.A(l), .B(j), .Y(men_men_n117_));
  AN2        u0089(.A(k), .B(i), .Y(men_men_n118_));
  NA2        u0090(.A(men_men_n118_), .B(men_men_n117_), .Y(men_men_n119_));
  NA2        u0091(.A(g), .B(e), .Y(men_men_n120_));
  NOi32      u0092(.An(c), .Bn(a), .C(d), .Y(men_men_n121_));
  NA2        u0093(.A(men_men_n121_), .B(men_men_n113_), .Y(men_men_n122_));
  NO4        u0094(.A(men_men_n122_), .B(men_men_n120_), .C(men_men_n119_), .D(men_men_n116_), .Y(men_men_n123_));
  NO3        u0095(.A(men_men_n123_), .B(men_men_n115_), .C(men_men_n106_), .Y(men_men_n124_));
  OAI210     u0096(.A0(men_men_n101_), .A1(men_men_n84_), .B0(men_men_n124_), .Y(men_men_n125_));
  NOi31      u0097(.An(k), .B(m), .C(j), .Y(men_men_n126_));
  NA3        u0098(.A(men_men_n126_), .B(men_men_n75_), .C(men_men_n74_), .Y(men_men_n127_));
  NOi31      u0099(.An(k), .B(m), .C(i), .Y(men_men_n128_));
  NA3        u0100(.A(men_men_n128_), .B(men_men_n78_), .C(men_men_n74_), .Y(men_men_n129_));
  NA2        u0101(.A(men_men_n129_), .B(men_men_n127_), .Y(men_men_n130_));
  NOi32      u0102(.An(f), .Bn(b), .C(e), .Y(men_men_n131_));
  NAi21      u0103(.An(g), .B(h), .Y(men_men_n132_));
  NAi21      u0104(.An(m), .B(n), .Y(men_men_n133_));
  NAi21      u0105(.An(j), .B(k), .Y(men_men_n134_));
  NO3        u0106(.A(men_men_n134_), .B(men_men_n133_), .C(men_men_n132_), .Y(men_men_n135_));
  NAi41      u0107(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n136_));
  NAi31      u0108(.An(j), .B(k), .C(h), .Y(men_men_n137_));
  NO3        u0109(.A(men_men_n137_), .B(men_men_n136_), .C(men_men_n133_), .Y(men_men_n138_));
  AOI210     u0110(.A0(men_men_n135_), .A1(men_men_n131_), .B0(men_men_n138_), .Y(men_men_n139_));
  NO2        u0111(.A(k), .B(j), .Y(men_men_n140_));
  NO2        u0112(.A(men_men_n140_), .B(men_men_n133_), .Y(men_men_n141_));
  AN2        u0113(.A(k), .B(j), .Y(men_men_n142_));
  NAi21      u0114(.An(c), .B(b), .Y(men_men_n143_));
  NA2        u0115(.A(f), .B(d), .Y(men_men_n144_));
  NO3        u0116(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n132_), .Y(men_men_n145_));
  NA2        u0117(.A(h), .B(c), .Y(men_men_n146_));
  NAi31      u0118(.An(f), .B(e), .C(b), .Y(men_men_n147_));
  NA2        u0119(.A(men_men_n145_), .B(men_men_n141_), .Y(men_men_n148_));
  NA2        u0120(.A(d), .B(b), .Y(men_men_n149_));
  NAi21      u0121(.An(e), .B(f), .Y(men_men_n150_));
  NO2        u0122(.A(men_men_n150_), .B(men_men_n149_), .Y(men_men_n151_));
  NA2        u0123(.A(b), .B(a), .Y(men_men_n152_));
  NAi21      u0124(.An(e), .B(g), .Y(men_men_n153_));
  NAi21      u0125(.An(c), .B(d), .Y(men_men_n154_));
  NAi31      u0126(.An(l), .B(k), .C(h), .Y(men_men_n155_));
  NO2        u0127(.A(men_men_n133_), .B(men_men_n155_), .Y(men_men_n156_));
  NA2        u0128(.A(men_men_n156_), .B(men_men_n151_), .Y(men_men_n157_));
  NAi41      u0129(.An(men_men_n130_), .B(men_men_n157_), .C(men_men_n148_), .D(men_men_n139_), .Y(men_men_n158_));
  NAi31      u0130(.An(e), .B(f), .C(b), .Y(men_men_n159_));
  NOi21      u0131(.An(g), .B(d), .Y(men_men_n160_));
  NO2        u0132(.A(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  NOi21      u0133(.An(h), .B(i), .Y(men_men_n162_));
  NOi21      u0134(.An(k), .B(m), .Y(men_men_n163_));
  NA3        u0135(.A(men_men_n163_), .B(men_men_n162_), .C(n), .Y(men_men_n164_));
  NOi21      u0136(.An(men_men_n161_), .B(men_men_n164_), .Y(men_men_n165_));
  NOi21      u0137(.An(h), .B(g), .Y(men_men_n166_));
  NO2        u0138(.A(men_men_n144_), .B(men_men_n143_), .Y(men_men_n167_));
  NAi31      u0139(.An(l), .B(j), .C(h), .Y(men_men_n168_));
  NO2        u0140(.A(men_men_n168_), .B(men_men_n47_), .Y(men_men_n169_));
  NA2        u0141(.A(men_men_n169_), .B(men_men_n63_), .Y(men_men_n170_));
  NOi32      u0142(.An(n), .Bn(k), .C(m), .Y(men_men_n171_));
  NA2        u0143(.A(l), .B(i), .Y(men_men_n172_));
  INV        u0144(.A(men_men_n170_), .Y(men_men_n173_));
  NAi31      u0145(.An(d), .B(f), .C(c), .Y(men_men_n174_));
  NAi31      u0146(.An(e), .B(f), .C(c), .Y(men_men_n175_));
  NA2        u0147(.A(men_men_n175_), .B(men_men_n174_), .Y(men_men_n176_));
  NA2        u0148(.A(j), .B(h), .Y(men_men_n177_));
  OR3        u0149(.A(n), .B(m), .C(k), .Y(men_men_n178_));
  NO2        u0150(.A(men_men_n178_), .B(men_men_n177_), .Y(men_men_n179_));
  NAi32      u0151(.An(m), .Bn(k), .C(n), .Y(men_men_n180_));
  NO2        u0152(.A(men_men_n180_), .B(men_men_n177_), .Y(men_men_n181_));
  AOI220     u0153(.A0(men_men_n181_), .A1(men_men_n161_), .B0(men_men_n179_), .B1(men_men_n176_), .Y(men_men_n182_));
  NO2        u0154(.A(n), .B(m), .Y(men_men_n183_));
  NA2        u0155(.A(men_men_n183_), .B(men_men_n48_), .Y(men_men_n184_));
  NAi21      u0156(.An(f), .B(e), .Y(men_men_n185_));
  NA2        u0157(.A(d), .B(c), .Y(men_men_n186_));
  NAi21      u0158(.An(d), .B(c), .Y(men_men_n187_));
  NAi31      u0159(.An(m), .B(n), .C(b), .Y(men_men_n188_));
  NA2        u0160(.A(k), .B(i), .Y(men_men_n189_));
  NAi21      u0161(.An(h), .B(f), .Y(men_men_n190_));
  NO2        u0162(.A(men_men_n188_), .B(men_men_n154_), .Y(men_men_n191_));
  NOi32      u0163(.An(f), .Bn(c), .C(d), .Y(men_men_n192_));
  NOi32      u0164(.An(f), .Bn(c), .C(e), .Y(men_men_n193_));
  NO2        u0165(.A(men_men_n193_), .B(men_men_n192_), .Y(men_men_n194_));
  NO3        u0166(.A(n), .B(m), .C(j), .Y(men_men_n195_));
  NA2        u0167(.A(men_men_n195_), .B(men_men_n114_), .Y(men_men_n196_));
  AO210      u0168(.A0(men_men_n196_), .A1(men_men_n184_), .B0(men_men_n194_), .Y(men_men_n197_));
  NA2        u0169(.A(men_men_n197_), .B(men_men_n182_), .Y(men_men_n198_));
  OR4        u0170(.A(men_men_n198_), .B(men_men_n173_), .C(men_men_n165_), .D(men_men_n158_), .Y(men_men_n199_));
  NO4        u0171(.A(men_men_n199_), .B(men_men_n125_), .C(men_men_n81_), .D(men_men_n51_), .Y(men_men_n200_));
  NA3        u0172(.A(m), .B(men_men_n112_), .C(j), .Y(men_men_n201_));
  NAi31      u0173(.An(n), .B(h), .C(g), .Y(men_men_n202_));
  NO2        u0174(.A(men_men_n202_), .B(men_men_n201_), .Y(men_men_n203_));
  NOi32      u0175(.An(m), .Bn(k), .C(l), .Y(men_men_n204_));
  NA3        u0176(.A(men_men_n204_), .B(men_men_n85_), .C(g), .Y(men_men_n205_));
  AN2        u0177(.A(i), .B(g), .Y(men_men_n206_));
  NA3        u0178(.A(men_men_n72_), .B(men_men_n206_), .C(men_men_n113_), .Y(men_men_n207_));
  INV        u0179(.A(men_men_n207_), .Y(men_men_n208_));
  NO2        u0180(.A(men_men_n208_), .B(men_men_n203_), .Y(men_men_n209_));
  NAi41      u0181(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n210_));
  INV        u0182(.A(men_men_n210_), .Y(men_men_n211_));
  INV        u0183(.A(f), .Y(men_men_n212_));
  INV        u0184(.A(g), .Y(men_men_n213_));
  NOi31      u0185(.An(i), .B(j), .C(h), .Y(men_men_n214_));
  NOi21      u0186(.An(l), .B(m), .Y(men_men_n215_));
  NA2        u0187(.A(men_men_n215_), .B(men_men_n214_), .Y(men_men_n216_));
  NO3        u0188(.A(men_men_n216_), .B(men_men_n213_), .C(men_men_n212_), .Y(men_men_n217_));
  NA2        u0189(.A(men_men_n217_), .B(men_men_n211_), .Y(men_men_n218_));
  OAI210     u0190(.A0(men_men_n209_), .A1(men_men_n32_), .B0(men_men_n218_), .Y(men_men_n219_));
  NOi21      u0191(.An(n), .B(m), .Y(men_men_n220_));
  NOi32      u0192(.An(l), .Bn(i), .C(j), .Y(men_men_n221_));
  NA2        u0193(.A(men_men_n221_), .B(men_men_n220_), .Y(men_men_n222_));
  OA220      u0194(.A0(men_men_n222_), .A1(men_men_n105_), .B0(men_men_n77_), .B1(men_men_n76_), .Y(men_men_n223_));
  NAi21      u0195(.An(j), .B(h), .Y(men_men_n224_));
  XN2        u0196(.A(i), .B(h), .Y(men_men_n225_));
  NA2        u0197(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  NOi31      u0198(.An(k), .B(n), .C(m), .Y(men_men_n227_));
  NOi31      u0199(.An(men_men_n227_), .B(men_men_n186_), .C(men_men_n185_), .Y(men_men_n228_));
  NA2        u0200(.A(men_men_n228_), .B(men_men_n226_), .Y(men_men_n229_));
  NAi31      u0201(.An(f), .B(e), .C(c), .Y(men_men_n230_));
  NO4        u0202(.A(men_men_n230_), .B(men_men_n178_), .C(men_men_n177_), .D(men_men_n55_), .Y(men_men_n231_));
  NA4        u0203(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n232_));
  NAi32      u0204(.An(m), .Bn(i), .C(k), .Y(men_men_n233_));
  NO3        u0205(.A(men_men_n233_), .B(men_men_n89_), .C(men_men_n232_), .Y(men_men_n234_));
  INV        u0206(.A(k), .Y(men_men_n235_));
  NO2        u0207(.A(men_men_n234_), .B(men_men_n231_), .Y(men_men_n236_));
  NAi21      u0208(.An(n), .B(a), .Y(men_men_n237_));
  NO2        u0209(.A(men_men_n237_), .B(men_men_n149_), .Y(men_men_n238_));
  NAi41      u0210(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n239_));
  NO2        u0211(.A(men_men_n239_), .B(e), .Y(men_men_n240_));
  NO3        u0212(.A(men_men_n150_), .B(men_men_n93_), .C(men_men_n92_), .Y(men_men_n241_));
  OAI210     u0213(.A0(men_men_n241_), .A1(men_men_n240_), .B0(men_men_n238_), .Y(men_men_n242_));
  AN4        u0214(.A(men_men_n242_), .B(men_men_n236_), .C(men_men_n229_), .D(men_men_n223_), .Y(men_men_n243_));
  OR2        u0215(.A(h), .B(g), .Y(men_men_n244_));
  NAi41      u0216(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n245_));
  NO2        u0217(.A(men_men_n245_), .B(men_men_n212_), .Y(men_men_n246_));
  NA2        u0218(.A(men_men_n163_), .B(men_men_n108_), .Y(men_men_n247_));
  NAi21      u0219(.An(men_men_n247_), .B(men_men_n246_), .Y(men_men_n248_));
  NO2        u0220(.A(n), .B(a), .Y(men_men_n249_));
  NAi31      u0221(.An(men_men_n239_), .B(men_men_n249_), .C(men_men_n103_), .Y(men_men_n250_));
  AN2        u0222(.A(men_men_n250_), .B(men_men_n248_), .Y(men_men_n251_));
  NAi21      u0223(.An(h), .B(i), .Y(men_men_n252_));
  NA2        u0224(.A(men_men_n183_), .B(k), .Y(men_men_n253_));
  NO2        u0225(.A(men_men_n253_), .B(men_men_n252_), .Y(men_men_n254_));
  NA2        u0226(.A(men_men_n254_), .B(men_men_n192_), .Y(men_men_n255_));
  NA2        u0227(.A(men_men_n255_), .B(men_men_n251_), .Y(men_men_n256_));
  NOi21      u0228(.An(g), .B(e), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n69_), .B(men_men_n71_), .Y(men_men_n258_));
  NOi32      u0230(.An(l), .Bn(j), .C(i), .Y(men_men_n259_));
  AOI210     u0231(.A0(men_men_n72_), .A1(men_men_n85_), .B0(men_men_n259_), .Y(men_men_n260_));
  NO2        u0232(.A(men_men_n252_), .B(men_men_n42_), .Y(men_men_n261_));
  NAi21      u0233(.An(f), .B(g), .Y(men_men_n262_));
  NO2        u0234(.A(men_men_n262_), .B(men_men_n61_), .Y(men_men_n263_));
  NO2        u0235(.A(men_men_n65_), .B(men_men_n117_), .Y(men_men_n264_));
  AOI220     u0236(.A0(men_men_n264_), .A1(men_men_n263_), .B0(men_men_n261_), .B1(men_men_n63_), .Y(men_men_n265_));
  INV        u0237(.A(men_men_n265_), .Y(men_men_n266_));
  NO3        u0238(.A(men_men_n134_), .B(men_men_n47_), .C(men_men_n43_), .Y(men_men_n267_));
  NOi41      u0239(.An(men_men_n243_), .B(men_men_n266_), .C(men_men_n256_), .D(men_men_n219_), .Y(men_men_n268_));
  NO3        u0240(.A(men_men_n203_), .B(men_men_n46_), .C(men_men_n39_), .Y(men_men_n269_));
  NO2        u0241(.A(men_men_n269_), .B(men_men_n111_), .Y(men_men_n270_));
  NA3        u0242(.A(men_men_n55_), .B(c), .C(b), .Y(men_men_n271_));
  NAi21      u0243(.An(h), .B(g), .Y(men_men_n272_));
  OR4        u0244(.A(men_men_n272_), .B(men_men_n271_), .C(men_men_n222_), .D(e), .Y(men_men_n273_));
  NAi31      u0245(.An(g), .B(k), .C(h), .Y(men_men_n274_));
  NAi31      u0246(.An(e), .B(d), .C(a), .Y(men_men_n275_));
  INV        u0247(.A(men_men_n273_), .Y(men_men_n276_));
  NA3        u0248(.A(men_men_n163_), .B(men_men_n162_), .C(men_men_n82_), .Y(men_men_n277_));
  NO2        u0249(.A(men_men_n277_), .B(men_men_n194_), .Y(men_men_n278_));
  INV        u0250(.A(men_men_n278_), .Y(men_men_n279_));
  NA3        u0251(.A(e), .B(c), .C(b), .Y(men_men_n280_));
  NAi32      u0252(.An(k), .Bn(i), .C(j), .Y(men_men_n281_));
  NAi21      u0253(.An(l), .B(k), .Y(men_men_n282_));
  NO2        u0254(.A(men_men_n282_), .B(men_men_n47_), .Y(men_men_n283_));
  NOi21      u0255(.An(l), .B(j), .Y(men_men_n284_));
  NA2        u0256(.A(men_men_n166_), .B(men_men_n284_), .Y(men_men_n285_));
  NA3        u0257(.A(men_men_n118_), .B(men_men_n117_), .C(g), .Y(men_men_n286_));
  OR3        u0258(.A(men_men_n69_), .B(men_men_n71_), .C(e), .Y(men_men_n287_));
  AOI210     u0259(.A0(men_men_n286_), .A1(men_men_n285_), .B0(men_men_n287_), .Y(men_men_n288_));
  INV        u0260(.A(men_men_n288_), .Y(men_men_n289_));
  NAi32      u0261(.An(j), .Bn(h), .C(i), .Y(men_men_n290_));
  NAi21      u0262(.An(m), .B(l), .Y(men_men_n291_));
  NO3        u0263(.A(men_men_n291_), .B(men_men_n290_), .C(men_men_n82_), .Y(men_men_n292_));
  NA2        u0264(.A(h), .B(g), .Y(men_men_n293_));
  NA2        u0265(.A(men_men_n171_), .B(men_men_n43_), .Y(men_men_n294_));
  NO2        u0266(.A(men_men_n294_), .B(men_men_n293_), .Y(men_men_n295_));
  NA2        u0267(.A(men_men_n295_), .B(men_men_n167_), .Y(men_men_n296_));
  NA3        u0268(.A(men_men_n296_), .B(men_men_n289_), .C(men_men_n279_), .Y(men_men_n297_));
  NO2        u0269(.A(men_men_n147_), .B(d), .Y(men_men_n298_));
  NO2        u0270(.A(men_men_n105_), .B(men_men_n102_), .Y(men_men_n299_));
  NAi32      u0271(.An(n), .Bn(m), .C(l), .Y(men_men_n300_));
  NO2        u0272(.A(men_men_n300_), .B(men_men_n290_), .Y(men_men_n301_));
  NO2        u0273(.A(men_men_n122_), .B(men_men_n116_), .Y(men_men_n302_));
  NAi31      u0274(.An(k), .B(l), .C(j), .Y(men_men_n303_));
  OAI210     u0275(.A0(men_men_n282_), .A1(j), .B0(men_men_n303_), .Y(men_men_n304_));
  NOi21      u0276(.An(men_men_n304_), .B(men_men_n120_), .Y(men_men_n305_));
  NA2        u0277(.A(men_men_n305_), .B(men_men_n302_), .Y(men_men_n306_));
  INV        u0278(.A(men_men_n306_), .Y(men_men_n307_));
  NO4        u0279(.A(men_men_n307_), .B(men_men_n297_), .C(men_men_n276_), .D(men_men_n270_), .Y(men_men_n308_));
  NA2        u0280(.A(men_men_n254_), .B(men_men_n193_), .Y(men_men_n309_));
  NAi21      u0281(.An(m), .B(k), .Y(men_men_n310_));
  NO2        u0282(.A(men_men_n225_), .B(men_men_n310_), .Y(men_men_n311_));
  NAi41      u0283(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n312_));
  NO2        u0284(.A(men_men_n312_), .B(men_men_n153_), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n313_), .B(men_men_n311_), .Y(men_men_n314_));
  NAi31      u0286(.An(i), .B(l), .C(h), .Y(men_men_n315_));
  NO4        u0287(.A(men_men_n315_), .B(men_men_n153_), .C(men_men_n69_), .D(men_men_n71_), .Y(men_men_n316_));
  NA2        u0288(.A(e), .B(c), .Y(men_men_n317_));
  NO3        u0289(.A(men_men_n317_), .B(n), .C(d), .Y(men_men_n318_));
  NOi21      u0290(.An(f), .B(h), .Y(men_men_n319_));
  NA2        u0291(.A(men_men_n319_), .B(men_men_n118_), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n320_), .B(men_men_n213_), .Y(men_men_n321_));
  NAi31      u0293(.An(d), .B(e), .C(b), .Y(men_men_n322_));
  NO2        u0294(.A(men_men_n133_), .B(men_men_n322_), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n323_), .B(men_men_n321_), .Y(men_men_n324_));
  NAi41      u0296(.An(men_men_n316_), .B(men_men_n324_), .C(men_men_n314_), .D(men_men_n309_), .Y(men_men_n325_));
  NO4        u0297(.A(men_men_n312_), .B(men_men_n77_), .C(men_men_n68_), .D(men_men_n213_), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n249_), .B(men_men_n103_), .Y(men_men_n327_));
  OR2        u0299(.A(men_men_n327_), .B(men_men_n205_), .Y(men_men_n328_));
  NOi31      u0300(.An(l), .B(n), .C(m), .Y(men_men_n329_));
  NA2        u0301(.A(men_men_n329_), .B(men_men_n214_), .Y(men_men_n330_));
  NO2        u0302(.A(men_men_n330_), .B(men_men_n194_), .Y(men_men_n331_));
  NAi32      u0303(.An(men_men_n331_), .Bn(men_men_n326_), .C(men_men_n328_), .Y(men_men_n332_));
  NAi32      u0304(.An(m), .Bn(j), .C(k), .Y(men_men_n333_));
  NAi41      u0305(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n334_));
  NOi31      u0306(.An(j), .B(m), .C(k), .Y(men_men_n335_));
  NO2        u0307(.A(men_men_n126_), .B(men_men_n335_), .Y(men_men_n336_));
  AN3        u0308(.A(h), .B(g), .C(f), .Y(men_men_n337_));
  NOi32      u0309(.An(m), .Bn(j), .C(l), .Y(men_men_n338_));
  NO2        u0310(.A(men_men_n338_), .B(men_men_n96_), .Y(men_men_n339_));
  NAi32      u0311(.An(men_men_n339_), .Bn(men_men_n202_), .C(men_men_n298_), .Y(men_men_n340_));
  NO2        u0312(.A(men_men_n291_), .B(men_men_n290_), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n216_), .B(g), .Y(men_men_n342_));
  NO2        u0314(.A(men_men_n159_), .B(men_men_n82_), .Y(men_men_n343_));
  AOI220     u0315(.A0(men_men_n343_), .A1(men_men_n342_), .B0(men_men_n246_), .B1(men_men_n341_), .Y(men_men_n344_));
  NA2        u0316(.A(men_men_n233_), .B(men_men_n77_), .Y(men_men_n345_));
  NA3        u0317(.A(men_men_n345_), .B(men_men_n337_), .C(men_men_n211_), .Y(men_men_n346_));
  NA3        u0318(.A(men_men_n346_), .B(men_men_n344_), .C(men_men_n340_), .Y(men_men_n347_));
  NA3        u0319(.A(h), .B(g), .C(f), .Y(men_men_n348_));
  NO2        u0320(.A(men_men_n348_), .B(men_men_n73_), .Y(men_men_n349_));
  NA2        u0321(.A(men_men_n334_), .B(men_men_n210_), .Y(men_men_n350_));
  NA2        u0322(.A(men_men_n166_), .B(e), .Y(men_men_n351_));
  NO2        u0323(.A(men_men_n351_), .B(men_men_n41_), .Y(men_men_n352_));
  AOI220     u0324(.A0(men_men_n352_), .A1(men_men_n302_), .B0(men_men_n350_), .B1(men_men_n349_), .Y(men_men_n353_));
  NOi32      u0325(.An(j), .Bn(g), .C(i), .Y(men_men_n354_));
  NA3        u0326(.A(men_men_n354_), .B(men_men_n282_), .C(men_men_n113_), .Y(men_men_n355_));
  OR2        u0327(.A(men_men_n111_), .B(men_men_n355_), .Y(men_men_n356_));
  NOi32      u0328(.An(e), .Bn(b), .C(a), .Y(men_men_n357_));
  AN2        u0329(.A(l), .B(j), .Y(men_men_n358_));
  NO2        u0330(.A(men_men_n310_), .B(men_men_n358_), .Y(men_men_n359_));
  NO3        u0331(.A(men_men_n312_), .B(men_men_n68_), .C(men_men_n213_), .Y(men_men_n360_));
  NA2        u0332(.A(men_men_n207_), .B(men_men_n35_), .Y(men_men_n361_));
  AOI220     u0333(.A0(men_men_n361_), .A1(men_men_n357_), .B0(men_men_n360_), .B1(men_men_n359_), .Y(men_men_n362_));
  NO2        u0334(.A(men_men_n322_), .B(n), .Y(men_men_n363_));
  NA2        u0335(.A(men_men_n206_), .B(k), .Y(men_men_n364_));
  NA3        u0336(.A(m), .B(men_men_n112_), .C(men_men_n212_), .Y(men_men_n365_));
  NO2        u0337(.A(men_men_n365_), .B(men_men_n364_), .Y(men_men_n366_));
  NAi41      u0338(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n367_));
  NA2        u0339(.A(men_men_n49_), .B(men_men_n113_), .Y(men_men_n368_));
  NO2        u0340(.A(men_men_n368_), .B(men_men_n367_), .Y(men_men_n369_));
  AOI220     u0341(.A0(men_men_n369_), .A1(b), .B0(men_men_n366_), .B1(men_men_n363_), .Y(men_men_n370_));
  NA4        u0342(.A(men_men_n370_), .B(men_men_n362_), .C(men_men_n356_), .D(men_men_n353_), .Y(men_men_n371_));
  NO4        u0343(.A(men_men_n371_), .B(men_men_n347_), .C(men_men_n332_), .D(men_men_n325_), .Y(men_men_n372_));
  NA4        u0344(.A(men_men_n372_), .B(men_men_n308_), .C(men_men_n268_), .D(men_men_n200_), .Y(men10));
  NA3        u0345(.A(m), .B(k), .C(i), .Y(men_men_n374_));
  NO3        u0346(.A(men_men_n374_), .B(j), .C(men_men_n213_), .Y(men_men_n375_));
  NOi21      u0347(.An(e), .B(f), .Y(men_men_n376_));
  NO4        u0348(.A(men_men_n154_), .B(men_men_n376_), .C(n), .D(men_men_n110_), .Y(men_men_n377_));
  NAi31      u0349(.An(b), .B(f), .C(c), .Y(men_men_n378_));
  INV        u0350(.A(men_men_n378_), .Y(men_men_n379_));
  NOi32      u0351(.An(k), .Bn(h), .C(j), .Y(men_men_n380_));
  NA2        u0352(.A(men_men_n380_), .B(men_men_n220_), .Y(men_men_n381_));
  NA2        u0353(.A(men_men_n164_), .B(men_men_n381_), .Y(men_men_n382_));
  AOI220     u0354(.A0(men_men_n382_), .A1(men_men_n379_), .B0(men_men_n377_), .B1(men_men_n375_), .Y(men_men_n383_));
  AN2        u0355(.A(j), .B(h), .Y(men_men_n384_));
  NO3        u0356(.A(n), .B(m), .C(k), .Y(men_men_n385_));
  NA2        u0357(.A(men_men_n385_), .B(men_men_n384_), .Y(men_men_n386_));
  NO3        u0358(.A(men_men_n386_), .B(men_men_n154_), .C(men_men_n212_), .Y(men_men_n387_));
  OR2        u0359(.A(m), .B(k), .Y(men_men_n388_));
  NO2        u0360(.A(men_men_n177_), .B(men_men_n388_), .Y(men_men_n389_));
  NA4        u0361(.A(n), .B(f), .C(c), .D(men_men_n116_), .Y(men_men_n390_));
  NOi21      u0362(.An(men_men_n389_), .B(men_men_n390_), .Y(men_men_n391_));
  NOi32      u0363(.An(d), .Bn(a), .C(c), .Y(men_men_n392_));
  NA2        u0364(.A(men_men_n392_), .B(men_men_n185_), .Y(men_men_n393_));
  NAi21      u0365(.An(i), .B(g), .Y(men_men_n394_));
  NAi31      u0366(.An(k), .B(m), .C(j), .Y(men_men_n395_));
  NO2        u0367(.A(men_men_n391_), .B(men_men_n387_), .Y(men_men_n396_));
  NO2        u0368(.A(men_men_n390_), .B(men_men_n291_), .Y(men_men_n397_));
  NOi32      u0369(.An(f), .Bn(d), .C(c), .Y(men_men_n398_));
  AOI220     u0370(.A0(men_men_n398_), .A1(men_men_n301_), .B0(men_men_n397_), .B1(men_men_n214_), .Y(men_men_n399_));
  NA3        u0371(.A(men_men_n399_), .B(men_men_n396_), .C(men_men_n383_), .Y(men_men_n400_));
  NO2        u0372(.A(men_men_n55_), .B(men_men_n116_), .Y(men_men_n401_));
  NA2        u0373(.A(men_men_n249_), .B(men_men_n401_), .Y(men_men_n402_));
  INV        u0374(.A(e), .Y(men_men_n403_));
  NA2        u0375(.A(men_men_n44_), .B(e), .Y(men_men_n404_));
  OAI220     u0376(.A0(men_men_n404_), .A1(men_men_n201_), .B0(men_men_n205_), .B1(men_men_n403_), .Y(men_men_n405_));
  AN2        u0377(.A(g), .B(e), .Y(men_men_n406_));
  NA3        u0378(.A(men_men_n406_), .B(men_men_n204_), .C(i), .Y(men_men_n407_));
  INV        u0379(.A(men_men_n407_), .Y(men_men_n408_));
  NO2        u0380(.A(men_men_n99_), .B(men_men_n403_), .Y(men_men_n409_));
  NO3        u0381(.A(men_men_n409_), .B(men_men_n408_), .C(men_men_n405_), .Y(men_men_n410_));
  NOi32      u0382(.An(h), .Bn(e), .C(g), .Y(men_men_n411_));
  NA3        u0383(.A(men_men_n411_), .B(men_men_n284_), .C(m), .Y(men_men_n412_));
  NOi21      u0384(.An(g), .B(h), .Y(men_men_n413_));
  AN3        u0385(.A(m), .B(l), .C(i), .Y(men_men_n414_));
  NA3        u0386(.A(men_men_n414_), .B(men_men_n413_), .C(e), .Y(men_men_n415_));
  AN3        u0387(.A(h), .B(g), .C(e), .Y(men_men_n416_));
  NA2        u0388(.A(men_men_n416_), .B(men_men_n96_), .Y(men_men_n417_));
  AN2        u0389(.A(men_men_n417_), .B(men_men_n415_), .Y(men_men_n418_));
  AOI210     u0390(.A0(men_men_n418_), .A1(men_men_n410_), .B0(men_men_n402_), .Y(men_men_n419_));
  NA3        u0391(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n420_));
  NO2        u0392(.A(men_men_n420_), .B(men_men_n402_), .Y(men_men_n421_));
  NAi31      u0393(.An(b), .B(c), .C(a), .Y(men_men_n422_));
  NO2        u0394(.A(men_men_n422_), .B(n), .Y(men_men_n423_));
  NA2        u0395(.A(men_men_n49_), .B(m), .Y(men_men_n424_));
  NO2        u0396(.A(men_men_n424_), .B(men_men_n150_), .Y(men_men_n425_));
  NA2        u0397(.A(men_men_n425_), .B(men_men_n423_), .Y(men_men_n426_));
  INV        u0398(.A(men_men_n426_), .Y(men_men_n427_));
  NO4        u0399(.A(men_men_n427_), .B(men_men_n421_), .C(men_men_n419_), .D(men_men_n400_), .Y(men_men_n428_));
  NA2        u0400(.A(i), .B(g), .Y(men_men_n429_));
  NO3        u0401(.A(men_men_n275_), .B(men_men_n429_), .C(c), .Y(men_men_n430_));
  NOi21      u0402(.An(a), .B(n), .Y(men_men_n431_));
  NOi21      u0403(.An(d), .B(c), .Y(men_men_n432_));
  NA2        u0404(.A(men_men_n432_), .B(men_men_n431_), .Y(men_men_n433_));
  NA3        u0405(.A(i), .B(g), .C(f), .Y(men_men_n434_));
  OR2        u0406(.A(men_men_n434_), .B(men_men_n67_), .Y(men_men_n435_));
  NA3        u0407(.A(men_men_n414_), .B(men_men_n413_), .C(men_men_n185_), .Y(men_men_n436_));
  AOI210     u0408(.A0(men_men_n436_), .A1(men_men_n435_), .B0(men_men_n433_), .Y(men_men_n437_));
  AOI210     u0409(.A0(men_men_n430_), .A1(men_men_n283_), .B0(men_men_n437_), .Y(men_men_n438_));
  OR2        u0410(.A(n), .B(m), .Y(men_men_n439_));
  NO2        u0411(.A(men_men_n439_), .B(men_men_n155_), .Y(men_men_n440_));
  NO2        u0412(.A(men_men_n186_), .B(men_men_n150_), .Y(men_men_n441_));
  OAI210     u0413(.A0(men_men_n440_), .A1(men_men_n179_), .B0(men_men_n441_), .Y(men_men_n442_));
  INV        u0414(.A(men_men_n368_), .Y(men_men_n443_));
  NA3        u0415(.A(men_men_n443_), .B(men_men_n357_), .C(d), .Y(men_men_n444_));
  NO2        u0416(.A(men_men_n422_), .B(men_men_n47_), .Y(men_men_n445_));
  NO3        u0417(.A(men_men_n62_), .B(men_men_n112_), .C(e), .Y(men_men_n446_));
  NAi21      u0418(.An(k), .B(j), .Y(men_men_n447_));
  NA2        u0419(.A(men_men_n252_), .B(men_men_n447_), .Y(men_men_n448_));
  NA3        u0420(.A(men_men_n448_), .B(men_men_n446_), .C(men_men_n445_), .Y(men_men_n449_));
  NAi21      u0421(.An(e), .B(d), .Y(men_men_n450_));
  INV        u0422(.A(men_men_n450_), .Y(men_men_n451_));
  NO2        u0423(.A(men_men_n253_), .B(men_men_n212_), .Y(men_men_n452_));
  NA3        u0424(.A(men_men_n452_), .B(men_men_n451_), .C(men_men_n226_), .Y(men_men_n453_));
  NA4        u0425(.A(men_men_n453_), .B(men_men_n449_), .C(men_men_n444_), .D(men_men_n442_), .Y(men_men_n454_));
  NO2        u0426(.A(men_men_n330_), .B(men_men_n212_), .Y(men_men_n455_));
  NA2        u0427(.A(men_men_n455_), .B(men_men_n451_), .Y(men_men_n456_));
  NOi31      u0428(.An(n), .B(m), .C(k), .Y(men_men_n457_));
  AOI220     u0429(.A0(men_men_n457_), .A1(men_men_n384_), .B0(men_men_n220_), .B1(men_men_n48_), .Y(men_men_n458_));
  NAi31      u0430(.An(g), .B(f), .C(c), .Y(men_men_n459_));
  INV        u0431(.A(men_men_n456_), .Y(men_men_n460_));
  NOi41      u0432(.An(men_men_n438_), .B(men_men_n460_), .C(men_men_n454_), .D(men_men_n266_), .Y(men_men_n461_));
  NOi32      u0433(.An(c), .Bn(a), .C(b), .Y(men_men_n462_));
  NA2        u0434(.A(men_men_n462_), .B(men_men_n113_), .Y(men_men_n463_));
  INV        u0435(.A(men_men_n274_), .Y(men_men_n464_));
  AN2        u0436(.A(e), .B(d), .Y(men_men_n465_));
  NA2        u0437(.A(men_men_n465_), .B(men_men_n464_), .Y(men_men_n466_));
  INV        u0438(.A(men_men_n150_), .Y(men_men_n467_));
  NO2        u0439(.A(men_men_n132_), .B(men_men_n41_), .Y(men_men_n468_));
  NO2        u0440(.A(men_men_n62_), .B(e), .Y(men_men_n469_));
  NA3        u0441(.A(men_men_n315_), .B(men_men_n168_), .C(men_men_n119_), .Y(men_men_n470_));
  AOI220     u0442(.A0(men_men_n470_), .A1(men_men_n469_), .B0(men_men_n468_), .B1(men_men_n467_), .Y(men_men_n471_));
  AOI210     u0443(.A0(men_men_n471_), .A1(men_men_n466_), .B0(men_men_n463_), .Y(men_men_n472_));
  NOi21      u0444(.An(a), .B(b), .Y(men_men_n473_));
  NA3        u0445(.A(e), .B(d), .C(c), .Y(men_men_n474_));
  NAi21      u0446(.An(men_men_n474_), .B(men_men_n473_), .Y(men_men_n475_));
  AOI210     u0447(.A0(men_men_n269_), .A1(men_men_n207_), .B0(men_men_n475_), .Y(men_men_n476_));
  NO4        u0448(.A(men_men_n190_), .B(men_men_n102_), .C(men_men_n52_), .D(b), .Y(men_men_n477_));
  NA2        u0449(.A(men_men_n379_), .B(men_men_n156_), .Y(men_men_n478_));
  OR2        u0450(.A(k), .B(j), .Y(men_men_n479_));
  NA2        u0451(.A(l), .B(k), .Y(men_men_n480_));
  NA3        u0452(.A(men_men_n480_), .B(men_men_n479_), .C(men_men_n220_), .Y(men_men_n481_));
  AOI210     u0453(.A0(men_men_n233_), .A1(men_men_n333_), .B0(men_men_n82_), .Y(men_men_n482_));
  NOi21      u0454(.An(men_men_n481_), .B(men_men_n482_), .Y(men_men_n483_));
  OR3        u0455(.A(men_men_n483_), .B(men_men_n146_), .C(men_men_n136_), .Y(men_men_n484_));
  NA2        u0456(.A(men_men_n129_), .B(men_men_n127_), .Y(men_men_n485_));
  NA2        u0457(.A(men_men_n392_), .B(men_men_n113_), .Y(men_men_n486_));
  NO4        u0458(.A(men_men_n486_), .B(men_men_n93_), .C(men_men_n112_), .D(e), .Y(men_men_n487_));
  NO3        u0459(.A(men_men_n487_), .B(men_men_n485_), .C(men_men_n316_), .Y(men_men_n488_));
  NA3        u0460(.A(men_men_n488_), .B(men_men_n484_), .C(men_men_n478_), .Y(men_men_n489_));
  NO4        u0461(.A(men_men_n489_), .B(men_men_n477_), .C(men_men_n476_), .D(men_men_n472_), .Y(men_men_n490_));
  NA2        u0462(.A(men_men_n66_), .B(men_men_n63_), .Y(men_men_n491_));
  NOi21      u0463(.An(d), .B(e), .Y(men_men_n492_));
  NO2        u0464(.A(men_men_n190_), .B(men_men_n52_), .Y(men_men_n493_));
  NAi31      u0465(.An(j), .B(l), .C(i), .Y(men_men_n494_));
  OAI210     u0466(.A0(men_men_n494_), .A1(men_men_n133_), .B0(men_men_n102_), .Y(men_men_n495_));
  NA3        u0467(.A(men_men_n495_), .B(men_men_n493_), .C(men_men_n492_), .Y(men_men_n496_));
  NO3        u0468(.A(men_men_n393_), .B(men_men_n339_), .C(men_men_n202_), .Y(men_men_n497_));
  NO2        u0469(.A(men_men_n393_), .B(men_men_n368_), .Y(men_men_n498_));
  NO3        u0470(.A(men_men_n498_), .B(men_men_n497_), .C(men_men_n299_), .Y(men_men_n499_));
  NA4        u0471(.A(men_men_n499_), .B(men_men_n496_), .C(men_men_n491_), .D(men_men_n243_), .Y(men_men_n500_));
  OAI210     u0472(.A0(men_men_n128_), .A1(men_men_n126_), .B0(n), .Y(men_men_n501_));
  NO2        u0473(.A(men_men_n501_), .B(men_men_n132_), .Y(men_men_n502_));
  OA210      u0474(.A0(men_men_n292_), .A1(men_men_n502_), .B0(men_men_n193_), .Y(men_men_n503_));
  XO2        u0475(.A(i), .B(h), .Y(men_men_n504_));
  NA3        u0476(.A(men_men_n504_), .B(men_men_n163_), .C(n), .Y(men_men_n505_));
  NAi41      u0477(.An(men_men_n292_), .B(men_men_n505_), .C(men_men_n458_), .D(men_men_n381_), .Y(men_men_n506_));
  NOi32      u0478(.An(men_men_n506_), .Bn(men_men_n469_), .C(men_men_n271_), .Y(men_men_n507_));
  NAi31      u0479(.An(c), .B(f), .C(d), .Y(men_men_n508_));
  AOI210     u0480(.A0(men_men_n277_), .A1(men_men_n196_), .B0(men_men_n508_), .Y(men_men_n509_));
  NOi21      u0481(.An(men_men_n80_), .B(men_men_n509_), .Y(men_men_n510_));
  NA3        u0482(.A(men_men_n377_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n511_));
  NA2        u0483(.A(men_men_n227_), .B(men_men_n108_), .Y(men_men_n512_));
  AOI210     u0484(.A0(men_men_n512_), .A1(men_men_n184_), .B0(men_men_n508_), .Y(men_men_n513_));
  AOI210     u0485(.A0(men_men_n355_), .A1(men_men_n35_), .B0(men_men_n475_), .Y(men_men_n514_));
  NOi31      u0486(.An(men_men_n511_), .B(men_men_n514_), .C(men_men_n513_), .Y(men_men_n515_));
  AN2        u0487(.A(men_men_n169_), .B(men_men_n63_), .Y(men_men_n516_));
  NA3        u0488(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n517_));
  INV        u0489(.A(men_men_n288_), .Y(men_men_n518_));
  NAi41      u0490(.An(men_men_n516_), .B(men_men_n518_), .C(men_men_n515_), .D(men_men_n510_), .Y(men_men_n519_));
  NO4        u0491(.A(men_men_n519_), .B(men_men_n507_), .C(men_men_n503_), .D(men_men_n500_), .Y(men_men_n520_));
  NA4        u0492(.A(men_men_n520_), .B(men_men_n490_), .C(men_men_n461_), .D(men_men_n428_), .Y(men11));
  NO2        u0493(.A(men_men_n69_), .B(f), .Y(men_men_n522_));
  NA2        u0494(.A(j), .B(g), .Y(men_men_n523_));
  NAi31      u0495(.An(i), .B(m), .C(l), .Y(men_men_n524_));
  NA3        u0496(.A(m), .B(k), .C(j), .Y(men_men_n525_));
  OAI220     u0497(.A0(men_men_n525_), .A1(men_men_n132_), .B0(men_men_n524_), .B1(men_men_n523_), .Y(men_men_n526_));
  NOi32      u0498(.An(e), .Bn(b), .C(f), .Y(men_men_n527_));
  NA2        u0499(.A(men_men_n259_), .B(men_men_n113_), .Y(men_men_n528_));
  NA2        u0500(.A(men_men_n44_), .B(j), .Y(men_men_n529_));
  NO2        u0501(.A(men_men_n529_), .B(men_men_n294_), .Y(men_men_n530_));
  NAi31      u0502(.An(d), .B(e), .C(a), .Y(men_men_n531_));
  NO2        u0503(.A(men_men_n531_), .B(n), .Y(men_men_n532_));
  AOI220     u0504(.A0(men_men_n532_), .A1(men_men_n100_), .B0(men_men_n530_), .B1(men_men_n527_), .Y(men_men_n533_));
  NAi41      u0505(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n534_));
  AN2        u0506(.A(men_men_n534_), .B(men_men_n367_), .Y(men_men_n535_));
  AOI210     u0507(.A0(men_men_n535_), .A1(men_men_n393_), .B0(men_men_n272_), .Y(men_men_n536_));
  NA2        u0508(.A(j), .B(i), .Y(men_men_n537_));
  NAi31      u0509(.An(n), .B(m), .C(k), .Y(men_men_n538_));
  NO3        u0510(.A(men_men_n538_), .B(men_men_n537_), .C(men_men_n112_), .Y(men_men_n539_));
  NO4        u0511(.A(n), .B(d), .C(men_men_n116_), .D(a), .Y(men_men_n540_));
  OR2        u0512(.A(n), .B(c), .Y(men_men_n541_));
  INV        u0513(.A(men_men_n540_), .Y(men_men_n542_));
  NOi32      u0514(.An(g), .Bn(f), .C(i), .Y(men_men_n543_));
  NA2        u0515(.A(men_men_n526_), .B(f), .Y(men_men_n544_));
  NO2        u0516(.A(men_men_n274_), .B(men_men_n47_), .Y(men_men_n545_));
  NO2        u0517(.A(men_men_n544_), .B(men_men_n542_), .Y(men_men_n546_));
  AOI210     u0518(.A0(men_men_n539_), .A1(men_men_n536_), .B0(men_men_n546_), .Y(men_men_n547_));
  NA2        u0519(.A(men_men_n142_), .B(men_men_n34_), .Y(men_men_n548_));
  OAI220     u0520(.A0(men_men_n548_), .A1(m), .B0(men_men_n529_), .B1(men_men_n233_), .Y(men_men_n549_));
  NOi41      u0521(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n550_));
  NAi32      u0522(.An(e), .Bn(b), .C(c), .Y(men_men_n551_));
  OR2        u0523(.A(men_men_n551_), .B(men_men_n82_), .Y(men_men_n552_));
  AN2        u0524(.A(men_men_n334_), .B(men_men_n312_), .Y(men_men_n553_));
  NA2        u0525(.A(men_men_n553_), .B(men_men_n552_), .Y(men_men_n554_));
  OA210      u0526(.A0(men_men_n554_), .A1(men_men_n550_), .B0(men_men_n549_), .Y(men_men_n555_));
  OAI220     u0527(.A0(men_men_n395_), .A1(men_men_n394_), .B0(men_men_n524_), .B1(men_men_n523_), .Y(men_men_n556_));
  NAi31      u0528(.An(d), .B(c), .C(a), .Y(men_men_n557_));
  NO2        u0529(.A(men_men_n557_), .B(n), .Y(men_men_n558_));
  NA3        u0530(.A(men_men_n558_), .B(men_men_n556_), .C(e), .Y(men_men_n559_));
  NO3        u0531(.A(men_men_n58_), .B(men_men_n47_), .C(men_men_n213_), .Y(men_men_n560_));
  NO2        u0532(.A(men_men_n230_), .B(men_men_n110_), .Y(men_men_n561_));
  NA2        u0533(.A(men_men_n560_), .B(men_men_n561_), .Y(men_men_n562_));
  NA2        u0534(.A(men_men_n562_), .B(men_men_n559_), .Y(men_men_n563_));
  NO2        u0535(.A(men_men_n275_), .B(n), .Y(men_men_n564_));
  NO2        u0536(.A(men_men_n423_), .B(men_men_n564_), .Y(men_men_n565_));
  NA2        u0537(.A(men_men_n556_), .B(f), .Y(men_men_n566_));
  NAi32      u0538(.An(d), .Bn(a), .C(b), .Y(men_men_n567_));
  NO2        u0539(.A(men_men_n567_), .B(men_men_n47_), .Y(men_men_n568_));
  NA2        u0540(.A(h), .B(f), .Y(men_men_n569_));
  NO2        u0541(.A(men_men_n569_), .B(men_men_n93_), .Y(men_men_n570_));
  NO3        u0542(.A(men_men_n180_), .B(men_men_n177_), .C(g), .Y(men_men_n571_));
  AOI220     u0543(.A0(men_men_n571_), .A1(men_men_n54_), .B0(men_men_n570_), .B1(men_men_n568_), .Y(men_men_n572_));
  OAI210     u0544(.A0(men_men_n566_), .A1(men_men_n565_), .B0(men_men_n572_), .Y(men_men_n573_));
  AN3        u0545(.A(j), .B(h), .C(g), .Y(men_men_n574_));
  NO2        u0546(.A(men_men_n149_), .B(c), .Y(men_men_n575_));
  NA3        u0547(.A(f), .B(d), .C(b), .Y(men_men_n576_));
  NO4        u0548(.A(men_men_n576_), .B(men_men_n180_), .C(men_men_n177_), .D(g), .Y(men_men_n577_));
  NO4        u0549(.A(men_men_n577_), .B(men_men_n573_), .C(men_men_n563_), .D(men_men_n555_), .Y(men_men_n578_));
  AN3        u0550(.A(men_men_n578_), .B(men_men_n547_), .C(men_men_n533_), .Y(men_men_n579_));
  INV        u0551(.A(k), .Y(men_men_n580_));
  NA3        u0552(.A(l), .B(men_men_n580_), .C(i), .Y(men_men_n581_));
  INV        u0553(.A(men_men_n581_), .Y(men_men_n582_));
  NA4        u0554(.A(men_men_n392_), .B(men_men_n413_), .C(men_men_n185_), .D(men_men_n113_), .Y(men_men_n583_));
  NAi32      u0555(.An(h), .Bn(f), .C(g), .Y(men_men_n584_));
  NAi41      u0556(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n585_));
  OAI210     u0557(.A0(men_men_n531_), .A1(n), .B0(men_men_n585_), .Y(men_men_n586_));
  NA2        u0558(.A(men_men_n586_), .B(m), .Y(men_men_n587_));
  NAi31      u0559(.An(h), .B(g), .C(f), .Y(men_men_n588_));
  OR3        u0560(.A(men_men_n588_), .B(men_men_n275_), .C(men_men_n47_), .Y(men_men_n589_));
  NA4        u0561(.A(men_men_n413_), .B(men_men_n121_), .C(men_men_n113_), .D(e), .Y(men_men_n590_));
  AN2        u0562(.A(men_men_n590_), .B(men_men_n589_), .Y(men_men_n591_));
  OA210      u0563(.A0(men_men_n587_), .A1(men_men_n584_), .B0(men_men_n591_), .Y(men_men_n592_));
  NA2        u0564(.A(men_men_n592_), .B(men_men_n583_), .Y(men_men_n593_));
  NAi31      u0565(.An(f), .B(h), .C(g), .Y(men_men_n594_));
  NO4        u0566(.A(men_men_n303_), .B(men_men_n594_), .C(men_men_n69_), .D(men_men_n71_), .Y(men_men_n595_));
  NOi32      u0567(.An(b), .Bn(a), .C(c), .Y(men_men_n596_));
  NOi41      u0568(.An(men_men_n596_), .B(men_men_n348_), .C(men_men_n65_), .D(men_men_n117_), .Y(men_men_n597_));
  OR2        u0569(.A(men_men_n597_), .B(men_men_n595_), .Y(men_men_n598_));
  NOi32      u0570(.An(d), .Bn(a), .C(e), .Y(men_men_n599_));
  NA2        u0571(.A(men_men_n599_), .B(men_men_n113_), .Y(men_men_n600_));
  NO2        u0572(.A(n), .B(c), .Y(men_men_n601_));
  NAi32      u0573(.An(n), .Bn(f), .C(m), .Y(men_men_n602_));
  NOi32      u0574(.An(e), .Bn(a), .C(d), .Y(men_men_n603_));
  AOI210     u0575(.A0(men_men_n29_), .A1(d), .B0(men_men_n603_), .Y(men_men_n604_));
  NO2        u0576(.A(men_men_n604_), .B(men_men_n548_), .Y(men_men_n605_));
  AOI210     u0577(.A0(men_men_n605_), .A1(men_men_n113_), .B0(men_men_n598_), .Y(men_men_n606_));
  OAI210     u0578(.A0(men_men_n248_), .A1(men_men_n85_), .B0(men_men_n606_), .Y(men_men_n607_));
  AOI210     u0579(.A0(men_men_n593_), .A1(men_men_n582_), .B0(men_men_n607_), .Y(men_men_n608_));
  NO3        u0580(.A(men_men_n310_), .B(men_men_n57_), .C(n), .Y(men_men_n609_));
  NA3        u0581(.A(men_men_n508_), .B(men_men_n175_), .C(men_men_n174_), .Y(men_men_n610_));
  NA2        u0582(.A(men_men_n459_), .B(men_men_n230_), .Y(men_men_n611_));
  OR2        u0583(.A(men_men_n611_), .B(men_men_n610_), .Y(men_men_n612_));
  NA2        u0584(.A(men_men_n72_), .B(men_men_n113_), .Y(men_men_n613_));
  NO2        u0585(.A(men_men_n613_), .B(men_men_n43_), .Y(men_men_n614_));
  AOI220     u0586(.A0(men_men_n614_), .A1(men_men_n536_), .B0(men_men_n612_), .B1(men_men_n609_), .Y(men_men_n615_));
  NO2        u0587(.A(men_men_n615_), .B(men_men_n85_), .Y(men_men_n616_));
  NA3        u0588(.A(men_men_n550_), .B(men_men_n335_), .C(men_men_n44_), .Y(men_men_n617_));
  NOi32      u0589(.An(e), .Bn(c), .C(f), .Y(men_men_n618_));
  NOi21      u0590(.An(f), .B(g), .Y(men_men_n619_));
  NO2        u0591(.A(men_men_n619_), .B(men_men_n210_), .Y(men_men_n620_));
  AOI220     u0592(.A0(men_men_n620_), .A1(men_men_n389_), .B0(men_men_n618_), .B1(men_men_n179_), .Y(men_men_n621_));
  NA3        u0593(.A(men_men_n621_), .B(men_men_n617_), .C(men_men_n182_), .Y(men_men_n622_));
  AOI210     u0594(.A0(men_men_n535_), .A1(men_men_n393_), .B0(men_men_n293_), .Y(men_men_n623_));
  NA2        u0595(.A(men_men_n623_), .B(men_men_n264_), .Y(men_men_n624_));
  NOi21      u0596(.An(j), .B(l), .Y(men_men_n625_));
  NAi21      u0597(.An(k), .B(h), .Y(men_men_n626_));
  NO2        u0598(.A(men_men_n626_), .B(men_men_n262_), .Y(men_men_n627_));
  NA2        u0599(.A(men_men_n627_), .B(men_men_n625_), .Y(men_men_n628_));
  OR2        u0600(.A(men_men_n628_), .B(men_men_n587_), .Y(men_men_n629_));
  NOi31      u0601(.An(m), .B(n), .C(k), .Y(men_men_n630_));
  NA2        u0602(.A(men_men_n625_), .B(men_men_n630_), .Y(men_men_n631_));
  NO2        u0603(.A(men_men_n275_), .B(men_men_n47_), .Y(men_men_n632_));
  NO2        u0604(.A(men_men_n303_), .B(men_men_n594_), .Y(men_men_n633_));
  NO2        u0605(.A(men_men_n531_), .B(men_men_n47_), .Y(men_men_n634_));
  AOI220     u0606(.A0(men_men_n634_), .A1(men_men_n633_), .B0(men_men_n632_), .B1(men_men_n570_), .Y(men_men_n635_));
  NA3        u0607(.A(men_men_n635_), .B(men_men_n629_), .C(men_men_n624_), .Y(men_men_n636_));
  NA2        u0608(.A(men_men_n108_), .B(men_men_n36_), .Y(men_men_n637_));
  NO2        u0609(.A(k), .B(men_men_n213_), .Y(men_men_n638_));
  NO2        u0610(.A(men_men_n527_), .B(men_men_n357_), .Y(men_men_n639_));
  NO2        u0611(.A(men_men_n639_), .B(n), .Y(men_men_n640_));
  NAi31      u0612(.An(men_men_n637_), .B(men_men_n640_), .C(men_men_n638_), .Y(men_men_n641_));
  NO2        u0613(.A(men_men_n529_), .B(men_men_n180_), .Y(men_men_n642_));
  NA3        u0614(.A(men_men_n551_), .B(men_men_n271_), .C(men_men_n147_), .Y(men_men_n643_));
  NA2        u0615(.A(men_men_n504_), .B(men_men_n163_), .Y(men_men_n644_));
  NO3        u0616(.A(men_men_n390_), .B(men_men_n644_), .C(men_men_n85_), .Y(men_men_n645_));
  AOI210     u0617(.A0(men_men_n643_), .A1(men_men_n642_), .B0(men_men_n645_), .Y(men_men_n646_));
  AN3        u0618(.A(f), .B(d), .C(b), .Y(men_men_n647_));
  OAI210     u0619(.A0(men_men_n647_), .A1(men_men_n131_), .B0(n), .Y(men_men_n648_));
  NA3        u0620(.A(men_men_n504_), .B(men_men_n163_), .C(men_men_n213_), .Y(men_men_n649_));
  AOI210     u0621(.A0(men_men_n648_), .A1(men_men_n232_), .B0(men_men_n649_), .Y(men_men_n650_));
  NAi31      u0622(.An(m), .B(n), .C(k), .Y(men_men_n651_));
  OR2        u0623(.A(men_men_n136_), .B(men_men_n57_), .Y(men_men_n652_));
  OAI210     u0624(.A0(men_men_n652_), .A1(men_men_n651_), .B0(men_men_n250_), .Y(men_men_n653_));
  OAI210     u0625(.A0(men_men_n653_), .A1(men_men_n650_), .B0(j), .Y(men_men_n654_));
  NA3        u0626(.A(men_men_n654_), .B(men_men_n646_), .C(men_men_n641_), .Y(men_men_n655_));
  NO4        u0627(.A(men_men_n655_), .B(men_men_n636_), .C(men_men_n622_), .D(men_men_n616_), .Y(men_men_n656_));
  NA2        u0628(.A(men_men_n377_), .B(men_men_n166_), .Y(men_men_n657_));
  NAi31      u0629(.An(g), .B(h), .C(f), .Y(men_men_n658_));
  OA210      u0630(.A0(men_men_n531_), .A1(n), .B0(men_men_n585_), .Y(men_men_n659_));
  NO2        u0631(.A(men_men_n659_), .B(men_men_n89_), .Y(men_men_n660_));
  INV        u0632(.A(men_men_n660_), .Y(men_men_n661_));
  AOI210     u0633(.A0(men_men_n661_), .A1(men_men_n657_), .B0(men_men_n525_), .Y(men_men_n662_));
  NO3        u0634(.A(g), .B(men_men_n212_), .C(men_men_n52_), .Y(men_men_n663_));
  NAi21      u0635(.An(h), .B(j), .Y(men_men_n664_));
  NO2        u0636(.A(men_men_n512_), .B(men_men_n85_), .Y(men_men_n665_));
  OAI210     u0637(.A0(men_men_n665_), .A1(men_men_n389_), .B0(men_men_n663_), .Y(men_men_n666_));
  OR2        u0638(.A(men_men_n69_), .B(men_men_n71_), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n596_), .B(men_men_n337_), .Y(men_men_n668_));
  OA220      u0640(.A0(men_men_n631_), .A1(men_men_n668_), .B0(men_men_n628_), .B1(men_men_n667_), .Y(men_men_n669_));
  NA3        u0641(.A(men_men_n522_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n670_));
  AN2        u0642(.A(h), .B(f), .Y(men_men_n671_));
  NA2        u0643(.A(men_men_n671_), .B(men_men_n37_), .Y(men_men_n672_));
  NA2        u0644(.A(men_men_n98_), .B(men_men_n44_), .Y(men_men_n673_));
  OAI220     u0645(.A0(men_men_n673_), .A1(men_men_n327_), .B0(men_men_n672_), .B1(men_men_n463_), .Y(men_men_n674_));
  AOI210     u0646(.A0(men_men_n567_), .A1(men_men_n422_), .B0(men_men_n47_), .Y(men_men_n675_));
  OAI220     u0647(.A0(men_men_n588_), .A1(men_men_n581_), .B0(men_men_n320_), .B1(men_men_n523_), .Y(men_men_n676_));
  AOI210     u0648(.A0(men_men_n676_), .A1(men_men_n675_), .B0(men_men_n674_), .Y(men_men_n677_));
  NA4        u0649(.A(men_men_n677_), .B(men_men_n670_), .C(men_men_n669_), .D(men_men_n666_), .Y(men_men_n678_));
  NO2        u0650(.A(men_men_n252_), .B(f), .Y(men_men_n679_));
  NO2        u0651(.A(men_men_n619_), .B(men_men_n57_), .Y(men_men_n680_));
  NO3        u0652(.A(men_men_n680_), .B(men_men_n679_), .C(men_men_n34_), .Y(men_men_n681_));
  NA2        u0653(.A(men_men_n323_), .B(men_men_n142_), .Y(men_men_n682_));
  NA2        u0654(.A(men_men_n133_), .B(men_men_n47_), .Y(men_men_n683_));
  NA2        u0655(.A(men_men_n357_), .B(men_men_n113_), .Y(men_men_n684_));
  OA220      u0656(.A0(men_men_n684_), .A1(men_men_n548_), .B0(men_men_n355_), .B1(men_men_n111_), .Y(men_men_n685_));
  OAI210     u0657(.A0(men_men_n682_), .A1(men_men_n681_), .B0(men_men_n685_), .Y(men_men_n686_));
  NO3        u0658(.A(men_men_n398_), .B(men_men_n193_), .C(men_men_n192_), .Y(men_men_n687_));
  NA2        u0659(.A(men_men_n687_), .B(men_men_n230_), .Y(men_men_n688_));
  NA3        u0660(.A(men_men_n688_), .B(men_men_n254_), .C(j), .Y(men_men_n689_));
  NO3        u0661(.A(men_men_n459_), .B(men_men_n177_), .C(i), .Y(men_men_n690_));
  NA2        u0662(.A(men_men_n462_), .B(men_men_n82_), .Y(men_men_n691_));
  NO4        u0663(.A(men_men_n525_), .B(men_men_n691_), .C(men_men_n132_), .D(men_men_n212_), .Y(men_men_n692_));
  INV        u0664(.A(men_men_n692_), .Y(men_men_n693_));
  NA4        u0665(.A(men_men_n693_), .B(men_men_n689_), .C(men_men_n511_), .D(men_men_n396_), .Y(men_men_n694_));
  NO4        u0666(.A(men_men_n694_), .B(men_men_n686_), .C(men_men_n678_), .D(men_men_n662_), .Y(men_men_n695_));
  NA4        u0667(.A(men_men_n695_), .B(men_men_n656_), .C(men_men_n608_), .D(men_men_n579_), .Y(men08));
  NO2        u0668(.A(k), .B(h), .Y(men_men_n697_));
  AO210      u0669(.A0(men_men_n252_), .A1(men_men_n447_), .B0(men_men_n697_), .Y(men_men_n698_));
  NO2        u0670(.A(men_men_n698_), .B(men_men_n291_), .Y(men_men_n699_));
  NA2        u0671(.A(men_men_n618_), .B(men_men_n82_), .Y(men_men_n700_));
  NA2        u0672(.A(men_men_n700_), .B(men_men_n459_), .Y(men_men_n701_));
  NA2        u0673(.A(men_men_n701_), .B(men_men_n699_), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n82_), .B(men_men_n110_), .Y(men_men_n703_));
  NO2        u0675(.A(men_men_n703_), .B(men_men_n53_), .Y(men_men_n704_));
  NA2        u0676(.A(men_men_n576_), .B(men_men_n232_), .Y(men_men_n705_));
  NA2        u0677(.A(men_men_n705_), .B(men_men_n342_), .Y(men_men_n706_));
  AOI210     u0678(.A0(men_men_n576_), .A1(men_men_n159_), .B0(men_men_n82_), .Y(men_men_n707_));
  NA4        u0679(.A(men_men_n215_), .B(men_men_n142_), .C(men_men_n43_), .D(h), .Y(men_men_n708_));
  AN2        u0680(.A(l), .B(k), .Y(men_men_n709_));
  NA3        u0681(.A(men_men_n706_), .B(men_men_n702_), .C(men_men_n344_), .Y(men_men_n710_));
  AN2        u0682(.A(men_men_n532_), .B(men_men_n94_), .Y(men_men_n711_));
  NO4        u0683(.A(men_men_n177_), .B(men_men_n388_), .C(men_men_n112_), .D(g), .Y(men_men_n712_));
  NA2        u0684(.A(men_men_n712_), .B(men_men_n705_), .Y(men_men_n713_));
  NO2        u0685(.A(men_men_n38_), .B(men_men_n212_), .Y(men_men_n714_));
  AOI220     u0686(.A0(men_men_n620_), .A1(men_men_n341_), .B0(men_men_n714_), .B1(men_men_n564_), .Y(men_men_n715_));
  NAi31      u0687(.An(men_men_n711_), .B(men_men_n715_), .C(men_men_n713_), .Y(men_men_n716_));
  NO2        u0688(.A(men_men_n535_), .B(men_men_n35_), .Y(men_men_n717_));
  OAI210     u0689(.A0(men_men_n551_), .A1(men_men_n45_), .B0(men_men_n652_), .Y(men_men_n718_));
  NO2        u0690(.A(men_men_n480_), .B(men_men_n133_), .Y(men_men_n719_));
  AOI210     u0691(.A0(men_men_n719_), .A1(men_men_n718_), .B0(men_men_n717_), .Y(men_men_n720_));
  NO3        u0692(.A(men_men_n310_), .B(men_men_n132_), .C(men_men_n41_), .Y(men_men_n721_));
  BUFFER     u0693(.A(men_men_n721_), .Y(men_men_n722_));
  NA2        u0694(.A(men_men_n698_), .B(men_men_n137_), .Y(men_men_n723_));
  AOI220     u0695(.A0(men_men_n723_), .A1(men_men_n397_), .B0(men_men_n722_), .B1(men_men_n74_), .Y(men_men_n724_));
  OAI210     u0696(.A0(men_men_n720_), .A1(men_men_n85_), .B0(men_men_n724_), .Y(men_men_n725_));
  NA3        u0697(.A(men_men_n688_), .B(men_men_n329_), .C(men_men_n380_), .Y(men_men_n726_));
  NA2        u0698(.A(men_men_n709_), .B(men_men_n220_), .Y(men_men_n727_));
  NO2        u0699(.A(men_men_n727_), .B(men_men_n322_), .Y(men_men_n728_));
  AOI210     u0700(.A0(men_men_n728_), .A1(men_men_n679_), .B0(men_men_n487_), .Y(men_men_n729_));
  NA3        u0701(.A(m), .B(l), .C(k), .Y(men_men_n730_));
  NO2        u0702(.A(men_men_n534_), .B(men_men_n272_), .Y(men_men_n731_));
  NOi21      u0703(.An(men_men_n731_), .B(men_men_n528_), .Y(men_men_n732_));
  NA4        u0704(.A(men_men_n113_), .B(l), .C(k), .D(men_men_n85_), .Y(men_men_n733_));
  NA3        u0705(.A(men_men_n121_), .B(men_men_n406_), .C(i), .Y(men_men_n734_));
  NO2        u0706(.A(men_men_n734_), .B(men_men_n733_), .Y(men_men_n735_));
  NO2        u0707(.A(men_men_n735_), .B(men_men_n732_), .Y(men_men_n736_));
  NA3        u0708(.A(men_men_n736_), .B(men_men_n729_), .C(men_men_n726_), .Y(men_men_n737_));
  NO4        u0709(.A(men_men_n737_), .B(men_men_n725_), .C(men_men_n716_), .D(men_men_n710_), .Y(men_men_n738_));
  NA2        u0710(.A(men_men_n620_), .B(men_men_n389_), .Y(men_men_n739_));
  NOi31      u0711(.An(g), .B(h), .C(f), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n634_), .B(men_men_n740_), .Y(men_men_n741_));
  AO210      u0713(.A0(men_men_n741_), .A1(men_men_n589_), .B0(men_men_n537_), .Y(men_men_n742_));
  NO3        u0714(.A(men_men_n393_), .B(men_men_n523_), .C(h), .Y(men_men_n743_));
  AOI210     u0715(.A0(men_men_n743_), .A1(men_men_n113_), .B0(men_men_n498_), .Y(men_men_n744_));
  NA4        u0716(.A(men_men_n744_), .B(men_men_n742_), .C(men_men_n739_), .D(men_men_n251_), .Y(men_men_n745_));
  NA2        u0717(.A(men_men_n709_), .B(men_men_n71_), .Y(men_men_n746_));
  NO4        u0718(.A(men_men_n687_), .B(men_men_n177_), .C(n), .D(i), .Y(men_men_n747_));
  NOi21      u0719(.An(h), .B(j), .Y(men_men_n748_));
  NA2        u0720(.A(men_men_n748_), .B(f), .Y(men_men_n749_));
  NO2        u0721(.A(men_men_n749_), .B(men_men_n245_), .Y(men_men_n750_));
  NO3        u0722(.A(men_men_n750_), .B(men_men_n747_), .C(men_men_n690_), .Y(men_men_n751_));
  OAI220     u0723(.A0(men_men_n751_), .A1(men_men_n746_), .B0(men_men_n591_), .B1(men_men_n58_), .Y(men_men_n752_));
  AOI210     u0724(.A0(men_men_n745_), .A1(l), .B0(men_men_n752_), .Y(men_men_n753_));
  NO2        u0725(.A(j), .B(i), .Y(men_men_n754_));
  NA3        u0726(.A(men_men_n754_), .B(men_men_n78_), .C(l), .Y(men_men_n755_));
  NA2        u0727(.A(men_men_n754_), .B(men_men_n33_), .Y(men_men_n756_));
  NA2        u0728(.A(men_men_n416_), .B(men_men_n121_), .Y(men_men_n757_));
  OA220      u0729(.A0(men_men_n757_), .A1(men_men_n756_), .B0(men_men_n755_), .B1(men_men_n587_), .Y(men_men_n758_));
  NO3        u0730(.A(men_men_n154_), .B(men_men_n47_), .C(men_men_n110_), .Y(men_men_n759_));
  NO3        u0731(.A(men_men_n541_), .B(men_men_n152_), .C(men_men_n71_), .Y(men_men_n760_));
  NO3        u0732(.A(men_men_n480_), .B(men_men_n434_), .C(j), .Y(men_men_n761_));
  OAI210     u0733(.A0(men_men_n760_), .A1(men_men_n759_), .B0(men_men_n761_), .Y(men_men_n762_));
  OAI210     u0734(.A0(men_men_n741_), .A1(men_men_n58_), .B0(men_men_n762_), .Y(men_men_n763_));
  NA2        u0735(.A(k), .B(j), .Y(men_men_n764_));
  NO3        u0736(.A(men_men_n291_), .B(men_men_n764_), .C(men_men_n40_), .Y(men_men_n765_));
  AOI210     u0737(.A0(men_men_n527_), .A1(n), .B0(men_men_n550_), .Y(men_men_n766_));
  NA2        u0738(.A(men_men_n766_), .B(men_men_n553_), .Y(men_men_n767_));
  AN3        u0739(.A(men_men_n767_), .B(men_men_n765_), .C(men_men_n97_), .Y(men_men_n768_));
  NO3        u0740(.A(men_men_n177_), .B(men_men_n388_), .C(men_men_n112_), .Y(men_men_n769_));
  AOI220     u0741(.A0(men_men_n769_), .A1(men_men_n246_), .B0(men_men_n611_), .B1(men_men_n301_), .Y(men_men_n770_));
  NAi31      u0742(.An(men_men_n604_), .B(men_men_n91_), .C(men_men_n82_), .Y(men_men_n771_));
  NA2        u0743(.A(men_men_n771_), .B(men_men_n770_), .Y(men_men_n772_));
  NO2        u0744(.A(men_men_n291_), .B(men_men_n137_), .Y(men_men_n773_));
  AOI220     u0745(.A0(men_men_n773_), .A1(men_men_n620_), .B0(men_men_n721_), .B1(men_men_n707_), .Y(men_men_n774_));
  NO2        u0746(.A(men_men_n730_), .B(men_men_n89_), .Y(men_men_n775_));
  NA2        u0747(.A(men_men_n775_), .B(men_men_n586_), .Y(men_men_n776_));
  NO2        u0748(.A(men_men_n588_), .B(men_men_n117_), .Y(men_men_n777_));
  OAI210     u0749(.A0(men_men_n777_), .A1(men_men_n761_), .B0(men_men_n675_), .Y(men_men_n778_));
  NA3        u0750(.A(men_men_n778_), .B(men_men_n776_), .C(men_men_n774_), .Y(men_men_n779_));
  OR4        u0751(.A(men_men_n779_), .B(men_men_n772_), .C(men_men_n768_), .D(men_men_n763_), .Y(men_men_n780_));
  NA3        u0752(.A(men_men_n766_), .B(men_men_n553_), .C(men_men_n552_), .Y(men_men_n781_));
  NA4        u0753(.A(men_men_n781_), .B(men_men_n215_), .C(men_men_n447_), .D(men_men_n34_), .Y(men_men_n782_));
  NO4        u0754(.A(men_men_n480_), .B(men_men_n429_), .C(j), .D(f), .Y(men_men_n783_));
  OAI220     u0755(.A0(men_men_n708_), .A1(men_men_n700_), .B0(men_men_n327_), .B1(men_men_n38_), .Y(men_men_n784_));
  AOI210     u0756(.A0(men_men_n783_), .A1(men_men_n258_), .B0(men_men_n784_), .Y(men_men_n785_));
  NA3        u0757(.A(men_men_n543_), .B(men_men_n284_), .C(h), .Y(men_men_n786_));
  NOi21      u0758(.An(men_men_n675_), .B(men_men_n786_), .Y(men_men_n787_));
  NO2        u0759(.A(men_men_n90_), .B(men_men_n45_), .Y(men_men_n788_));
  NO2        u0760(.A(men_men_n755_), .B(men_men_n667_), .Y(men_men_n789_));
  AOI210     u0761(.A0(men_men_n788_), .A1(men_men_n640_), .B0(men_men_n789_), .Y(men_men_n790_));
  NAi41      u0762(.An(men_men_n787_), .B(men_men_n790_), .C(men_men_n785_), .D(men_men_n782_), .Y(men_men_n791_));
  BUFFER     u0763(.A(men_men_n94_), .Y(men_men_n792_));
  AOI220     u0764(.A0(men_men_n792_), .A1(men_men_n238_), .B0(men_men_n761_), .B1(men_men_n632_), .Y(men_men_n793_));
  NO2        u0765(.A(men_men_n659_), .B(men_men_n71_), .Y(men_men_n794_));
  AOI210     u0766(.A0(men_men_n783_), .A1(men_men_n794_), .B0(men_men_n331_), .Y(men_men_n795_));
  OAI210     u0767(.A0(men_men_n730_), .A1(men_men_n658_), .B0(men_men_n517_), .Y(men_men_n796_));
  NA3        u0768(.A(men_men_n249_), .B(men_men_n55_), .C(b), .Y(men_men_n797_));
  AOI220     u0769(.A0(men_men_n601_), .A1(men_men_n29_), .B0(men_men_n462_), .B1(men_men_n82_), .Y(men_men_n798_));
  NA2        u0770(.A(men_men_n798_), .B(men_men_n797_), .Y(men_men_n799_));
  NO2        u0771(.A(men_men_n786_), .B(men_men_n486_), .Y(men_men_n800_));
  AOI210     u0772(.A0(men_men_n799_), .A1(men_men_n796_), .B0(men_men_n800_), .Y(men_men_n801_));
  NA3        u0773(.A(men_men_n801_), .B(men_men_n795_), .C(men_men_n793_), .Y(men_men_n802_));
  NOi41      u0774(.An(men_men_n758_), .B(men_men_n802_), .C(men_men_n791_), .D(men_men_n780_), .Y(men_men_n803_));
  OR3        u0775(.A(men_men_n708_), .B(men_men_n232_), .C(g), .Y(men_men_n804_));
  NO3        u0776(.A(men_men_n336_), .B(men_men_n293_), .C(men_men_n112_), .Y(men_men_n805_));
  NA2        u0777(.A(men_men_n805_), .B(men_men_n767_), .Y(men_men_n806_));
  NA2        u0778(.A(men_men_n44_), .B(men_men_n52_), .Y(men_men_n807_));
  NO3        u0779(.A(men_men_n807_), .B(men_men_n756_), .C(men_men_n275_), .Y(men_men_n808_));
  NO3        u0780(.A(men_men_n523_), .B(men_men_n92_), .C(h), .Y(men_men_n809_));
  AOI210     u0781(.A0(men_men_n809_), .A1(men_men_n704_), .B0(men_men_n808_), .Y(men_men_n810_));
  NA4        u0782(.A(men_men_n810_), .B(men_men_n806_), .C(men_men_n804_), .D(men_men_n399_), .Y(men_men_n811_));
  OR2        u0783(.A(men_men_n658_), .B(men_men_n90_), .Y(men_men_n812_));
  NOi31      u0784(.An(b), .B(d), .C(a), .Y(men_men_n813_));
  NO2        u0785(.A(men_men_n813_), .B(men_men_n599_), .Y(men_men_n814_));
  NO2        u0786(.A(men_men_n814_), .B(n), .Y(men_men_n815_));
  NOi21      u0787(.An(men_men_n798_), .B(men_men_n815_), .Y(men_men_n816_));
  OAI220     u0788(.A0(men_men_n816_), .A1(men_men_n812_), .B0(men_men_n786_), .B1(men_men_n600_), .Y(men_men_n817_));
  NO2        u0789(.A(men_men_n551_), .B(men_men_n82_), .Y(men_men_n818_));
  NO3        u0790(.A(men_men_n619_), .B(men_men_n322_), .C(men_men_n117_), .Y(men_men_n819_));
  NOi21      u0791(.An(men_men_n819_), .B(men_men_n164_), .Y(men_men_n820_));
  AOI210     u0792(.A0(men_men_n805_), .A1(men_men_n818_), .B0(men_men_n820_), .Y(men_men_n821_));
  OAI210     u0793(.A0(men_men_n708_), .A1(men_men_n390_), .B0(men_men_n821_), .Y(men_men_n822_));
  NO2        u0794(.A(men_men_n687_), .B(n), .Y(men_men_n823_));
  AOI220     u0795(.A0(men_men_n773_), .A1(men_men_n663_), .B0(men_men_n823_), .B1(men_men_n699_), .Y(men_men_n824_));
  NO2        u0796(.A(men_men_n317_), .B(men_men_n237_), .Y(men_men_n825_));
  OAI210     u0797(.A0(men_men_n94_), .A1(men_men_n91_), .B0(men_men_n825_), .Y(men_men_n826_));
  NA2        u0798(.A(men_men_n121_), .B(men_men_n82_), .Y(men_men_n827_));
  AOI210     u0799(.A0(men_men_n420_), .A1(men_men_n412_), .B0(men_men_n827_), .Y(men_men_n828_));
  NAi21      u0800(.An(men_men_n828_), .B(men_men_n826_), .Y(men_men_n829_));
  NA2        u0801(.A(men_men_n728_), .B(men_men_n34_), .Y(men_men_n830_));
  NAi21      u0802(.An(men_men_n733_), .B(men_men_n430_), .Y(men_men_n831_));
  NO2        u0803(.A(men_men_n272_), .B(i), .Y(men_men_n832_));
  NA2        u0804(.A(men_men_n712_), .B(men_men_n343_), .Y(men_men_n833_));
  AN2        u0805(.A(men_men_n833_), .B(men_men_n831_), .Y(men_men_n834_));
  NAi41      u0806(.An(men_men_n829_), .B(men_men_n834_), .C(men_men_n830_), .D(men_men_n824_), .Y(men_men_n835_));
  NO4        u0807(.A(men_men_n835_), .B(men_men_n822_), .C(men_men_n817_), .D(men_men_n811_), .Y(men_men_n836_));
  NA4        u0808(.A(men_men_n836_), .B(men_men_n803_), .C(men_men_n753_), .D(men_men_n738_), .Y(men09));
  INV        u0809(.A(men_men_n122_), .Y(men_men_n838_));
  NA2        u0810(.A(f), .B(e), .Y(men_men_n839_));
  NO2        u0811(.A(men_men_n225_), .B(men_men_n112_), .Y(men_men_n840_));
  NA2        u0812(.A(men_men_n840_), .B(g), .Y(men_men_n841_));
  NA4        u0813(.A(men_men_n303_), .B(men_men_n168_), .C(men_men_n260_), .D(men_men_n119_), .Y(men_men_n842_));
  AOI210     u0814(.A0(men_men_n842_), .A1(g), .B0(men_men_n468_), .Y(men_men_n843_));
  AOI210     u0815(.A0(men_men_n843_), .A1(men_men_n841_), .B0(men_men_n839_), .Y(men_men_n844_));
  NA2        u0816(.A(men_men_n440_), .B(e), .Y(men_men_n845_));
  NO2        u0817(.A(men_men_n845_), .B(men_men_n508_), .Y(men_men_n846_));
  AOI210     u0818(.A0(men_men_n844_), .A1(men_men_n838_), .B0(men_men_n846_), .Y(men_men_n847_));
  NA3        u0819(.A(m), .B(l), .C(i), .Y(men_men_n848_));
  OAI220     u0820(.A0(men_men_n588_), .A1(men_men_n848_), .B0(men_men_n348_), .B1(men_men_n524_), .Y(men_men_n849_));
  NAi21      u0821(.An(men_men_n849_), .B(men_men_n435_), .Y(men_men_n850_));
  NA3        u0822(.A(men_men_n812_), .B(men_men_n566_), .C(men_men_n517_), .Y(men_men_n851_));
  OA210      u0823(.A0(men_men_n851_), .A1(men_men_n850_), .B0(men_men_n815_), .Y(men_men_n852_));
  INV        u0824(.A(men_men_n334_), .Y(men_men_n853_));
  NO2        u0825(.A(men_men_n128_), .B(men_men_n126_), .Y(men_men_n854_));
  NOi31      u0826(.An(k), .B(m), .C(l), .Y(men_men_n855_));
  NO2        u0827(.A(men_men_n335_), .B(men_men_n855_), .Y(men_men_n856_));
  AOI210     u0828(.A0(men_men_n856_), .A1(men_men_n854_), .B0(men_men_n594_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n797_), .B(men_men_n327_), .Y(men_men_n858_));
  NA2        u0830(.A(men_men_n337_), .B(men_men_n338_), .Y(men_men_n859_));
  OAI210     u0831(.A0(men_men_n205_), .A1(men_men_n212_), .B0(men_men_n859_), .Y(men_men_n860_));
  AOI220     u0832(.A0(men_men_n860_), .A1(men_men_n858_), .B0(men_men_n857_), .B1(men_men_n853_), .Y(men_men_n861_));
  NA2        u0833(.A(men_men_n172_), .B(men_men_n114_), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n862_), .B(men_men_n698_), .Y(men_men_n863_));
  NA3        u0835(.A(men_men_n863_), .B(men_men_n191_), .C(men_men_n31_), .Y(men_men_n864_));
  NA4        u0836(.A(men_men_n864_), .B(men_men_n861_), .C(men_men_n621_), .D(men_men_n80_), .Y(men_men_n865_));
  NO2        u0837(.A(men_men_n584_), .B(men_men_n494_), .Y(men_men_n866_));
  NOi21      u0838(.An(f), .B(d), .Y(men_men_n867_));
  NA2        u0839(.A(men_men_n867_), .B(m), .Y(men_men_n868_));
  NOi32      u0840(.An(g), .Bn(f), .C(d), .Y(men_men_n869_));
  NA4        u0841(.A(men_men_n869_), .B(men_men_n601_), .C(men_men_n29_), .D(m), .Y(men_men_n870_));
  NA2        u0842(.A(men_men_n303_), .B(men_men_n119_), .Y(men_men_n871_));
  AN2        u0843(.A(f), .B(d), .Y(men_men_n872_));
  NA3        u0844(.A(men_men_n473_), .B(men_men_n872_), .C(men_men_n82_), .Y(men_men_n873_));
  NO3        u0845(.A(men_men_n873_), .B(men_men_n71_), .C(men_men_n213_), .Y(men_men_n874_));
  NO2        u0846(.A(men_men_n281_), .B(men_men_n52_), .Y(men_men_n875_));
  NA2        u0847(.A(men_men_n871_), .B(men_men_n874_), .Y(men_men_n876_));
  NAi21      u0848(.An(men_men_n485_), .B(men_men_n876_), .Y(men_men_n877_));
  NO4        u0849(.A(men_men_n619_), .B(men_men_n133_), .C(men_men_n322_), .D(men_men_n155_), .Y(men_men_n878_));
  NO2        u0850(.A(men_men_n651_), .B(men_men_n322_), .Y(men_men_n879_));
  AN2        u0851(.A(men_men_n879_), .B(men_men_n679_), .Y(men_men_n880_));
  NO3        u0852(.A(men_men_n880_), .B(men_men_n878_), .C(men_men_n234_), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n599_), .B(men_men_n82_), .Y(men_men_n882_));
  NO2        u0854(.A(men_men_n859_), .B(men_men_n882_), .Y(men_men_n883_));
  NA3        u0855(.A(men_men_n163_), .B(men_men_n108_), .C(men_men_n107_), .Y(men_men_n884_));
  OAI220     u0856(.A0(men_men_n873_), .A1(men_men_n424_), .B0(men_men_n334_), .B1(men_men_n884_), .Y(men_men_n885_));
  NOi31      u0857(.An(men_men_n223_), .B(men_men_n885_), .C(men_men_n883_), .Y(men_men_n886_));
  NA2        u0858(.A(c), .B(men_men_n116_), .Y(men_men_n887_));
  NO2        u0859(.A(men_men_n887_), .B(men_men_n403_), .Y(men_men_n888_));
  NA3        u0860(.A(men_men_n888_), .B(men_men_n506_), .C(f), .Y(men_men_n889_));
  OR2        u0861(.A(men_men_n658_), .B(men_men_n538_), .Y(men_men_n890_));
  INV        u0862(.A(men_men_n890_), .Y(men_men_n891_));
  NA2        u0863(.A(men_men_n814_), .B(men_men_n111_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n892_), .B(men_men_n891_), .Y(men_men_n893_));
  NA4        u0865(.A(men_men_n893_), .B(men_men_n889_), .C(men_men_n886_), .D(men_men_n881_), .Y(men_men_n894_));
  NO4        u0866(.A(men_men_n894_), .B(men_men_n877_), .C(men_men_n865_), .D(men_men_n852_), .Y(men_men_n895_));
  OR2        u0867(.A(men_men_n873_), .B(men_men_n71_), .Y(men_men_n896_));
  NA2        u0868(.A(men_men_n840_), .B(g), .Y(men_men_n897_));
  AOI210     u0869(.A0(men_men_n897_), .A1(men_men_n285_), .B0(men_men_n896_), .Y(men_men_n898_));
  NO2        u0870(.A(men_men_n137_), .B(men_men_n133_), .Y(men_men_n899_));
  NO2        u0871(.A(men_men_n230_), .B(men_men_n224_), .Y(men_men_n900_));
  AOI220     u0872(.A0(men_men_n900_), .A1(men_men_n227_), .B0(men_men_n298_), .B1(men_men_n899_), .Y(men_men_n901_));
  NO2        u0873(.A(men_men_n424_), .B(men_men_n839_), .Y(men_men_n902_));
  NA2        u0874(.A(men_men_n902_), .B(men_men_n558_), .Y(men_men_n903_));
  NA2        u0875(.A(men_men_n903_), .B(men_men_n901_), .Y(men_men_n904_));
  NA2        u0876(.A(e), .B(d), .Y(men_men_n905_));
  OAI220     u0877(.A0(men_men_n905_), .A1(c), .B0(men_men_n317_), .B1(d), .Y(men_men_n906_));
  NA3        u0878(.A(men_men_n906_), .B(men_men_n452_), .C(men_men_n504_), .Y(men_men_n907_));
  AOI210     u0879(.A0(men_men_n512_), .A1(men_men_n184_), .B0(men_men_n230_), .Y(men_men_n908_));
  AOI210     u0880(.A0(men_men_n620_), .A1(men_men_n341_), .B0(men_men_n908_), .Y(men_men_n909_));
  NA3        u0881(.A(men_men_n171_), .B(men_men_n83_), .C(men_men_n34_), .Y(men_men_n910_));
  NA3        u0882(.A(men_men_n910_), .B(men_men_n909_), .C(men_men_n907_), .Y(men_men_n911_));
  NO3        u0883(.A(men_men_n911_), .B(men_men_n904_), .C(men_men_n898_), .Y(men_men_n912_));
  OR2        u0884(.A(men_men_n700_), .B(men_men_n216_), .Y(men_men_n913_));
  OAI220     u0885(.A0(men_men_n619_), .A1(men_men_n57_), .B0(men_men_n293_), .B1(j), .Y(men_men_n914_));
  AOI220     u0886(.A0(men_men_n914_), .A1(men_men_n879_), .B0(men_men_n609_), .B1(men_men_n618_), .Y(men_men_n915_));
  OAI210     u0887(.A0(men_men_n845_), .A1(men_men_n174_), .B0(men_men_n915_), .Y(men_men_n916_));
  AOI210     u0888(.A0(men_men_n118_), .A1(men_men_n117_), .B0(men_men_n259_), .Y(men_men_n917_));
  NO2        u0889(.A(men_men_n917_), .B(men_men_n870_), .Y(men_men_n918_));
  AO210      u0890(.A0(men_men_n858_), .A1(men_men_n849_), .B0(men_men_n918_), .Y(men_men_n919_));
  NO2        u0891(.A(men_men_n919_), .B(men_men_n916_), .Y(men_men_n920_));
  AO220      u0892(.A0(men_men_n452_), .A1(men_men_n748_), .B0(men_men_n179_), .B1(f), .Y(men_men_n921_));
  OAI210     u0893(.A0(men_men_n921_), .A1(men_men_n455_), .B0(men_men_n906_), .Y(men_men_n922_));
  NA2        u0894(.A(men_men_n851_), .B(men_men_n704_), .Y(men_men_n923_));
  AN4        u0895(.A(men_men_n923_), .B(men_men_n922_), .C(men_men_n920_), .D(men_men_n913_), .Y(men_men_n924_));
  NA4        u0896(.A(men_men_n924_), .B(men_men_n912_), .C(men_men_n895_), .D(men_men_n847_), .Y(men12));
  NO2        u0897(.A(men_men_n450_), .B(c), .Y(men_men_n926_));
  NO4        u0898(.A(men_men_n439_), .B(men_men_n252_), .C(men_men_n580_), .D(men_men_n213_), .Y(men_men_n927_));
  NA2        u0899(.A(men_men_n927_), .B(men_men_n926_), .Y(men_men_n928_));
  NO2        u0900(.A(men_men_n450_), .B(men_men_n116_), .Y(men_men_n929_));
  NO2        u0901(.A(men_men_n854_), .B(men_men_n348_), .Y(men_men_n930_));
  NO2        u0902(.A(men_men_n658_), .B(men_men_n374_), .Y(men_men_n931_));
  NA2        u0903(.A(men_men_n930_), .B(men_men_n929_), .Y(men_men_n932_));
  NA3        u0904(.A(men_men_n932_), .B(men_men_n928_), .C(men_men_n438_), .Y(men_men_n933_));
  AOI210     u0905(.A0(men_men_n233_), .A1(men_men_n333_), .B0(men_men_n202_), .Y(men_men_n934_));
  OR2        u0906(.A(men_men_n934_), .B(men_men_n927_), .Y(men_men_n935_));
  AOI210     u0907(.A0(men_men_n330_), .A1(men_men_n386_), .B0(men_men_n213_), .Y(men_men_n936_));
  OAI210     u0908(.A0(men_men_n936_), .A1(men_men_n935_), .B0(men_men_n398_), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n637_), .B(men_men_n262_), .Y(men_men_n938_));
  NO2        u0910(.A(men_men_n588_), .B(men_men_n848_), .Y(men_men_n939_));
  AOI220     u0911(.A0(men_men_n939_), .A1(men_men_n564_), .B0(men_men_n825_), .B1(men_men_n938_), .Y(men_men_n940_));
  NO2        u0912(.A(men_men_n154_), .B(men_men_n237_), .Y(men_men_n941_));
  NA3        u0913(.A(men_men_n941_), .B(men_men_n240_), .C(i), .Y(men_men_n942_));
  NA3        u0914(.A(men_men_n942_), .B(men_men_n940_), .C(men_men_n937_), .Y(men_men_n943_));
  OR2        u0915(.A(men_men_n318_), .B(men_men_n929_), .Y(men_men_n944_));
  NA2        u0916(.A(men_men_n944_), .B(men_men_n349_), .Y(men_men_n945_));
  NO3        u0917(.A(men_men_n133_), .B(men_men_n155_), .C(men_men_n213_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n946_), .B(men_men_n527_), .Y(men_men_n947_));
  NA4        u0919(.A(men_men_n440_), .B(men_men_n432_), .C(men_men_n185_), .D(g), .Y(men_men_n948_));
  NA3        u0920(.A(men_men_n948_), .B(men_men_n947_), .C(men_men_n945_), .Y(men_men_n949_));
  NO3        u0921(.A(men_men_n949_), .B(men_men_n943_), .C(men_men_n933_), .Y(men_men_n950_));
  NO2        u0922(.A(men_men_n365_), .B(men_men_n364_), .Y(men_men_n951_));
  INV        u0923(.A(men_men_n585_), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n551_), .B(men_men_n147_), .Y(men_men_n953_));
  NOi21      u0925(.An(men_men_n34_), .B(men_men_n651_), .Y(men_men_n954_));
  AOI220     u0926(.A0(men_men_n954_), .A1(men_men_n953_), .B0(men_men_n952_), .B1(men_men_n951_), .Y(men_men_n955_));
  OAI210     u0927(.A0(men_men_n250_), .A1(men_men_n43_), .B0(men_men_n955_), .Y(men_men_n956_));
  NA2        u0928(.A(men_men_n430_), .B(men_men_n264_), .Y(men_men_n957_));
  NO3        u0929(.A(men_men_n827_), .B(men_men_n87_), .C(men_men_n403_), .Y(men_men_n958_));
  NAi31      u0930(.An(men_men_n958_), .B(men_men_n957_), .C(men_men_n314_), .Y(men_men_n959_));
  NO2        u0931(.A(men_men_n47_), .B(men_men_n43_), .Y(men_men_n960_));
  NO2        u0932(.A(men_men_n501_), .B(men_men_n293_), .Y(men_men_n961_));
  INV        u0933(.A(men_men_n961_), .Y(men_men_n962_));
  NO2        u0934(.A(men_men_n962_), .B(men_men_n147_), .Y(men_men_n963_));
  NA2        u0935(.A(men_men_n630_), .B(men_men_n358_), .Y(men_men_n964_));
  OAI210     u0936(.A0(men_men_n734_), .A1(men_men_n964_), .B0(men_men_n362_), .Y(men_men_n965_));
  NO4        u0937(.A(men_men_n965_), .B(men_men_n963_), .C(men_men_n959_), .D(men_men_n956_), .Y(men_men_n966_));
  NA2        u0938(.A(men_men_n341_), .B(g), .Y(men_men_n967_));
  NA2        u0939(.A(men_men_n166_), .B(i), .Y(men_men_n968_));
  NA2        u0940(.A(men_men_n414_), .B(men_men_n37_), .Y(men_men_n969_));
  NO2        u0941(.A(men_men_n147_), .B(men_men_n82_), .Y(men_men_n970_));
  OR2        u0942(.A(men_men_n970_), .B(men_men_n550_), .Y(men_men_n971_));
  NA2        u0943(.A(men_men_n551_), .B(men_men_n378_), .Y(men_men_n972_));
  AOI210     u0944(.A0(men_men_n972_), .A1(n), .B0(men_men_n971_), .Y(men_men_n973_));
  OAI220     u0945(.A0(men_men_n973_), .A1(men_men_n967_), .B0(men_men_n969_), .B1(men_men_n327_), .Y(men_men_n974_));
  NO2        u0946(.A(men_men_n658_), .B(men_men_n494_), .Y(men_men_n975_));
  NA3        u0947(.A(men_men_n337_), .B(men_men_n625_), .C(i), .Y(men_men_n976_));
  OAI210     u0948(.A0(men_men_n434_), .A1(men_men_n303_), .B0(men_men_n976_), .Y(men_men_n977_));
  OAI220     u0949(.A0(men_men_n977_), .A1(men_men_n975_), .B0(men_men_n675_), .B1(men_men_n760_), .Y(men_men_n978_));
  NA2        u0950(.A(men_men_n603_), .B(men_men_n113_), .Y(men_men_n979_));
  OR3        u0951(.A(men_men_n303_), .B(men_men_n429_), .C(f), .Y(men_men_n980_));
  NA3        u0952(.A(men_men_n625_), .B(men_men_n78_), .C(i), .Y(men_men_n981_));
  OA220      u0953(.A0(men_men_n981_), .A1(men_men_n979_), .B0(men_men_n980_), .B1(men_men_n587_), .Y(men_men_n982_));
  NA3        u0954(.A(men_men_n319_), .B(men_men_n118_), .C(g), .Y(men_men_n983_));
  AOI210     u0955(.A0(men_men_n672_), .A1(men_men_n983_), .B0(m), .Y(men_men_n984_));
  OAI210     u0956(.A0(men_men_n984_), .A1(men_men_n930_), .B0(men_men_n318_), .Y(men_men_n985_));
  NA2        u0957(.A(men_men_n691_), .B(men_men_n882_), .Y(men_men_n986_));
  INV        u0958(.A(men_men_n435_), .Y(men_men_n987_));
  NA2        u0959(.A(men_men_n221_), .B(men_men_n75_), .Y(men_men_n988_));
  NA3        u0960(.A(men_men_n988_), .B(men_men_n981_), .C(men_men_n980_), .Y(men_men_n989_));
  AOI220     u0961(.A0(men_men_n989_), .A1(men_men_n258_), .B0(men_men_n987_), .B1(men_men_n986_), .Y(men_men_n990_));
  NA4        u0962(.A(men_men_n990_), .B(men_men_n985_), .C(men_men_n982_), .D(men_men_n978_), .Y(men_men_n991_));
  NA2        u0963(.A(men_men_n660_), .B(men_men_n86_), .Y(men_men_n992_));
  NO2        u0964(.A(men_men_n458_), .B(men_men_n213_), .Y(men_men_n993_));
  AOI220     u0965(.A0(men_men_n993_), .A1(men_men_n379_), .B0(men_men_n944_), .B1(men_men_n217_), .Y(men_men_n994_));
  AOI220     u0966(.A0(men_men_n931_), .A1(men_men_n941_), .B0(men_men_n586_), .B1(men_men_n88_), .Y(men_men_n995_));
  NA3        u0967(.A(men_men_n995_), .B(men_men_n994_), .C(men_men_n992_), .Y(men_men_n996_));
  OAI210     u0968(.A0(men_men_n987_), .A1(men_men_n939_), .B0(men_men_n540_), .Y(men_men_n997_));
  AOI210     u0969(.A0(men_men_n415_), .A1(men_men_n407_), .B0(men_men_n827_), .Y(men_men_n998_));
  OAI210     u0970(.A0(men_men_n365_), .A1(men_men_n364_), .B0(men_men_n109_), .Y(men_men_n999_));
  AOI210     u0971(.A0(men_men_n999_), .A1(men_men_n532_), .B0(men_men_n998_), .Y(men_men_n1000_));
  NA2        u0972(.A(men_men_n984_), .B(men_men_n929_), .Y(men_men_n1001_));
  NA2        u0973(.A(men_men_n642_), .B(men_men_n527_), .Y(men_men_n1002_));
  NA4        u0974(.A(men_men_n1002_), .B(men_men_n1001_), .C(men_men_n1000_), .D(men_men_n997_), .Y(men_men_n1003_));
  NO4        u0975(.A(men_men_n1003_), .B(men_men_n996_), .C(men_men_n991_), .D(men_men_n974_), .Y(men_men_n1004_));
  NAi31      u0976(.An(men_men_n143_), .B(men_men_n416_), .C(n), .Y(men_men_n1005_));
  NO3        u0977(.A(men_men_n126_), .B(men_men_n335_), .C(men_men_n855_), .Y(men_men_n1006_));
  NO2        u0978(.A(men_men_n1006_), .B(men_men_n1005_), .Y(men_men_n1007_));
  NA2        u0979(.A(men_men_n230_), .B(men_men_n175_), .Y(men_men_n1008_));
  NO3        u0980(.A(men_men_n301_), .B(men_men_n440_), .C(men_men_n179_), .Y(men_men_n1009_));
  NOi31      u0981(.An(men_men_n1008_), .B(men_men_n1009_), .C(men_men_n213_), .Y(men_men_n1010_));
  NAi21      u0982(.An(men_men_n551_), .B(men_men_n993_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n433_), .B(men_men_n882_), .Y(men_men_n1012_));
  NO3        u0984(.A(men_men_n434_), .B(men_men_n303_), .C(men_men_n71_), .Y(men_men_n1013_));
  AOI220     u0985(.A0(men_men_n1013_), .A1(men_men_n1012_), .B0(men_men_n477_), .B1(g), .Y(men_men_n1014_));
  NA2        u0986(.A(men_men_n1014_), .B(men_men_n1011_), .Y(men_men_n1015_));
  OAI220     u0987(.A0(men_men_n1005_), .A1(men_men_n233_), .B0(men_men_n976_), .B1(men_men_n600_), .Y(men_men_n1016_));
  NA2        u0988(.A(men_men_n934_), .B(men_men_n926_), .Y(men_men_n1017_));
  NO3        u0989(.A(men_men_n541_), .B(men_men_n152_), .C(men_men_n212_), .Y(men_men_n1018_));
  OAI210     u0990(.A0(men_men_n1018_), .A1(men_men_n522_), .B0(men_men_n375_), .Y(men_men_n1019_));
  OAI210     u0991(.A0(men_men_n931_), .A1(men_men_n939_), .B0(men_men_n423_), .Y(men_men_n1020_));
  NA4        u0992(.A(men_men_n1020_), .B(men_men_n1019_), .C(men_men_n1017_), .D(men_men_n617_), .Y(men_men_n1021_));
  OAI210     u0993(.A0(men_men_n934_), .A1(men_men_n927_), .B0(men_men_n1008_), .Y(men_men_n1022_));
  NA3        u0994(.A(men_men_n972_), .B(men_men_n482_), .C(men_men_n44_), .Y(men_men_n1023_));
  AOI210     u0995(.A0(men_men_n377_), .A1(men_men_n375_), .B0(men_men_n326_), .Y(men_men_n1024_));
  NA4        u0996(.A(men_men_n1024_), .B(men_men_n1023_), .C(men_men_n1022_), .D(men_men_n273_), .Y(men_men_n1025_));
  OR3        u0997(.A(men_men_n1025_), .B(men_men_n1021_), .C(men_men_n1016_), .Y(men_men_n1026_));
  NO4        u0998(.A(men_men_n1026_), .B(men_men_n1015_), .C(men_men_n1010_), .D(men_men_n1007_), .Y(men_men_n1027_));
  NA4        u0999(.A(men_men_n1027_), .B(men_men_n1004_), .C(men_men_n966_), .D(men_men_n950_), .Y(men13));
  AN2        u1000(.A(c), .B(b), .Y(men_men_n1029_));
  NA3        u1001(.A(men_men_n249_), .B(men_men_n1029_), .C(m), .Y(men_men_n1030_));
  NA2        u1002(.A(men_men_n492_), .B(f), .Y(men_men_n1031_));
  NO4        u1003(.A(men_men_n1031_), .B(men_men_n1030_), .C(j), .D(men_men_n581_), .Y(men_men_n1032_));
  NA2        u1004(.A(men_men_n264_), .B(men_men_n1029_), .Y(men_men_n1033_));
  NO4        u1005(.A(men_men_n1033_), .B(men_men_n1031_), .C(men_men_n968_), .D(a), .Y(men_men_n1034_));
  NAi32      u1006(.An(d), .Bn(c), .C(e), .Y(men_men_n1035_));
  NA2        u1007(.A(men_men_n142_), .B(men_men_n43_), .Y(men_men_n1036_));
  NO4        u1008(.A(men_men_n1036_), .B(men_men_n1035_), .C(men_men_n588_), .D(men_men_n300_), .Y(men_men_n1037_));
  NA2        u1009(.A(men_men_n664_), .B(men_men_n224_), .Y(men_men_n1038_));
  NA2        u1010(.A(men_men_n406_), .B(men_men_n212_), .Y(men_men_n1039_));
  AN2        u1011(.A(d), .B(c), .Y(men_men_n1040_));
  NA2        u1012(.A(men_men_n1040_), .B(men_men_n116_), .Y(men_men_n1041_));
  NO4        u1013(.A(men_men_n1041_), .B(men_men_n1039_), .C(men_men_n180_), .D(men_men_n172_), .Y(men_men_n1042_));
  NA2        u1014(.A(men_men_n492_), .B(c), .Y(men_men_n1043_));
  NO4        u1015(.A(men_men_n1036_), .B(men_men_n584_), .C(men_men_n1043_), .D(men_men_n300_), .Y(men_men_n1044_));
  AO210      u1016(.A0(men_men_n1042_), .A1(men_men_n1038_), .B0(men_men_n1044_), .Y(men_men_n1045_));
  OR4        u1017(.A(men_men_n1045_), .B(men_men_n1037_), .C(men_men_n1034_), .D(men_men_n1032_), .Y(men_men_n1046_));
  NAi32      u1018(.An(f), .Bn(e), .C(c), .Y(men_men_n1047_));
  NO2        u1019(.A(men_men_n1047_), .B(men_men_n149_), .Y(men_men_n1048_));
  NA2        u1020(.A(men_men_n1048_), .B(g), .Y(men_men_n1049_));
  OR3        u1021(.A(men_men_n224_), .B(men_men_n180_), .C(men_men_n172_), .Y(men_men_n1050_));
  NO2        u1022(.A(men_men_n1050_), .B(men_men_n1049_), .Y(men_men_n1051_));
  NO2        u1023(.A(men_men_n1043_), .B(men_men_n300_), .Y(men_men_n1052_));
  NO2        u1024(.A(j), .B(men_men_n43_), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n627_), .B(men_men_n1053_), .Y(men_men_n1054_));
  NOi21      u1026(.An(men_men_n1052_), .B(men_men_n1054_), .Y(men_men_n1055_));
  NO2        u1027(.A(men_men_n764_), .B(men_men_n112_), .Y(men_men_n1056_));
  NOi41      u1028(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1057_));
  NA2        u1029(.A(men_men_n1057_), .B(men_men_n1056_), .Y(men_men_n1058_));
  NO2        u1030(.A(men_men_n1058_), .B(men_men_n1049_), .Y(men_men_n1059_));
  OR3        u1031(.A(e), .B(d), .C(c), .Y(men_men_n1060_));
  NA3        u1032(.A(k), .B(j), .C(i), .Y(men_men_n1061_));
  NO3        u1033(.A(men_men_n1061_), .B(men_men_n300_), .C(men_men_n89_), .Y(men_men_n1062_));
  NOi21      u1034(.An(men_men_n1062_), .B(men_men_n1060_), .Y(men_men_n1063_));
  OR4        u1035(.A(men_men_n1063_), .B(men_men_n1059_), .C(men_men_n1055_), .D(men_men_n1051_), .Y(men_men_n1064_));
  NA3        u1036(.A(men_men_n465_), .B(men_men_n329_), .C(men_men_n52_), .Y(men_men_n1065_));
  NO2        u1037(.A(men_men_n1065_), .B(men_men_n1054_), .Y(men_men_n1066_));
  NO4        u1038(.A(men_men_n1065_), .B(men_men_n584_), .C(men_men_n447_), .D(men_men_n43_), .Y(men_men_n1067_));
  NO2        u1039(.A(f), .B(c), .Y(men_men_n1068_));
  NOi21      u1040(.An(men_men_n1068_), .B(men_men_n439_), .Y(men_men_n1069_));
  NA2        u1041(.A(men_men_n1069_), .B(men_men_n55_), .Y(men_men_n1070_));
  OR2        u1042(.A(k), .B(i), .Y(men_men_n1071_));
  NO3        u1043(.A(men_men_n1071_), .B(men_men_n244_), .C(l), .Y(men_men_n1072_));
  NOi31      u1044(.An(men_men_n1072_), .B(men_men_n1070_), .C(j), .Y(men_men_n1073_));
  OR3        u1045(.A(men_men_n1073_), .B(men_men_n1067_), .C(men_men_n1066_), .Y(men_men_n1074_));
  OR3        u1046(.A(men_men_n1074_), .B(men_men_n1064_), .C(men_men_n1046_), .Y(men02));
  OR2        u1047(.A(l), .B(k), .Y(men_men_n1076_));
  OR3        u1048(.A(h), .B(g), .C(f), .Y(men_men_n1077_));
  OR3        u1049(.A(n), .B(m), .C(i), .Y(men_men_n1078_));
  NO4        u1050(.A(men_men_n1078_), .B(men_men_n1077_), .C(men_men_n1076_), .D(men_men_n1060_), .Y(men_men_n1079_));
  NOi31      u1051(.An(e), .B(d), .C(c), .Y(men_men_n1080_));
  AOI210     u1052(.A0(men_men_n1062_), .A1(men_men_n1080_), .B0(men_men_n1037_), .Y(men_men_n1081_));
  AN3        u1053(.A(g), .B(f), .C(c), .Y(men_men_n1082_));
  NA3        u1054(.A(men_men_n1082_), .B(men_men_n465_), .C(h), .Y(men_men_n1083_));
  OR2        u1055(.A(men_men_n1061_), .B(men_men_n300_), .Y(men_men_n1084_));
  OR2        u1056(.A(men_men_n1084_), .B(men_men_n1083_), .Y(men_men_n1085_));
  NO3        u1057(.A(men_men_n1065_), .B(men_men_n1036_), .C(men_men_n584_), .Y(men_men_n1086_));
  NO2        u1058(.A(men_men_n1086_), .B(men_men_n1051_), .Y(men_men_n1087_));
  NA3        u1059(.A(l), .B(k), .C(j), .Y(men_men_n1088_));
  NA2        u1060(.A(i), .B(h), .Y(men_men_n1089_));
  NO3        u1061(.A(men_men_n1089_), .B(men_men_n1088_), .C(men_men_n133_), .Y(men_men_n1090_));
  NO3        u1062(.A(men_men_n144_), .B(men_men_n280_), .C(men_men_n213_), .Y(men_men_n1091_));
  AOI210     u1063(.A0(men_men_n1091_), .A1(men_men_n1090_), .B0(men_men_n1055_), .Y(men_men_n1092_));
  NA3        u1064(.A(c), .B(b), .C(a), .Y(men_men_n1093_));
  NO3        u1065(.A(men_men_n1093_), .B(men_men_n905_), .C(men_men_n212_), .Y(men_men_n1094_));
  NO3        u1066(.A(men_men_n1061_), .B(men_men_n47_), .C(men_men_n112_), .Y(men_men_n1095_));
  AOI210     u1067(.A0(men_men_n1095_), .A1(men_men_n1094_), .B0(men_men_n1066_), .Y(men_men_n1096_));
  AN4        u1068(.A(men_men_n1096_), .B(men_men_n1092_), .C(men_men_n1087_), .D(men_men_n1085_), .Y(men_men_n1097_));
  NO2        u1069(.A(men_men_n1041_), .B(men_men_n1039_), .Y(men_men_n1098_));
  NA2        u1070(.A(men_men_n1058_), .B(men_men_n1050_), .Y(men_men_n1099_));
  AOI210     u1071(.A0(men_men_n1099_), .A1(men_men_n1098_), .B0(men_men_n1032_), .Y(men_men_n1100_));
  NAi41      u1072(.An(men_men_n1079_), .B(men_men_n1100_), .C(men_men_n1097_), .D(men_men_n1081_), .Y(men03));
  NO2        u1073(.A(men_men_n524_), .B(men_men_n594_), .Y(men_men_n1102_));
  NA4        u1074(.A(men_men_n86_), .B(men_men_n85_), .C(g), .D(men_men_n212_), .Y(men_men_n1103_));
  NA4        u1075(.A(men_men_n574_), .B(m), .C(men_men_n112_), .D(men_men_n212_), .Y(men_men_n1104_));
  NA2        u1076(.A(men_men_n1104_), .B(men_men_n1103_), .Y(men_men_n1105_));
  NO3        u1077(.A(men_men_n1105_), .B(men_men_n1102_), .C(men_men_n999_), .Y(men_men_n1106_));
  NOi41      u1078(.An(men_men_n812_), .B(men_men_n860_), .C(men_men_n850_), .D(men_men_n714_), .Y(men_men_n1107_));
  OAI220     u1079(.A0(men_men_n1107_), .A1(men_men_n691_), .B0(men_men_n1106_), .B1(men_men_n585_), .Y(men_men_n1108_));
  NOi31      u1080(.An(i), .B(k), .C(j), .Y(men_men_n1109_));
  NA4        u1081(.A(men_men_n1109_), .B(men_men_n1080_), .C(men_men_n337_), .D(men_men_n329_), .Y(men_men_n1110_));
  OAI210     u1082(.A0(men_men_n827_), .A1(men_men_n417_), .B0(men_men_n1110_), .Y(men_men_n1111_));
  NOi31      u1083(.An(m), .B(n), .C(f), .Y(men_men_n1112_));
  NA2        u1084(.A(men_men_n1112_), .B(men_men_n49_), .Y(men_men_n1113_));
  AN2        u1085(.A(e), .B(c), .Y(men_men_n1114_));
  NA2        u1086(.A(men_men_n1114_), .B(a), .Y(men_men_n1115_));
  OAI220     u1087(.A0(men_men_n1115_), .A1(men_men_n1113_), .B0(men_men_n890_), .B1(men_men_n422_), .Y(men_men_n1116_));
  NA2        u1088(.A(men_men_n504_), .B(l), .Y(men_men_n1117_));
  NOi31      u1089(.An(men_men_n869_), .B(men_men_n1030_), .C(men_men_n1117_), .Y(men_men_n1118_));
  NO4        u1090(.A(men_men_n1118_), .B(men_men_n1116_), .C(men_men_n1111_), .D(men_men_n998_), .Y(men_men_n1119_));
  NO2        u1091(.A(men_men_n280_), .B(a), .Y(men_men_n1120_));
  INV        u1092(.A(men_men_n1037_), .Y(men_men_n1121_));
  NO2        u1093(.A(men_men_n1089_), .B(men_men_n480_), .Y(men_men_n1122_));
  NO2        u1094(.A(men_men_n85_), .B(g), .Y(men_men_n1123_));
  AOI210     u1095(.A0(men_men_n1123_), .A1(men_men_n1122_), .B0(men_men_n1072_), .Y(men_men_n1124_));
  OR2        u1096(.A(men_men_n1124_), .B(men_men_n1070_), .Y(men_men_n1125_));
  NA3        u1097(.A(men_men_n1125_), .B(men_men_n1121_), .C(men_men_n1119_), .Y(men_men_n1126_));
  NO4        u1098(.A(men_men_n1126_), .B(men_men_n1108_), .C(men_men_n829_), .D(men_men_n563_), .Y(men_men_n1127_));
  NA2        u1099(.A(c), .B(b), .Y(men_men_n1128_));
  NO2        u1100(.A(men_men_n703_), .B(men_men_n1128_), .Y(men_men_n1129_));
  OAI210     u1101(.A0(men_men_n868_), .A1(men_men_n843_), .B0(men_men_n410_), .Y(men_men_n1130_));
  NA2        u1102(.A(men_men_n1130_), .B(men_men_n1129_), .Y(men_men_n1131_));
  NAi21      u1103(.An(men_men_n418_), .B(men_men_n1129_), .Y(men_men_n1132_));
  OAI210     u1104(.A0(men_men_n545_), .A1(men_men_n39_), .B0(men_men_n1120_), .Y(men_men_n1133_));
  NA2        u1105(.A(men_men_n1133_), .B(men_men_n1132_), .Y(men_men_n1134_));
  INV        u1106(.A(men_men_n119_), .Y(men_men_n1135_));
  NA2        u1107(.A(men_men_n1135_), .B(g), .Y(men_men_n1136_));
  NAi21      u1108(.An(f), .B(d), .Y(men_men_n1137_));
  NO2        u1109(.A(men_men_n1137_), .B(men_men_n1093_), .Y(men_men_n1138_));
  INV        u1110(.A(men_men_n1138_), .Y(men_men_n1139_));
  AOI210     u1111(.A0(men_men_n1136_), .A1(men_men_n285_), .B0(men_men_n1139_), .Y(men_men_n1140_));
  AOI210     u1112(.A0(men_men_n1140_), .A1(men_men_n113_), .B0(men_men_n1134_), .Y(men_men_n1141_));
  NO2        u1113(.A(men_men_n186_), .B(men_men_n237_), .Y(men_men_n1142_));
  NA2        u1114(.A(men_men_n1142_), .B(m), .Y(men_men_n1143_));
  NA3        u1115(.A(men_men_n917_), .B(men_men_n1117_), .C(men_men_n168_), .Y(men_men_n1144_));
  NA2        u1116(.A(men_men_n1144_), .B(men_men_n469_), .Y(men_men_n1145_));
  NO2        u1117(.A(men_men_n1145_), .B(men_men_n1143_), .Y(men_men_n1146_));
  NA2        u1118(.A(men_men_n558_), .B(men_men_n405_), .Y(men_men_n1147_));
  NA2        u1119(.A(men_men_n162_), .B(men_men_n33_), .Y(men_men_n1148_));
  AOI210     u1120(.A0(men_men_n964_), .A1(men_men_n1148_), .B0(men_men_n213_), .Y(men_men_n1149_));
  NA2        u1121(.A(men_men_n1149_), .B(men_men_n1138_), .Y(men_men_n1150_));
  NO2        u1122(.A(men_men_n368_), .B(men_men_n367_), .Y(men_men_n1151_));
  INV        u1123(.A(men_men_n958_), .Y(men_men_n1152_));
  NAi41      u1124(.An(men_men_n1151_), .B(men_men_n1152_), .C(men_men_n1150_), .D(men_men_n1147_), .Y(men_men_n1153_));
  NO2        u1125(.A(men_men_n1153_), .B(men_men_n1146_), .Y(men_men_n1154_));
  NA4        u1126(.A(men_men_n1154_), .B(men_men_n1141_), .C(men_men_n1131_), .D(men_men_n1127_), .Y(men00));
  AOI210     u1127(.A0(men_men_n902_), .A1(men_men_n941_), .B0(men_men_n1111_), .Y(men_men_n1156_));
  NO3        u1128(.A(men_men_n1086_), .B(men_men_n958_), .C(men_men_n711_), .Y(men_men_n1157_));
  NA3        u1129(.A(men_men_n1157_), .B(men_men_n1156_), .C(men_men_n1000_), .Y(men_men_n1158_));
  NA2        u1130(.A(men_men_n506_), .B(f), .Y(men_men_n1159_));
  OAI210     u1131(.A0(men_men_n1006_), .A1(men_men_n40_), .B0(men_men_n644_), .Y(men_men_n1160_));
  NA3        u1132(.A(men_men_n1160_), .B(men_men_n257_), .C(n), .Y(men_men_n1161_));
  AOI210     u1133(.A0(men_men_n1161_), .A1(men_men_n1159_), .B0(men_men_n1041_), .Y(men_men_n1162_));
  NO3        u1134(.A(men_men_n1162_), .B(men_men_n1158_), .C(men_men_n1064_), .Y(men_men_n1163_));
  NA3        u1135(.A(men_men_n171_), .B(men_men_n44_), .C(men_men_n43_), .Y(men_men_n1164_));
  NA3        u1136(.A(d), .B(men_men_n52_), .C(b), .Y(men_men_n1165_));
  NOi31      u1137(.An(n), .B(m), .C(i), .Y(men_men_n1166_));
  NA3        u1138(.A(men_men_n1166_), .B(men_men_n647_), .C(men_men_n49_), .Y(men_men_n1167_));
  OAI210     u1139(.A0(men_men_n1165_), .A1(men_men_n1164_), .B0(men_men_n1167_), .Y(men_men_n1168_));
  NO2        u1140(.A(men_men_n1168_), .B(men_men_n1151_), .Y(men_men_n1169_));
  NO4        u1141(.A(men_men_n483_), .B(men_men_n351_), .C(men_men_n1128_), .D(men_men_n55_), .Y(men_men_n1170_));
  OR2        u1142(.A(men_men_n381_), .B(men_men_n136_), .Y(men_men_n1171_));
  NO2        u1143(.A(h), .B(g), .Y(men_men_n1172_));
  NA4        u1144(.A(men_men_n495_), .B(men_men_n465_), .C(men_men_n1172_), .D(men_men_n1029_), .Y(men_men_n1173_));
  OAI220     u1145(.A0(men_men_n524_), .A1(men_men_n594_), .B0(men_men_n90_), .B1(men_men_n89_), .Y(men_men_n1174_));
  AOI220     u1146(.A0(men_men_n1174_), .A1(men_men_n532_), .B0(men_men_n946_), .B1(men_men_n575_), .Y(men_men_n1175_));
  AOI220     u1147(.A0(men_men_n311_), .A1(men_men_n246_), .B0(men_men_n181_), .B1(men_men_n151_), .Y(men_men_n1176_));
  NA4        u1148(.A(men_men_n1176_), .B(men_men_n1175_), .C(men_men_n1173_), .D(men_men_n1171_), .Y(men_men_n1177_));
  NO3        u1149(.A(men_men_n1177_), .B(men_men_n1170_), .C(men_men_n266_), .Y(men_men_n1178_));
  INV        u1150(.A(men_men_n316_), .Y(men_men_n1179_));
  AOI210     u1151(.A0(men_men_n246_), .A1(men_men_n341_), .B0(men_men_n577_), .Y(men_men_n1180_));
  NA3        u1152(.A(men_men_n1180_), .B(men_men_n1179_), .C(men_men_n157_), .Y(men_men_n1181_));
  NO2        u1153(.A(men_men_n239_), .B(men_men_n185_), .Y(men_men_n1182_));
  NA2        u1154(.A(men_men_n1182_), .B(men_men_n423_), .Y(men_men_n1183_));
  NA3        u1155(.A(men_men_n183_), .B(men_men_n112_), .C(g), .Y(men_men_n1184_));
  NA3        u1156(.A(men_men_n465_), .B(men_men_n40_), .C(f), .Y(men_men_n1185_));
  NOi31      u1157(.An(men_men_n875_), .B(men_men_n1185_), .C(men_men_n1184_), .Y(men_men_n1186_));
  NAi31      u1158(.An(men_men_n188_), .B(men_men_n866_), .C(men_men_n465_), .Y(men_men_n1187_));
  NAi31      u1159(.An(men_men_n1186_), .B(men_men_n1187_), .C(men_men_n1183_), .Y(men_men_n1188_));
  NO2        u1160(.A(men_men_n274_), .B(men_men_n71_), .Y(men_men_n1189_));
  NO3        u1161(.A(men_men_n422_), .B(men_men_n839_), .C(n), .Y(men_men_n1190_));
  AOI210     u1162(.A0(men_men_n1190_), .A1(men_men_n1189_), .B0(men_men_n1079_), .Y(men_men_n1191_));
  NAi31      u1163(.An(men_men_n1044_), .B(men_men_n1191_), .C(men_men_n70_), .Y(men_men_n1192_));
  NO4        u1164(.A(men_men_n1192_), .B(men_men_n1188_), .C(men_men_n1181_), .D(men_men_n516_), .Y(men_men_n1193_));
  AN3        u1165(.A(men_men_n1193_), .B(men_men_n1178_), .C(men_men_n1169_), .Y(men_men_n1194_));
  NA2        u1166(.A(men_men_n532_), .B(men_men_n100_), .Y(men_men_n1195_));
  NA3        u1167(.A(men_men_n1112_), .B(men_men_n603_), .C(men_men_n464_), .Y(men_men_n1196_));
  NA4        u1168(.A(men_men_n1196_), .B(men_men_n559_), .C(men_men_n1195_), .D(men_men_n242_), .Y(men_men_n1197_));
  NA2        u1169(.A(men_men_n1105_), .B(men_men_n532_), .Y(men_men_n1198_));
  NA2        u1170(.A(men_men_n1198_), .B(men_men_n289_), .Y(men_men_n1199_));
  OAI210     u1171(.A0(men_men_n463_), .A1(men_men_n120_), .B0(men_men_n870_), .Y(men_men_n1200_));
  AOI220     u1172(.A0(men_men_n1200_), .A1(men_men_n1144_), .B0(men_men_n558_), .B1(men_men_n405_), .Y(men_men_n1201_));
  OR4        u1173(.A(men_men_n1041_), .B(men_men_n272_), .C(men_men_n222_), .D(e), .Y(men_men_n1202_));
  NA2        u1174(.A(n), .B(e), .Y(men_men_n1203_));
  NO2        u1175(.A(men_men_n1203_), .B(men_men_n149_), .Y(men_men_n1204_));
  OAI210     u1176(.A0(men_men_n352_), .A1(men_men_n305_), .B0(men_men_n445_), .Y(men_men_n1205_));
  NA3        u1177(.A(men_men_n1205_), .B(men_men_n1202_), .C(men_men_n1201_), .Y(men_men_n1206_));
  AOI210     u1178(.A0(men_men_n1204_), .A1(men_men_n857_), .B0(men_men_n828_), .Y(men_men_n1207_));
  NA2        u1179(.A(men_men_n954_), .B(men_men_n575_), .Y(men_men_n1208_));
  NO2        u1180(.A(men_men_n64_), .B(h), .Y(men_men_n1209_));
  NO3        u1181(.A(men_men_n1041_), .B(men_men_n1039_), .C(men_men_n727_), .Y(men_men_n1210_));
  INV        u1182(.A(men_men_n133_), .Y(men_men_n1211_));
  AN2        u1183(.A(men_men_n1211_), .B(men_men_n1091_), .Y(men_men_n1212_));
  OAI210     u1184(.A0(men_men_n1212_), .A1(men_men_n1210_), .B0(men_men_n1209_), .Y(men_men_n1213_));
  NA3        u1185(.A(men_men_n1213_), .B(men_men_n1208_), .C(men_men_n1207_), .Y(men_men_n1214_));
  NO4        u1186(.A(men_men_n1214_), .B(men_men_n1206_), .C(men_men_n1199_), .D(men_men_n1197_), .Y(men_men_n1215_));
  NA2        u1187(.A(men_men_n844_), .B(men_men_n759_), .Y(men_men_n1216_));
  NA4        u1188(.A(men_men_n1216_), .B(men_men_n1215_), .C(men_men_n1194_), .D(men_men_n1163_), .Y(men01));
  AN2        u1189(.A(men_men_n1019_), .B(men_men_n1017_), .Y(men_men_n1218_));
  NO3        u1190(.A(men_men_n808_), .B(men_men_n800_), .C(men_men_n278_), .Y(men_men_n1219_));
  NA2        u1191(.A(men_men_n391_), .B(i), .Y(men_men_n1220_));
  NA3        u1192(.A(men_men_n1220_), .B(men_men_n1219_), .C(men_men_n1218_), .Y(men_men_n1221_));
  NA2        u1193(.A(men_men_n586_), .B(men_men_n88_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n551_), .B(men_men_n271_), .Y(men_men_n1223_));
  NA2        u1195(.A(men_men_n961_), .B(men_men_n1223_), .Y(men_men_n1224_));
  NA4        u1196(.A(men_men_n1224_), .B(men_men_n1222_), .C(men_men_n915_), .D(men_men_n328_), .Y(men_men_n1225_));
  NA2        u1197(.A(men_men_n43_), .B(f), .Y(men_men_n1226_));
  NA2        u1198(.A(men_men_n709_), .B(men_men_n95_), .Y(men_men_n1227_));
  NO2        u1199(.A(men_men_n1227_), .B(men_men_n1226_), .Y(men_men_n1228_));
  NO2        u1200(.A(men_men_n786_), .B(men_men_n600_), .Y(men_men_n1229_));
  AOI210     u1201(.A0(men_men_n1228_), .A1(men_men_n632_), .B0(men_men_n1229_), .Y(men_men_n1230_));
  INV        u1202(.A(men_men_n118_), .Y(men_men_n1231_));
  OR2        u1203(.A(men_men_n1231_), .B(men_men_n583_), .Y(men_men_n1232_));
  NAi41      u1204(.An(men_men_n165_), .B(men_men_n1232_), .C(men_men_n1230_), .D(men_men_n901_), .Y(men_men_n1233_));
  NO3        u1205(.A(men_men_n787_), .B(men_men_n674_), .C(men_men_n509_), .Y(men_men_n1234_));
  NA4        u1206(.A(men_men_n709_), .B(men_men_n95_), .C(men_men_n43_), .D(men_men_n212_), .Y(men_men_n1235_));
  OA220      u1207(.A0(men_men_n1235_), .A1(men_men_n667_), .B0(men_men_n196_), .B1(men_men_n194_), .Y(men_men_n1236_));
  NA3        u1208(.A(men_men_n1236_), .B(men_men_n1234_), .C(men_men_n139_), .Y(men_men_n1237_));
  NO4        u1209(.A(men_men_n1237_), .B(men_men_n1233_), .C(men_men_n1225_), .D(men_men_n1221_), .Y(men_men_n1238_));
  NA2        u1210(.A(men_men_n295_), .B(men_men_n527_), .Y(men_men_n1239_));
  NA2        u1211(.A(men_men_n535_), .B(men_men_n393_), .Y(men_men_n1240_));
  NOi21      u1212(.An(men_men_n560_), .B(men_men_n580_), .Y(men_men_n1241_));
  NA2        u1213(.A(men_men_n1241_), .B(men_men_n1240_), .Y(men_men_n1242_));
  AN3        u1214(.A(m), .B(l), .C(k), .Y(men_men_n1243_));
  OAI210     u1215(.A0(men_men_n354_), .A1(men_men_n34_), .B0(men_men_n1243_), .Y(men_men_n1244_));
  NA2        u1216(.A(men_men_n204_), .B(men_men_n34_), .Y(men_men_n1245_));
  AO210      u1217(.A0(men_men_n1245_), .A1(men_men_n1244_), .B0(men_men_n327_), .Y(men_men_n1246_));
  NA3        u1218(.A(men_men_n1246_), .B(men_men_n1242_), .C(men_men_n1239_), .Y(men_men_n1247_));
  INV        u1219(.A(men_men_n598_), .Y(men_men_n1248_));
  OAI210     u1220(.A0(men_men_n1231_), .A1(men_men_n592_), .B0(men_men_n1248_), .Y(men_men_n1249_));
  NA2        u1221(.A(men_men_n277_), .B(men_men_n196_), .Y(men_men_n1250_));
  NA2        u1222(.A(men_men_n1250_), .B(men_men_n663_), .Y(men_men_n1251_));
  NO3        u1223(.A(men_men_n827_), .B(men_men_n205_), .C(men_men_n403_), .Y(men_men_n1252_));
  NO2        u1224(.A(men_men_n1252_), .B(men_men_n958_), .Y(men_men_n1253_));
  OAI210     u1225(.A0(men_men_n1228_), .A1(men_men_n321_), .B0(men_men_n675_), .Y(men_men_n1254_));
  NA4        u1226(.A(men_men_n1254_), .B(men_men_n1253_), .C(men_men_n1251_), .D(men_men_n790_), .Y(men_men_n1255_));
  NO3        u1227(.A(men_men_n1255_), .B(men_men_n1249_), .C(men_men_n1247_), .Y(men_men_n1256_));
  NA2        u1228(.A(men_men_n502_), .B(men_men_n54_), .Y(men_men_n1257_));
  NO2        u1229(.A(men_men_n1235_), .B(men_men_n979_), .Y(men_men_n1258_));
  NO2        u1230(.A(men_men_n1258_), .B(men_men_n1168_), .Y(men_men_n1259_));
  NA3        u1231(.A(men_men_n1259_), .B(men_men_n1257_), .C(men_men_n758_), .Y(men_men_n1260_));
  NO2        u1232(.A(men_men_n968_), .B(men_men_n232_), .Y(men_men_n1261_));
  NA2        u1233(.A(men_men_n570_), .B(men_men_n568_), .Y(men_men_n1262_));
  NO3        u1234(.A(men_men_n77_), .B(men_men_n293_), .C(men_men_n43_), .Y(men_men_n1263_));
  NA2        u1235(.A(men_men_n1263_), .B(men_men_n550_), .Y(men_men_n1264_));
  NA3        u1236(.A(men_men_n1264_), .B(men_men_n1262_), .C(men_men_n669_), .Y(men_men_n1265_));
  NA2        u1237(.A(men_men_n1263_), .B(men_men_n818_), .Y(men_men_n1266_));
  NA2        u1238(.A(men_men_n1266_), .B(men_men_n383_), .Y(men_men_n1267_));
  NO3        u1239(.A(men_men_n1267_), .B(men_men_n1265_), .C(men_men_n1260_), .Y(men_men_n1268_));
  NO2        u1240(.A(men_men_n132_), .B(men_men_n43_), .Y(men_men_n1269_));
  NO2        u1241(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n1270_));
  AO220      u1242(.A0(men_men_n1270_), .A1(men_men_n620_), .B0(men_men_n1269_), .B1(men_men_n707_), .Y(men_men_n1271_));
  NA2        u1243(.A(men_men_n1271_), .B(men_men_n335_), .Y(men_men_n1272_));
  INV        u1244(.A(men_men_n136_), .Y(men_men_n1273_));
  NO3        u1245(.A(men_men_n1089_), .B(men_men_n180_), .C(men_men_n85_), .Y(men_men_n1274_));
  AOI220     u1246(.A0(men_men_n1274_), .A1(men_men_n1273_), .B0(men_men_n1263_), .B1(men_men_n970_), .Y(men_men_n1275_));
  NA2        u1247(.A(men_men_n1275_), .B(men_men_n1272_), .Y(men_men_n1276_));
  NO2        u1248(.A(men_men_n611_), .B(men_men_n610_), .Y(men_men_n1277_));
  NO4        u1249(.A(men_men_n1089_), .B(men_men_n1277_), .C(men_men_n178_), .D(men_men_n85_), .Y(men_men_n1278_));
  NO3        u1250(.A(men_men_n1278_), .B(men_men_n1276_), .C(men_men_n636_), .Y(men_men_n1279_));
  NA4        u1251(.A(men_men_n1279_), .B(men_men_n1268_), .C(men_men_n1256_), .D(men_men_n1238_), .Y(men06));
  NO2        u1252(.A(men_men_n404_), .B(men_men_n557_), .Y(men_men_n1281_));
  INV        u1253(.A(men_men_n733_), .Y(men_men_n1282_));
  OAI210     u1254(.A0(men_men_n1282_), .A1(men_men_n267_), .B0(men_men_n1281_), .Y(men_men_n1283_));
  NO2        u1255(.A(men_men_n224_), .B(men_men_n102_), .Y(men_men_n1284_));
  OAI210     u1256(.A0(men_men_n1284_), .A1(men_men_n1274_), .B0(men_men_n379_), .Y(men_men_n1285_));
  NO3        u1257(.A(men_men_n596_), .B(men_men_n813_), .C(men_men_n599_), .Y(men_men_n1286_));
  OR2        u1258(.A(men_men_n1286_), .B(men_men_n890_), .Y(men_men_n1287_));
  NA3        u1259(.A(men_men_n1287_), .B(men_men_n1285_), .C(men_men_n1283_), .Y(men_men_n1288_));
  NO3        u1260(.A(men_men_n1288_), .B(men_men_n1265_), .C(men_men_n256_), .Y(men_men_n1289_));
  NO2        u1261(.A(men_men_n293_), .B(men_men_n43_), .Y(men_men_n1290_));
  AOI210     u1262(.A0(men_men_n1290_), .A1(men_men_n971_), .B0(men_men_n1261_), .Y(men_men_n1291_));
  AOI210     u1263(.A0(men_men_n1290_), .A1(men_men_n554_), .B0(men_men_n1271_), .Y(men_men_n1292_));
  AOI210     u1264(.A0(men_men_n1292_), .A1(men_men_n1291_), .B0(men_men_n333_), .Y(men_men_n1293_));
  INV        u1265(.A(men_men_n673_), .Y(men_men_n1294_));
  NA2        u1266(.A(men_men_n1294_), .B(men_men_n640_), .Y(men_men_n1295_));
  NO2        u1267(.A(men_men_n512_), .B(men_men_n175_), .Y(men_men_n1296_));
  NOi21      u1268(.An(men_men_n138_), .B(men_men_n43_), .Y(men_men_n1297_));
  NO2        u1269(.A(men_men_n604_), .B(men_men_n1113_), .Y(men_men_n1298_));
  OAI210     u1270(.A0(men_men_n459_), .A1(men_men_n247_), .B0(men_men_n910_), .Y(men_men_n1299_));
  NO4        u1271(.A(men_men_n1299_), .B(men_men_n1298_), .C(men_men_n1297_), .D(men_men_n1296_), .Y(men_men_n1300_));
  OR2        u1272(.A(men_men_n597_), .B(men_men_n595_), .Y(men_men_n1301_));
  INV        u1273(.A(men_men_n1301_), .Y(men_men_n1302_));
  NA3        u1274(.A(men_men_n1302_), .B(men_men_n1300_), .C(men_men_n1295_), .Y(men_men_n1303_));
  NO2        u1275(.A(men_men_n749_), .B(men_men_n364_), .Y(men_men_n1304_));
  NO3        u1276(.A(men_men_n675_), .B(men_men_n760_), .C(men_men_n632_), .Y(men_men_n1305_));
  NOi21      u1277(.An(men_men_n1304_), .B(men_men_n1305_), .Y(men_men_n1306_));
  AN2        u1278(.A(men_men_n954_), .B(men_men_n643_), .Y(men_men_n1307_));
  NO4        u1279(.A(men_men_n1307_), .B(men_men_n1306_), .C(men_men_n1303_), .D(men_men_n1293_), .Y(men_men_n1308_));
  NO2        u1280(.A(men_men_n807_), .B(men_men_n275_), .Y(men_men_n1309_));
  OAI220     u1281(.A0(men_men_n733_), .A1(men_men_n45_), .B0(men_men_n224_), .B1(men_men_n613_), .Y(men_men_n1310_));
  OAI210     u1282(.A0(men_men_n275_), .A1(c), .B0(men_men_n639_), .Y(men_men_n1311_));
  AOI220     u1283(.A0(men_men_n1311_), .A1(men_men_n1310_), .B0(men_men_n1309_), .B1(men_men_n267_), .Y(men_men_n1312_));
  OAI220     u1284(.A0(men_men_n700_), .A1(men_men_n247_), .B0(men_men_n508_), .B1(men_men_n512_), .Y(men_men_n1313_));
  OAI210     u1285(.A0(l), .A1(i), .B0(k), .Y(men_men_n1314_));
  NO3        u1286(.A(men_men_n1314_), .B(men_men_n594_), .C(j), .Y(men_men_n1315_));
  NOi21      u1287(.An(men_men_n1315_), .B(men_men_n667_), .Y(men_men_n1316_));
  NO3        u1288(.A(men_men_n1316_), .B(men_men_n1313_), .C(men_men_n1116_), .Y(men_men_n1317_));
  NA3        u1289(.A(men_men_n1317_), .B(men_men_n1312_), .C(men_men_n1208_), .Y(men_men_n1318_));
  NOi31      u1290(.An(men_men_n1286_), .B(men_men_n462_), .C(men_men_n392_), .Y(men_men_n1319_));
  OR3        u1291(.A(men_men_n1319_), .B(men_men_n786_), .C(men_men_n538_), .Y(men_men_n1320_));
  OR3        u1292(.A(men_men_n367_), .B(men_men_n224_), .C(men_men_n613_), .Y(men_men_n1321_));
  AOI210     u1293(.A0(men_men_n570_), .A1(men_men_n445_), .B0(men_men_n369_), .Y(men_men_n1322_));
  NA2        u1294(.A(men_men_n1315_), .B(men_men_n794_), .Y(men_men_n1323_));
  NA4        u1295(.A(men_men_n1323_), .B(men_men_n1322_), .C(men_men_n1321_), .D(men_men_n1320_), .Y(men_men_n1324_));
  NA2        u1296(.A(men_men_n1304_), .B(men_men_n759_), .Y(men_men_n1325_));
  AN2        u1297(.A(men_men_n927_), .B(men_men_n926_), .Y(men_men_n1326_));
  NO4        u1298(.A(men_men_n1326_), .B(men_men_n880_), .C(men_men_n498_), .D(men_men_n477_), .Y(men_men_n1327_));
  NA3        u1299(.A(men_men_n1327_), .B(men_men_n1325_), .C(men_men_n1266_), .Y(men_men_n1328_));
  NAi21      u1300(.An(j), .B(i), .Y(men_men_n1329_));
  NO4        u1301(.A(men_men_n1277_), .B(men_men_n1329_), .C(men_men_n439_), .D(men_men_n235_), .Y(men_men_n1330_));
  NO4        u1302(.A(men_men_n1330_), .B(men_men_n1328_), .C(men_men_n1324_), .D(men_men_n1318_), .Y(men_men_n1331_));
  NA4        u1303(.A(men_men_n1331_), .B(men_men_n1308_), .C(men_men_n1289_), .D(men_men_n1279_), .Y(men07));
  NAi32      u1304(.An(m), .Bn(b), .C(n), .Y(men_men_n1333_));
  NO3        u1305(.A(men_men_n1333_), .B(g), .C(f), .Y(men_men_n1334_));
  OAI210     u1306(.A0(men_men_n315_), .A1(men_men_n479_), .B0(men_men_n1334_), .Y(men_men_n1335_));
  NAi21      u1307(.An(f), .B(c), .Y(men_men_n1336_));
  OR2        u1308(.A(e), .B(d), .Y(men_men_n1337_));
  OAI220     u1309(.A0(men_men_n1337_), .A1(men_men_n1336_), .B0(men_men_n626_), .B1(men_men_n317_), .Y(men_men_n1338_));
  NA3        u1310(.A(men_men_n1338_), .B(men_men_n1053_), .C(men_men_n183_), .Y(men_men_n1339_));
  NOi31      u1311(.An(n), .B(m), .C(b), .Y(men_men_n1340_));
  NO3        u1312(.A(men_men_n133_), .B(men_men_n447_), .C(h), .Y(men_men_n1341_));
  NA2        u1313(.A(men_men_n1339_), .B(men_men_n1335_), .Y(men_men_n1342_));
  NOi41      u1314(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1343_));
  NA2        u1315(.A(men_men_n1091_), .B(men_men_n220_), .Y(men_men_n1344_));
  NO2        u1316(.A(men_men_n1344_), .B(men_men_n57_), .Y(men_men_n1345_));
  NO2        u1317(.A(k), .B(i), .Y(men_men_n1346_));
  NA3        u1318(.A(men_men_n1346_), .B(men_men_n900_), .C(men_men_n183_), .Y(men_men_n1347_));
  NA2        u1319(.A(men_men_n85_), .B(men_men_n43_), .Y(men_men_n1348_));
  NO2        u1320(.A(men_men_n1047_), .B(men_men_n439_), .Y(men_men_n1349_));
  NA3        u1321(.A(men_men_n1349_), .B(men_men_n1348_), .C(men_men_n213_), .Y(men_men_n1350_));
  NO2        u1322(.A(men_men_n1061_), .B(men_men_n300_), .Y(men_men_n1351_));
  NA2        u1323(.A(men_men_n539_), .B(men_men_n78_), .Y(men_men_n1352_));
  NA2        u1324(.A(men_men_n1209_), .B(men_men_n283_), .Y(men_men_n1353_));
  NA4        u1325(.A(men_men_n1353_), .B(men_men_n1352_), .C(men_men_n1350_), .D(men_men_n1347_), .Y(men_men_n1354_));
  NO3        u1326(.A(men_men_n1354_), .B(men_men_n1345_), .C(men_men_n1342_), .Y(men_men_n1355_));
  NO3        u1327(.A(e), .B(d), .C(c), .Y(men_men_n1356_));
  OAI210     u1328(.A0(men_men_n133_), .A1(men_men_n213_), .B0(men_men_n602_), .Y(men_men_n1357_));
  NA2        u1329(.A(men_men_n1357_), .B(men_men_n1356_), .Y(men_men_n1358_));
  INV        u1330(.A(men_men_n1358_), .Y(men_men_n1359_));
  OR2        u1331(.A(h), .B(f), .Y(men_men_n1360_));
  NO3        u1332(.A(n), .B(m), .C(i), .Y(men_men_n1361_));
  OAI210     u1333(.A0(men_men_n1114_), .A1(men_men_n160_), .B0(men_men_n1361_), .Y(men_men_n1362_));
  NO2        u1334(.A(i), .B(g), .Y(men_men_n1363_));
  OR3        u1335(.A(men_men_n1363_), .B(men_men_n1333_), .C(men_men_n68_), .Y(men_men_n1364_));
  OAI220     u1336(.A0(men_men_n1364_), .A1(men_men_n479_), .B0(men_men_n1362_), .B1(men_men_n1360_), .Y(men_men_n1365_));
  NA3        u1337(.A(men_men_n697_), .B(men_men_n683_), .C(men_men_n112_), .Y(men_men_n1366_));
  NA3        u1338(.A(men_men_n1340_), .B(men_men_n1056_), .C(men_men_n671_), .Y(men_men_n1367_));
  AOI210     u1339(.A0(men_men_n1367_), .A1(men_men_n1366_), .B0(men_men_n43_), .Y(men_men_n1368_));
  NA2        u1340(.A(men_men_n1361_), .B(men_men_n638_), .Y(men_men_n1369_));
  NO2        u1341(.A(l), .B(k), .Y(men_men_n1370_));
  NOi41      u1342(.An(men_men_n543_), .B(men_men_n1370_), .C(men_men_n474_), .D(men_men_n439_), .Y(men_men_n1371_));
  NO3        u1343(.A(men_men_n439_), .B(d), .C(c), .Y(men_men_n1372_));
  NO4        u1344(.A(men_men_n1371_), .B(men_men_n1368_), .C(men_men_n1365_), .D(men_men_n1359_), .Y(men_men_n1373_));
  NO2        u1345(.A(men_men_n150_), .B(h), .Y(men_men_n1374_));
  NO2        u1346(.A(men_men_n1071_), .B(l), .Y(men_men_n1375_));
  NO2        u1347(.A(g), .B(c), .Y(men_men_n1376_));
  NA3        u1348(.A(men_men_n1376_), .B(men_men_n144_), .C(men_men_n189_), .Y(men_men_n1377_));
  NO2        u1349(.A(men_men_n1377_), .B(men_men_n1375_), .Y(men_men_n1378_));
  NA2        u1350(.A(men_men_n1378_), .B(men_men_n183_), .Y(men_men_n1379_));
  NO2        u1351(.A(men_men_n450_), .B(a), .Y(men_men_n1380_));
  NA3        u1352(.A(men_men_n1380_), .B(k), .C(men_men_n113_), .Y(men_men_n1381_));
  NO2        u1353(.A(i), .B(h), .Y(men_men_n1382_));
  NA2        u1354(.A(men_men_n1382_), .B(men_men_n220_), .Y(men_men_n1383_));
  AOI210     u1355(.A0(men_men_n1137_), .A1(h), .B0(men_men_n411_), .Y(men_men_n1384_));
  NA2        u1356(.A(men_men_n140_), .B(men_men_n220_), .Y(men_men_n1385_));
  AOI210     u1357(.A0(men_men_n257_), .A1(men_men_n116_), .B0(men_men_n527_), .Y(men_men_n1386_));
  OAI220     u1358(.A0(men_men_n1386_), .A1(men_men_n1383_), .B0(men_men_n1385_), .B1(men_men_n1384_), .Y(men_men_n1387_));
  NO2        u1359(.A(men_men_n756_), .B(men_men_n190_), .Y(men_men_n1388_));
  NOi31      u1360(.An(m), .B(n), .C(b), .Y(men_men_n1389_));
  NOi31      u1361(.An(f), .B(d), .C(c), .Y(men_men_n1390_));
  NA2        u1362(.A(men_men_n1390_), .B(men_men_n1389_), .Y(men_men_n1391_));
  INV        u1363(.A(men_men_n1391_), .Y(men_men_n1392_));
  NO3        u1364(.A(men_men_n1392_), .B(men_men_n1388_), .C(men_men_n1387_), .Y(men_men_n1393_));
  NA2        u1365(.A(men_men_n1082_), .B(men_men_n465_), .Y(men_men_n1394_));
  NO4        u1366(.A(men_men_n1394_), .B(men_men_n1056_), .C(men_men_n439_), .D(men_men_n43_), .Y(men_men_n1395_));
  OAI210     u1367(.A0(men_men_n186_), .A1(men_men_n523_), .B0(men_men_n1057_), .Y(men_men_n1396_));
  NO3        u1368(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1397_));
  INV        u1369(.A(men_men_n1396_), .Y(men_men_n1398_));
  NO2        u1370(.A(men_men_n1398_), .B(men_men_n1395_), .Y(men_men_n1399_));
  AN4        u1371(.A(men_men_n1399_), .B(men_men_n1393_), .C(men_men_n1381_), .D(men_men_n1379_), .Y(men_men_n1400_));
  NA2        u1372(.A(men_men_n1340_), .B(men_men_n376_), .Y(men_men_n1401_));
  NO2        u1373(.A(men_men_n1401_), .B(men_men_n1038_), .Y(men_men_n1402_));
  NA2        u1374(.A(men_men_n1372_), .B(men_men_n214_), .Y(men_men_n1403_));
  NO2        u1375(.A(men_men_n190_), .B(b), .Y(men_men_n1404_));
  AOI220     u1376(.A0(men_men_n1166_), .A1(men_men_n1404_), .B0(men_men_n1090_), .B1(men_men_n1394_), .Y(men_men_n1405_));
  NO2        u1377(.A(i), .B(men_men_n212_), .Y(men_men_n1406_));
  NA4        u1378(.A(men_men_n1142_), .B(men_men_n1406_), .C(men_men_n103_), .D(m), .Y(men_men_n1407_));
  NAi41      u1379(.An(men_men_n1402_), .B(men_men_n1407_), .C(men_men_n1405_), .D(men_men_n1403_), .Y(men_men_n1408_));
  NO4        u1380(.A(men_men_n133_), .B(g), .C(f), .D(e), .Y(men_men_n1409_));
  NA3        u1381(.A(men_men_n1346_), .B(men_men_n284_), .C(h), .Y(men_men_n1410_));
  OR2        u1382(.A(e), .B(a), .Y(men_men_n1411_));
  NO2        u1383(.A(men_men_n1337_), .B(men_men_n1336_), .Y(men_men_n1412_));
  AOI210     u1384(.A0(men_men_n30_), .A1(h), .B0(men_men_n1412_), .Y(men_men_n1413_));
  NO2        u1385(.A(men_men_n1413_), .B(men_men_n1078_), .Y(men_men_n1414_));
  NA2        u1386(.A(men_men_n1343_), .B(men_men_n1370_), .Y(men_men_n1415_));
  INV        u1387(.A(men_men_n1415_), .Y(men_men_n1416_));
  OR3        u1388(.A(men_men_n538_), .B(men_men_n537_), .C(men_men_n112_), .Y(men_men_n1417_));
  NA2        u1389(.A(men_men_n1112_), .B(men_men_n403_), .Y(men_men_n1418_));
  OAI220     u1390(.A0(men_men_n1418_), .A1(men_men_n432_), .B0(men_men_n1417_), .B1(men_men_n293_), .Y(men_men_n1419_));
  AO210      u1391(.A0(men_men_n1419_), .A1(men_men_n116_), .B0(men_men_n1416_), .Y(men_men_n1420_));
  NO3        u1392(.A(men_men_n1420_), .B(men_men_n1414_), .C(men_men_n1408_), .Y(men_men_n1421_));
  NA4        u1393(.A(men_men_n1421_), .B(men_men_n1400_), .C(men_men_n1373_), .D(men_men_n1355_), .Y(men_men_n1422_));
  NA2        u1394(.A(men_men_n376_), .B(men_men_n52_), .Y(men_men_n1423_));
  AOI210     u1395(.A0(men_men_n1423_), .A1(men_men_n1047_), .B0(men_men_n1369_), .Y(men_men_n1424_));
  NO2        u1396(.A(men_men_n1083_), .B(men_men_n1078_), .Y(men_men_n1425_));
  NO2        u1397(.A(men_men_n1425_), .B(men_men_n1424_), .Y(men_men_n1426_));
  NO2        u1398(.A(men_men_n388_), .B(j), .Y(men_men_n1427_));
  NA3        u1399(.A(men_men_n1397_), .B(men_men_n1337_), .C(men_men_n1112_), .Y(men_men_n1428_));
  NAi41      u1400(.An(men_men_n1382_), .B(men_men_n1069_), .C(men_men_n172_), .D(men_men_n153_), .Y(men_men_n1429_));
  NA2        u1401(.A(men_men_n1429_), .B(men_men_n1428_), .Y(men_men_n1430_));
  NA3        u1402(.A(g), .B(men_men_n1427_), .C(men_men_n162_), .Y(men_men_n1431_));
  INV        u1403(.A(men_men_n1431_), .Y(men_men_n1432_));
  NO3        u1404(.A(men_men_n749_), .B(men_men_n178_), .C(men_men_n406_), .Y(men_men_n1433_));
  NO3        u1405(.A(men_men_n1433_), .B(men_men_n1432_), .C(men_men_n1430_), .Y(men_men_n1434_));
  OR2        u1406(.A(n), .B(i), .Y(men_men_n1435_));
  OAI210     u1407(.A0(men_men_n1435_), .A1(men_men_n1068_), .B0(men_men_n47_), .Y(men_men_n1436_));
  AOI220     u1408(.A0(men_men_n1436_), .A1(men_men_n1172_), .B0(men_men_n832_), .B1(men_men_n195_), .Y(men_men_n1437_));
  INV        u1409(.A(men_men_n1437_), .Y(men_men_n1438_));
  NA2        u1410(.A(men_men_n1404_), .B(men_men_n41_), .Y(men_men_n1439_));
  NO2        u1411(.A(men_men_n224_), .B(k), .Y(men_men_n1440_));
  NO2        u1412(.A(men_men_n1439_), .B(men_men_n180_), .Y(men_men_n1441_));
  NO2        u1413(.A(men_men_n1441_), .B(men_men_n1438_), .Y(men_men_n1442_));
  INV        u1414(.A(men_men_n47_), .Y(men_men_n1443_));
  NO3        u1415(.A(men_men_n1093_), .B(men_men_n1337_), .C(men_men_n47_), .Y(men_men_n1444_));
  NA2        u1416(.A(men_men_n1094_), .B(men_men_n1443_), .Y(men_men_n1445_));
  NO2        u1417(.A(men_men_n1078_), .B(h), .Y(men_men_n1446_));
  NA3        u1418(.A(men_men_n1446_), .B(d), .C(men_men_n1039_), .Y(men_men_n1447_));
  OAI220     u1419(.A0(men_men_n1447_), .A1(c), .B0(men_men_n1445_), .B1(j), .Y(men_men_n1448_));
  NA2        u1420(.A(men_men_n183_), .B(men_men_n112_), .Y(men_men_n1449_));
  AOI210     u1421(.A0(men_men_n523_), .A1(h), .B0(men_men_n65_), .Y(men_men_n1450_));
  NA2        u1422(.A(men_men_n1450_), .B(men_men_n1380_), .Y(men_men_n1451_));
  NO2        u1423(.A(men_men_n1329_), .B(men_men_n178_), .Y(men_men_n1452_));
  NOi21      u1424(.An(d), .B(f), .Y(men_men_n1453_));
  NO3        u1425(.A(men_men_n1390_), .B(men_men_n1453_), .C(men_men_n40_), .Y(men_men_n1454_));
  NA2        u1426(.A(men_men_n1454_), .B(men_men_n1452_), .Y(men_men_n1455_));
  NO2        u1427(.A(men_men_n1337_), .B(f), .Y(men_men_n1456_));
  NO2        u1428(.A(men_men_n293_), .B(c), .Y(men_men_n1457_));
  NA2        u1429(.A(men_men_n1457_), .B(men_men_n539_), .Y(men_men_n1458_));
  NA3        u1430(.A(men_men_n1458_), .B(men_men_n1455_), .C(men_men_n1451_), .Y(men_men_n1459_));
  NO2        u1431(.A(men_men_n1459_), .B(men_men_n1448_), .Y(men_men_n1460_));
  NA4        u1432(.A(men_men_n1460_), .B(men_men_n1442_), .C(men_men_n1434_), .D(men_men_n1426_), .Y(men_men_n1461_));
  NO3        u1433(.A(men_men_n1082_), .B(men_men_n1068_), .C(men_men_n40_), .Y(men_men_n1462_));
  NO2        u1434(.A(men_men_n465_), .B(men_men_n293_), .Y(men_men_n1463_));
  OAI210     u1435(.A0(men_men_n1463_), .A1(men_men_n1462_), .B0(men_men_n1351_), .Y(men_men_n1464_));
  OAI210     u1436(.A0(men_men_n1409_), .A1(men_men_n1340_), .B0(men_men_n887_), .Y(men_men_n1465_));
  OAI220     u1437(.A0(men_men_n1035_), .A1(men_men_n133_), .B0(men_men_n664_), .B1(men_men_n178_), .Y(men_men_n1466_));
  NA2        u1438(.A(men_men_n1466_), .B(men_men_n619_), .Y(men_men_n1467_));
  NA3        u1439(.A(men_men_n1467_), .B(men_men_n1465_), .C(men_men_n1464_), .Y(men_men_n1468_));
  NA2        u1440(.A(men_men_n1376_), .B(men_men_n1453_), .Y(men_men_n1469_));
  NO2        u1441(.A(men_men_n1469_), .B(m), .Y(men_men_n1470_));
  NA3        u1442(.A(men_men_n1091_), .B(men_men_n108_), .C(men_men_n220_), .Y(men_men_n1471_));
  NO2        u1443(.A(men_men_n154_), .B(men_men_n185_), .Y(men_men_n1472_));
  OAI210     u1444(.A0(men_men_n1472_), .A1(men_men_n110_), .B0(men_men_n1389_), .Y(men_men_n1473_));
  NA2        u1445(.A(men_men_n1473_), .B(men_men_n1471_), .Y(men_men_n1474_));
  NO3        u1446(.A(men_men_n1474_), .B(men_men_n1470_), .C(men_men_n1468_), .Y(men_men_n1475_));
  NO2        u1447(.A(men_men_n1336_), .B(e), .Y(men_men_n1476_));
  NA2        u1448(.A(men_men_n1476_), .B(men_men_n401_), .Y(men_men_n1477_));
  OAI210     u1449(.A0(men_men_n1456_), .A1(men_men_n1123_), .B0(men_men_n630_), .Y(men_men_n1478_));
  OR3        u1450(.A(men_men_n1440_), .B(men_men_n1209_), .C(men_men_n133_), .Y(men_men_n1479_));
  OAI220     u1451(.A0(men_men_n1479_), .A1(men_men_n1477_), .B0(men_men_n1478_), .B1(men_men_n441_), .Y(men_men_n1480_));
  NO3        u1452(.A(men_men_n1417_), .B(men_men_n348_), .C(a), .Y(men_men_n1481_));
  NO2        u1453(.A(men_men_n1481_), .B(men_men_n1480_), .Y(men_men_n1482_));
  NO2        u1454(.A(men_men_n185_), .B(c), .Y(men_men_n1483_));
  OAI210     u1455(.A0(men_men_n1483_), .A1(men_men_n1476_), .B0(men_men_n183_), .Y(men_men_n1484_));
  AOI220     u1456(.A0(men_men_n1484_), .A1(men_men_n1070_), .B0(men_men_n529_), .B1(men_men_n364_), .Y(men_men_n1485_));
  NA2        u1457(.A(men_men_n537_), .B(g), .Y(men_men_n1486_));
  AOI210     u1458(.A0(men_men_n1486_), .A1(men_men_n1372_), .B0(men_men_n1444_), .Y(men_men_n1487_));
  NA2        u1459(.A(men_men_n1123_), .B(a), .Y(men_men_n1488_));
  OAI220     u1460(.A0(men_men_n1488_), .A1(men_men_n65_), .B0(men_men_n1487_), .B1(men_men_n212_), .Y(men_men_n1489_));
  AOI210     u1461(.A0(men_men_n905_), .A1(men_men_n413_), .B0(men_men_n104_), .Y(men_men_n1490_));
  OR2        u1462(.A(men_men_n1490_), .B(men_men_n537_), .Y(men_men_n1491_));
  NO2        u1463(.A(men_men_n1491_), .B(men_men_n178_), .Y(men_men_n1492_));
  NA4        u1464(.A(men_men_n1091_), .B(men_men_n1088_), .C(men_men_n220_), .D(men_men_n64_), .Y(men_men_n1493_));
  NA2        u1465(.A(men_men_n1341_), .B(men_men_n186_), .Y(men_men_n1494_));
  NO2        u1466(.A(men_men_n47_), .B(l), .Y(men_men_n1495_));
  OAI210     u1467(.A0(men_men_n1411_), .A1(men_men_n867_), .B0(men_men_n479_), .Y(men_men_n1496_));
  OAI210     u1468(.A0(men_men_n1496_), .A1(men_men_n1094_), .B0(men_men_n1495_), .Y(men_men_n1497_));
  NO2        u1469(.A(men_men_n252_), .B(g), .Y(men_men_n1498_));
  NO2        u1470(.A(m), .B(i), .Y(men_men_n1499_));
  BUFFER     u1471(.A(men_men_n1499_), .Y(men_men_n1500_));
  AOI220     u1472(.A0(men_men_n1500_), .A1(men_men_n1374_), .B0(men_men_n1069_), .B1(men_men_n1498_), .Y(men_men_n1501_));
  NA4        u1473(.A(men_men_n1501_), .B(men_men_n1497_), .C(men_men_n1494_), .D(men_men_n1493_), .Y(men_men_n1502_));
  NO4        u1474(.A(men_men_n1502_), .B(men_men_n1492_), .C(men_men_n1489_), .D(men_men_n1485_), .Y(men_men_n1503_));
  NA3        u1475(.A(men_men_n1503_), .B(men_men_n1482_), .C(men_men_n1475_), .Y(men_men_n1504_));
  NA3        u1476(.A(men_men_n960_), .B(men_men_n140_), .C(men_men_n44_), .Y(men_men_n1505_));
  NO2        u1477(.A(men_men_n151_), .B(men_men_n1505_), .Y(men_men_n1506_));
  INV        u1478(.A(men_men_n187_), .Y(men_men_n1507_));
  NA2        u1479(.A(men_men_n1507_), .B(men_men_n1446_), .Y(men_men_n1508_));
  AO210      u1480(.A0(men_men_n134_), .A1(l), .B0(men_men_n1401_), .Y(men_men_n1509_));
  NO2        u1481(.A(men_men_n68_), .B(c), .Y(men_men_n1510_));
  NO4        u1482(.A(men_men_n1360_), .B(men_men_n188_), .C(men_men_n447_), .D(men_men_n43_), .Y(men_men_n1511_));
  AOI210     u1483(.A0(men_men_n1452_), .A1(men_men_n1510_), .B0(men_men_n1511_), .Y(men_men_n1512_));
  NA3        u1484(.A(men_men_n1512_), .B(men_men_n1509_), .C(men_men_n1508_), .Y(men_men_n1513_));
  NO2        u1485(.A(men_men_n1513_), .B(men_men_n1506_), .Y(men_men_n1514_));
  NO4        u1486(.A(men_men_n224_), .B(men_men_n188_), .C(men_men_n257_), .D(k), .Y(men_men_n1515_));
  AOI210     u1487(.A0(men_men_n160_), .A1(men_men_n52_), .B0(men_men_n1476_), .Y(men_men_n1516_));
  NO2        u1488(.A(men_men_n1516_), .B(men_men_n1449_), .Y(men_men_n1517_));
  NO2        u1489(.A(men_men_n1505_), .B(men_men_n110_), .Y(men_men_n1518_));
  NOi21      u1490(.An(men_men_n1341_), .B(e), .Y(men_men_n1519_));
  NO4        u1491(.A(men_men_n1519_), .B(men_men_n1518_), .C(men_men_n1517_), .D(men_men_n1515_), .Y(men_men_n1520_));
  AOI220     u1492(.A0(men_men_n1499_), .A1(men_men_n638_), .B0(men_men_n1053_), .B1(men_men_n163_), .Y(men_men_n1521_));
  NOi31      u1493(.An(men_men_n30_), .B(men_men_n1521_), .C(n), .Y(men_men_n1522_));
  INV        u1494(.A(men_men_n1522_), .Y(men_men_n1523_));
  NA2        u1495(.A(men_men_n55_), .B(a), .Y(men_men_n1524_));
  NO2        u1496(.A(men_men_n1418_), .B(men_men_n1524_), .Y(men_men_n1525_));
  NA4        u1497(.A(men_men_n1539_), .B(men_men_n1523_), .C(men_men_n1520_), .D(men_men_n1514_), .Y(men_men_n1526_));
  OR4        u1498(.A(men_men_n1526_), .B(men_men_n1504_), .C(men_men_n1461_), .D(men_men_n1422_), .Y(men04));
  NOi31      u1499(.An(men_men_n1409_), .B(men_men_n1410_), .C(men_men_n1041_), .Y(men_men_n1528_));
  NA2        u1500(.A(men_men_n1456_), .B(men_men_n832_), .Y(men_men_n1529_));
  NO4        u1501(.A(men_men_n1529_), .B(men_men_n1030_), .C(men_men_n480_), .D(j), .Y(men_men_n1530_));
  OR3        u1502(.A(men_men_n1530_), .B(men_men_n1528_), .C(men_men_n1059_), .Y(men_men_n1531_));
  NO3        u1503(.A(men_men_n1348_), .B(men_men_n89_), .C(k), .Y(men_men_n1532_));
  AOI210     u1504(.A0(men_men_n1532_), .A1(men_men_n1052_), .B0(men_men_n1186_), .Y(men_men_n1533_));
  NA2        u1505(.A(men_men_n1533_), .B(men_men_n1213_), .Y(men_men_n1534_));
  NO4        u1506(.A(men_men_n1534_), .B(men_men_n1531_), .C(men_men_n1067_), .D(men_men_n1046_), .Y(men_men_n1535_));
  NA4        u1507(.A(men_men_n1535_), .B(men_men_n1125_), .C(men_men_n1110_), .D(men_men_n1097_), .Y(men05));
  INV        u1508(.A(men_men_n1525_), .Y(men_men_n1539_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule