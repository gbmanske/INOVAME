library verilog;
use verilog.vl_types.all;
entity contador4bits_vlg_vec_tst is
end contador4bits_vlg_vec_tst;
