//Benchmark atmr_intb_466_0.0313

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n350_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n404_, ori_ori_n405_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n373_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n435_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n363_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  NO3        o027(.A(ori_ori_n49_), .B(x11), .C(x09), .Y(ori_ori_n50_));
  INV        o028(.A(x09), .Y(ori_ori_n51_));
  NO2        o029(.A(x10), .B(x02), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(x07), .Y(ori_ori_n54_));
  OAI210     o032(.A0(ori_ori_n54_), .A1(ori_ori_n50_), .B0(ori_ori_n47_), .Y(ori_ori_n55_));
  NOi21      o033(.An(x01), .B(x09), .Y(ori_ori_n56_));
  INV        o034(.A(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(ori_ori_n51_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n56_), .Y(ori_ori_n59_));
  NA2        o037(.A(x09), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  INV        o038(.A(x07), .Y(ori_ori_n61_));
  INV        o039(.A(ori_ori_n59_), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n63_), .B(ori_ori_n24_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(ori_ori_n62_), .Y(ori_ori_n65_));
  NA2        o043(.A(ori_ori_n61_), .B(ori_ori_n48_), .Y(ori_ori_n66_));
  OAI210     o044(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n66_), .Y(ori_ori_n67_));
  AOI220     o045(.A0(ori_ori_n67_), .A1(ori_ori_n59_), .B0(ori_ori_n65_), .B1(ori_ori_n31_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(ori_ori_n68_), .A1(ori_ori_n55_), .B0(x05), .Y(ori_ori_n69_));
  NA2        o047(.A(x09), .B(x05), .Y(ori_ori_n70_));
  NA2        o048(.A(x10), .B(x06), .Y(ori_ori_n71_));
  NA3        o049(.A(ori_ori_n71_), .B(ori_ori_n70_), .C(ori_ori_n28_), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n61_), .B(ori_ori_n41_), .Y(ori_ori_n73_));
  OAI210     o051(.A0(ori_ori_n72_), .A1(x11), .B0(x03), .Y(ori_ori_n74_));
  NOi31      o052(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n75_));
  INV        o053(.A(x07), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n24_), .Y(ori_ori_n77_));
  NO2        o055(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n78_), .B(ori_ori_n36_), .Y(ori_ori_n79_));
  OAI210     o057(.A0(ori_ori_n78_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n80_));
  AOI210     o058(.A0(ori_ori_n79_), .A1(ori_ori_n48_), .B0(ori_ori_n80_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n82_));
  NO2        o060(.A(x08), .B(x01), .Y(ori_ori_n83_));
  OAI210     o061(.A0(ori_ori_n83_), .A1(ori_ori_n82_), .B0(ori_ori_n35_), .Y(ori_ori_n84_));
  NA2        o062(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n85_));
  NO3        o063(.A(ori_ori_n84_), .B(ori_ori_n81_), .C(ori_ori_n77_), .Y(ori_ori_n86_));
  AN2        o064(.A(ori_ori_n86_), .B(ori_ori_n74_), .Y(ori_ori_n87_));
  INV        o065(.A(ori_ori_n84_), .Y(ori_ori_n88_));
  NA2        o066(.A(x11), .B(x00), .Y(ori_ori_n89_));
  NO2        o067(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n90_));
  NOi21      o068(.An(ori_ori_n89_), .B(ori_ori_n90_), .Y(ori_ori_n91_));
  INV        o069(.A(ori_ori_n91_), .Y(ori_ori_n92_));
  NOi21      o070(.An(x01), .B(x10), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n29_), .B(ori_ori_n57_), .Y(ori_ori_n94_));
  NO3        o072(.A(ori_ori_n94_), .B(ori_ori_n93_), .C(x06), .Y(ori_ori_n95_));
  NA2        o073(.A(ori_ori_n95_), .B(ori_ori_n27_), .Y(ori_ori_n96_));
  OAI210     o074(.A0(ori_ori_n92_), .A1(x07), .B0(ori_ori_n96_), .Y(ori_ori_n97_));
  NO3        o075(.A(ori_ori_n97_), .B(ori_ori_n87_), .C(ori_ori_n69_), .Y(ori01));
  INV        o076(.A(x12), .Y(ori_ori_n99_));
  INV        o077(.A(x13), .Y(ori_ori_n100_));
  NA2        o078(.A(x08), .B(x04), .Y(ori_ori_n101_));
  NO2        o079(.A(x10), .B(x01), .Y(ori_ori_n102_));
  NO2        o080(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n103_), .B(ori_ori_n102_), .Y(ori_ori_n104_));
  NA2        o082(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n105_));
  NO2        o083(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n106_));
  NOi21      o084(.An(ori_ori_n106_), .B(ori_ori_n58_), .Y(ori_ori_n107_));
  INV        o085(.A(x13), .Y(ori_ori_n108_));
  NA2        o086(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n109_));
  NA2        o087(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n110_));
  NO2        o088(.A(ori_ori_n110_), .B(x05), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n35_), .B(ori_ori_n57_), .Y(ori_ori_n112_));
  AOI210     o090(.A0(ori_ori_n57_), .A1(ori_ori_n79_), .B0(ori_ori_n107_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n113_), .B(ori_ori_n71_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n115_));
  NA2        o093(.A(x10), .B(ori_ori_n57_), .Y(ori_ori_n116_));
  NA2        o094(.A(ori_ori_n116_), .B(ori_ori_n115_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n119_));
  NA3        o097(.A(ori_ori_n119_), .B(ori_ori_n118_), .C(x13), .Y(ori_ori_n120_));
  NO2        o098(.A(ori_ori_n60_), .B(x05), .Y(ori_ori_n121_));
  NOi31      o099(.An(ori_ori_n120_), .B(ori_ori_n121_), .C(ori_ori_n117_), .Y(ori_ori_n122_));
  NO3        o100(.A(ori_ori_n122_), .B(x06), .C(x03), .Y(ori_ori_n123_));
  NO2        o101(.A(ori_ori_n123_), .B(ori_ori_n114_), .Y(ori_ori_n124_));
  NA2        o102(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n125_));
  OAI210     o103(.A0(ori_ori_n83_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n126_), .B(ori_ori_n125_), .Y(ori_ori_n127_));
  NO2        o105(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n129_));
  AOI210     o107(.A0(ori_ori_n129_), .A1(ori_ori_n49_), .B0(ori_ori_n128_), .Y(ori_ori_n130_));
  AN2        o108(.A(ori_ori_n130_), .B(ori_ori_n127_), .Y(ori_ori_n131_));
  NO2        o109(.A(x09), .B(x05), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n132_), .B(ori_ori_n47_), .Y(ori_ori_n133_));
  AOI210     o111(.A0(ori_ori_n133_), .A1(ori_ori_n104_), .B0(ori_ori_n49_), .Y(ori_ori_n134_));
  NA2        o112(.A(x09), .B(x00), .Y(ori_ori_n135_));
  NA2        o113(.A(ori_ori_n106_), .B(ori_ori_n135_), .Y(ori_ori_n136_));
  NO2        o114(.A(ori_ori_n134_), .B(ori_ori_n131_), .Y(ori_ori_n137_));
  NO2        o115(.A(x03), .B(x02), .Y(ori_ori_n138_));
  NA2        o116(.A(ori_ori_n84_), .B(ori_ori_n100_), .Y(ori_ori_n139_));
  OAI210     o117(.A0(ori_ori_n139_), .A1(ori_ori_n107_), .B0(ori_ori_n138_), .Y(ori_ori_n140_));
  OA210      o118(.A0(ori_ori_n137_), .A1(x11), .B0(ori_ori_n140_), .Y(ori_ori_n141_));
  OAI210     o119(.A0(ori_ori_n124_), .A1(ori_ori_n23_), .B0(ori_ori_n141_), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n104_), .B(ori_ori_n40_), .Y(ori_ori_n143_));
  NAi21      o121(.An(x06), .B(x10), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n143_), .B(ori_ori_n41_), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n146_));
  NA2        o124(.A(ori_ori_n100_), .B(x01), .Y(ori_ori_n147_));
  NO2        o125(.A(ori_ori_n147_), .B(x08), .Y(ori_ori_n148_));
  OAI210     o126(.A0(x05), .A1(ori_ori_n148_), .B0(ori_ori_n51_), .Y(ori_ori_n149_));
  AOI210     o127(.A0(ori_ori_n149_), .A1(ori_ori_n146_), .B0(ori_ori_n48_), .Y(ori_ori_n150_));
  AOI210     o128(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n151_));
  OAI210     o129(.A0(ori_ori_n150_), .A1(ori_ori_n145_), .B0(ori_ori_n151_), .Y(ori_ori_n152_));
  NA2        o130(.A(x04), .B(x02), .Y(ori_ori_n153_));
  NA2        o131(.A(x10), .B(x05), .Y(ori_ori_n154_));
  NO2        o132(.A(x09), .B(x01), .Y(ori_ori_n155_));
  NO3        o133(.A(ori_ori_n155_), .B(ori_ori_n102_), .C(ori_ori_n31_), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n156_), .B(x00), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n106_), .B(x08), .Y(ori_ori_n158_));
  INV        o136(.A(ori_ori_n157_), .Y(ori_ori_n159_));
  NAi21      o137(.An(ori_ori_n153_), .B(ori_ori_n159_), .Y(ori_ori_n160_));
  INV        o138(.A(ori_ori_n25_), .Y(ori_ori_n161_));
  NAi21      o139(.An(x13), .B(x00), .Y(ori_ori_n162_));
  AOI210     o140(.A0(ori_ori_n29_), .A1(ori_ori_n48_), .B0(ori_ori_n162_), .Y(ori_ori_n163_));
  AOI220     o141(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(ori_ori_n164_));
  OAI210     o142(.A0(ori_ori_n154_), .A1(ori_ori_n35_), .B0(ori_ori_n164_), .Y(ori_ori_n165_));
  AN2        o143(.A(ori_ori_n165_), .B(ori_ori_n163_), .Y(ori_ori_n166_));
  AN2        o144(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n94_), .B(x06), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n162_), .B(ori_ori_n36_), .Y(ori_ori_n169_));
  INV        o147(.A(ori_ori_n169_), .Y(ori_ori_n170_));
  NO2        o148(.A(ori_ori_n168_), .B(ori_ori_n167_), .Y(ori_ori_n171_));
  OAI210     o149(.A0(ori_ori_n171_), .A1(ori_ori_n166_), .B0(ori_ori_n161_), .Y(ori_ori_n172_));
  NOi21      o150(.An(x09), .B(x00), .Y(ori_ori_n173_));
  NO3        o151(.A(ori_ori_n82_), .B(ori_ori_n173_), .C(ori_ori_n47_), .Y(ori_ori_n174_));
  NA2        o152(.A(ori_ori_n174_), .B(ori_ori_n116_), .Y(ori_ori_n175_));
  NA2        o153(.A(x10), .B(x08), .Y(ori_ori_n176_));
  INV        o154(.A(ori_ori_n176_), .Y(ori_ori_n177_));
  NA2        o155(.A(x06), .B(x05), .Y(ori_ori_n178_));
  OAI210     o156(.A0(ori_ori_n178_), .A1(ori_ori_n35_), .B0(ori_ori_n99_), .Y(ori_ori_n179_));
  AOI210     o157(.A0(ori_ori_n177_), .A1(ori_ori_n58_), .B0(ori_ori_n179_), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n180_), .B(ori_ori_n175_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n100_), .B(x12), .Y(ori_ori_n182_));
  AOI210     o160(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n182_), .Y(ori_ori_n183_));
  NA2        o161(.A(ori_ori_n93_), .B(ori_ori_n51_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n185_));
  NA2        o163(.A(ori_ori_n185_), .B(x02), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n183_), .B(ori_ori_n181_), .Y(ori_ori_n187_));
  NA4        o165(.A(ori_ori_n187_), .B(ori_ori_n172_), .C(ori_ori_n160_), .D(ori_ori_n152_), .Y(ori_ori_n188_));
  AOI210     o166(.A0(ori_ori_n142_), .A1(ori_ori_n99_), .B0(ori_ori_n188_), .Y(ori_ori_n189_));
  INV        o167(.A(ori_ori_n72_), .Y(ori_ori_n190_));
  NA2        o168(.A(ori_ori_n190_), .B(ori_ori_n127_), .Y(ori_ori_n191_));
  NA2        o169(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n192_));
  NA2        o170(.A(ori_ori_n192_), .B(ori_ori_n126_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n115_), .B(x06), .Y(ori_ori_n194_));
  INV        o172(.A(ori_ori_n194_), .Y(ori_ori_n195_));
  AOI210     o173(.A0(ori_ori_n195_), .A1(ori_ori_n191_), .B0(x12), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n75_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n93_), .B(x06), .Y(ori_ori_n198_));
  AOI210     o176(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n51_), .Y(ori_ori_n199_));
  NO3        o177(.A(ori_ori_n199_), .B(ori_ori_n198_), .C(ori_ori_n41_), .Y(ori_ori_n200_));
  INV        o178(.A(ori_ori_n129_), .Y(ori_ori_n201_));
  OAI210     o179(.A0(ori_ori_n201_), .A1(ori_ori_n200_), .B0(x02), .Y(ori_ori_n202_));
  AOI210     o180(.A0(ori_ori_n202_), .A1(ori_ori_n57_), .B0(ori_ori_n23_), .Y(ori_ori_n203_));
  OAI210     o181(.A0(ori_ori_n196_), .A1(ori_ori_n57_), .B0(ori_ori_n203_), .Y(ori_ori_n204_));
  INV        o182(.A(ori_ori_n129_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n51_), .B(x03), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n100_), .B(x03), .Y(ori_ori_n207_));
  INV        o185(.A(ori_ori_n144_), .Y(ori_ori_n208_));
  NOi21      o186(.An(x13), .B(x04), .Y(ori_ori_n209_));
  NO3        o187(.A(ori_ori_n209_), .B(ori_ori_n75_), .C(ori_ori_n173_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n210_), .B(x05), .Y(ori_ori_n211_));
  AOI220     o189(.A0(ori_ori_n211_), .A1(ori_ori_n405_), .B0(ori_ori_n208_), .B1(ori_ori_n57_), .Y(ori_ori_n212_));
  INV        o190(.A(ori_ori_n212_), .Y(ori_ori_n213_));
  INV        o191(.A(ori_ori_n90_), .Y(ori_ori_n214_));
  NO2        o192(.A(ori_ori_n214_), .B(x12), .Y(ori_ori_n215_));
  NA2        o193(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n216_));
  NO2        o194(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n217_));
  OAI210     o195(.A0(ori_ori_n217_), .A1(ori_ori_n165_), .B0(ori_ori_n163_), .Y(ori_ori_n218_));
  NO2        o196(.A(x06), .B(x00), .Y(ori_ori_n219_));
  NO2        o197(.A(ori_ori_n219_), .B(ori_ori_n41_), .Y(ori_ori_n220_));
  OAI210     o198(.A0(ori_ori_n101_), .A1(ori_ori_n135_), .B0(ori_ori_n71_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  NA2        o200(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n223_));
  NA2        o201(.A(ori_ori_n223_), .B(x03), .Y(ori_ori_n224_));
  OA210      o202(.A0(ori_ori_n224_), .A1(ori_ori_n222_), .B0(ori_ori_n218_), .Y(ori_ori_n225_));
  NA2        o203(.A(x13), .B(ori_ori_n99_), .Y(ori_ori_n226_));
  NA3        o204(.A(ori_ori_n226_), .B(ori_ori_n179_), .C(ori_ori_n91_), .Y(ori_ori_n227_));
  OAI210     o205(.A0(ori_ori_n225_), .A1(ori_ori_n216_), .B0(ori_ori_n227_), .Y(ori_ori_n228_));
  AOI210     o206(.A0(ori_ori_n215_), .A1(ori_ori_n213_), .B0(ori_ori_n228_), .Y(ori_ori_n229_));
  AOI210     o207(.A0(ori_ori_n229_), .A1(ori_ori_n204_), .B0(x07), .Y(ori_ori_n230_));
  NA2        o208(.A(ori_ori_n70_), .B(ori_ori_n29_), .Y(ori_ori_n231_));
  NOi31      o209(.An(ori_ori_n125_), .B(ori_ori_n209_), .C(ori_ori_n173_), .Y(ori_ori_n232_));
  NO2        o210(.A(ori_ori_n232_), .B(ori_ori_n231_), .Y(ori_ori_n233_));
  NO2        o211(.A(x08), .B(x05), .Y(ori_ori_n234_));
  OAI210     o212(.A0(ori_ori_n75_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n235_));
  INV        o213(.A(ori_ori_n235_), .Y(ori_ori_n236_));
  NO2        o214(.A(x12), .B(x02), .Y(ori_ori_n237_));
  INV        o215(.A(ori_ori_n237_), .Y(ori_ori_n238_));
  NO2        o216(.A(ori_ori_n238_), .B(ori_ori_n214_), .Y(ori_ori_n239_));
  OA210      o217(.A0(ori_ori_n236_), .A1(ori_ori_n233_), .B0(ori_ori_n239_), .Y(ori_ori_n240_));
  NA2        o218(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n241_));
  NO2        o219(.A(ori_ori_n241_), .B(x01), .Y(ori_ori_n242_));
  NOi21      o220(.An(ori_ori_n83_), .B(ori_ori_n109_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n243_), .B(ori_ori_n242_), .Y(ori_ori_n244_));
  AOI210     o222(.A0(ori_ori_n244_), .A1(ori_ori_n120_), .B0(ori_ori_n29_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n100_), .B(x04), .Y(ori_ori_n246_));
  NO2        o224(.A(x02), .B(ori_ori_n108_), .Y(ori_ori_n247_));
  NO3        o225(.A(ori_ori_n89_), .B(x12), .C(x03), .Y(ori_ori_n248_));
  OAI210     o226(.A0(ori_ori_n247_), .A1(ori_ori_n245_), .B0(ori_ori_n248_), .Y(ori_ori_n249_));
  AOI210     o227(.A0(ori_ori_n184_), .A1(ori_ori_n178_), .B0(ori_ori_n101_), .Y(ori_ori_n250_));
  NOi21      o228(.An(ori_ori_n231_), .B(ori_ori_n198_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n252_));
  OAI210     o230(.A0(ori_ori_n251_), .A1(ori_ori_n250_), .B0(ori_ori_n252_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n58_), .B(x05), .Y(ori_ori_n254_));
  NO3        o232(.A(ori_ori_n254_), .B(ori_ori_n199_), .C(ori_ori_n168_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n216_), .B(ori_ori_n28_), .Y(ori_ori_n256_));
  OAI210     o234(.A0(ori_ori_n255_), .A1(ori_ori_n205_), .B0(ori_ori_n256_), .Y(ori_ori_n257_));
  NA3        o235(.A(ori_ori_n257_), .B(ori_ori_n253_), .C(ori_ori_n249_), .Y(ori_ori_n258_));
  NO3        o236(.A(ori_ori_n258_), .B(ori_ori_n240_), .C(ori_ori_n230_), .Y(ori_ori_n259_));
  OAI210     o237(.A0(ori_ori_n189_), .A1(ori_ori_n61_), .B0(ori_ori_n259_), .Y(ori02));
  NOi21      o238(.An(ori_ori_n210_), .B(ori_ori_n155_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n100_), .B(ori_ori_n35_), .Y(ori_ori_n262_));
  NA3        o240(.A(ori_ori_n262_), .B(ori_ori_n177_), .C(ori_ori_n56_), .Y(ori_ori_n263_));
  OAI210     o241(.A0(ori_ori_n261_), .A1(ori_ori_n32_), .B0(ori_ori_n263_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n264_), .B(ori_ori_n154_), .Y(ori_ori_n265_));
  INV        o243(.A(ori_ori_n154_), .Y(ori_ori_n266_));
  INV        o244(.A(ori_ori_n199_), .Y(ori_ori_n267_));
  OAI220     o245(.A0(ori_ori_n267_), .A1(ori_ori_n100_), .B0(ori_ori_n84_), .B1(ori_ori_n51_), .Y(ori_ori_n268_));
  AOI220     o246(.A0(ori_ori_n268_), .A1(ori_ori_n266_), .B0(ori_ori_n139_), .B1(ori_ori_n138_), .Y(ori_ori_n269_));
  AOI210     o247(.A0(ori_ori_n269_), .A1(ori_ori_n265_), .B0(ori_ori_n48_), .Y(ori_ori_n270_));
  NO2        o248(.A(x05), .B(x02), .Y(ori_ori_n271_));
  OAI210     o249(.A0(ori_ori_n193_), .A1(ori_ori_n173_), .B0(ori_ori_n271_), .Y(ori_ori_n272_));
  AOI220     o250(.A0(ori_ori_n234_), .A1(ori_ori_n58_), .B0(ori_ori_n56_), .B1(ori_ori_n36_), .Y(ori_ori_n273_));
  NOi21      o251(.An(ori_ori_n262_), .B(ori_ori_n273_), .Y(ori_ori_n274_));
  AOI210     o252(.A0(ori_ori_n209_), .A1(ori_ori_n78_), .B0(ori_ori_n274_), .Y(ori_ori_n275_));
  AOI210     o253(.A0(ori_ori_n275_), .A1(ori_ori_n272_), .B0(ori_ori_n129_), .Y(ori_ori_n276_));
  NO2        o254(.A(ori_ori_n223_), .B(ori_ori_n47_), .Y(ori_ori_n277_));
  NA2        o255(.A(ori_ori_n277_), .B(ori_ori_n211_), .Y(ori_ori_n278_));
  OAI210     o256(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n279_));
  NA2        o257(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n280_));
  OA210      o258(.A0(ori_ori_n280_), .A1(x08), .B0(ori_ori_n133_), .Y(ori_ori_n281_));
  AOI210     o259(.A0(ori_ori_n281_), .A1(ori_ori_n126_), .B0(ori_ori_n279_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n282_), .B(ori_ori_n94_), .Y(ori_ori_n283_));
  NA3        o261(.A(ori_ori_n94_), .B(ori_ori_n83_), .C(ori_ori_n206_), .Y(ori_ori_n284_));
  NA3        o262(.A(ori_ori_n93_), .B(ori_ori_n82_), .C(ori_ori_n42_), .Y(ori_ori_n285_));
  AOI210     o263(.A0(ori_ori_n285_), .A1(ori_ori_n284_), .B0(x04), .Y(ori_ori_n286_));
  INV        o264(.A(ori_ori_n138_), .Y(ori_ori_n287_));
  NO2        o265(.A(ori_ori_n287_), .B(ori_ori_n117_), .Y(ori_ori_n288_));
  AOI210     o266(.A0(ori_ori_n288_), .A1(x13), .B0(ori_ori_n286_), .Y(ori_ori_n289_));
  NA3        o267(.A(ori_ori_n289_), .B(ori_ori_n283_), .C(ori_ori_n278_), .Y(ori_ori_n290_));
  NO3        o268(.A(ori_ori_n290_), .B(ori_ori_n276_), .C(ori_ori_n270_), .Y(ori_ori_n291_));
  NA2        o269(.A(ori_ori_n128_), .B(x03), .Y(ori_ori_n292_));
  INV        o270(.A(ori_ori_n162_), .Y(ori_ori_n293_));
  AOI220     o271(.A0(x08), .A1(ori_ori_n293_), .B0(ori_ori_n185_), .B1(x08), .Y(ori_ori_n294_));
  OAI210     o272(.A0(ori_ori_n294_), .A1(ori_ori_n254_), .B0(ori_ori_n292_), .Y(ori_ori_n295_));
  NA2        o273(.A(ori_ori_n295_), .B(ori_ori_n102_), .Y(ori_ori_n296_));
  NA2        o274(.A(ori_ori_n153_), .B(ori_ori_n147_), .Y(ori_ori_n297_));
  AN2        o275(.A(ori_ori_n297_), .B(ori_ori_n158_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n118_), .B(ori_ori_n28_), .Y(ori_ori_n299_));
  OAI210     o277(.A0(ori_ori_n299_), .A1(ori_ori_n298_), .B0(ori_ori_n103_), .Y(ori_ori_n300_));
  NA2        o278(.A(ori_ori_n246_), .B(ori_ori_n99_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n99_), .B(ori_ori_n41_), .Y(ori_ori_n302_));
  NA3        o280(.A(ori_ori_n302_), .B(ori_ori_n301_), .C(ori_ori_n117_), .Y(ori_ori_n303_));
  NA4        o281(.A(ori_ori_n303_), .B(ori_ori_n300_), .C(ori_ori_n296_), .D(ori_ori_n48_), .Y(ori_ori_n304_));
  INV        o282(.A(ori_ori_n185_), .Y(ori_ori_n305_));
  NA2        o283(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n306_));
  OAI220     o284(.A0(ori_ori_n306_), .A1(ori_ori_n404_), .B0(ori_ori_n305_), .B1(ori_ori_n59_), .Y(ori_ori_n307_));
  NA2        o285(.A(ori_ori_n307_), .B(x02), .Y(ori_ori_n308_));
  INV        o286(.A(ori_ori_n217_), .Y(ori_ori_n309_));
  NA2        o287(.A(ori_ori_n182_), .B(x04), .Y(ori_ori_n310_));
  NO2        o288(.A(ori_ori_n310_), .B(ori_ori_n309_), .Y(ori_ori_n311_));
  NO3        o289(.A(ori_ori_n164_), .B(x13), .C(ori_ori_n31_), .Y(ori_ori_n312_));
  OAI210     o290(.A0(ori_ori_n312_), .A1(ori_ori_n311_), .B0(ori_ori_n94_), .Y(ori_ori_n313_));
  NO3        o291(.A(ori_ori_n182_), .B(ori_ori_n146_), .C(ori_ori_n52_), .Y(ori_ori_n314_));
  OAI210     o292(.A0(ori_ori_n135_), .A1(ori_ori_n36_), .B0(ori_ori_n99_), .Y(ori_ori_n315_));
  OAI210     o293(.A0(ori_ori_n315_), .A1(ori_ori_n174_), .B0(ori_ori_n314_), .Y(ori_ori_n316_));
  NA4        o294(.A(ori_ori_n316_), .B(ori_ori_n313_), .C(ori_ori_n308_), .D(x06), .Y(ori_ori_n317_));
  NA2        o295(.A(x09), .B(x03), .Y(ori_ori_n318_));
  OAI220     o296(.A0(ori_ori_n318_), .A1(ori_ori_n116_), .B0(ori_ori_n192_), .B1(ori_ori_n63_), .Y(ori_ori_n319_));
  OAI220     o297(.A0(ori_ori_n147_), .A1(x09), .B0(x08), .B1(ori_ori_n41_), .Y(ori_ori_n320_));
  NO3        o298(.A(ori_ori_n254_), .B(ori_ori_n115_), .C(x08), .Y(ori_ori_n321_));
  AOI210     o299(.A0(ori_ori_n320_), .A1(ori_ori_n205_), .B0(ori_ori_n321_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n323_));
  NO3        o301(.A(ori_ori_n106_), .B(ori_ori_n116_), .C(ori_ori_n38_), .Y(ori_ori_n324_));
  AOI210     o302(.A0(ori_ori_n314_), .A1(ori_ori_n323_), .B0(ori_ori_n324_), .Y(ori_ori_n325_));
  OAI210     o303(.A0(ori_ori_n322_), .A1(ori_ori_n28_), .B0(ori_ori_n325_), .Y(ori_ori_n326_));
  AO220      o304(.A0(ori_ori_n326_), .A1(x04), .B0(ori_ori_n319_), .B1(x05), .Y(ori_ori_n327_));
  AOI210     o305(.A0(ori_ori_n317_), .A1(ori_ori_n304_), .B0(ori_ori_n327_), .Y(ori_ori_n328_));
  OAI210     o306(.A0(ori_ori_n291_), .A1(x12), .B0(ori_ori_n328_), .Y(ori03));
  OR2        o307(.A(ori_ori_n42_), .B(ori_ori_n206_), .Y(ori_ori_n330_));
  AOI210     o308(.A0(ori_ori_n139_), .A1(ori_ori_n99_), .B0(ori_ori_n330_), .Y(ori_ori_n331_));
  AO210      o309(.A0(ori_ori_n309_), .A1(ori_ori_n85_), .B0(ori_ori_n310_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n182_), .B(ori_ori_n138_), .Y(ori_ori_n333_));
  NA3        o311(.A(ori_ori_n333_), .B(ori_ori_n332_), .C(ori_ori_n186_), .Y(ori_ori_n334_));
  OAI210     o312(.A0(ori_ori_n334_), .A1(ori_ori_n331_), .B0(x05), .Y(ori_ori_n335_));
  NA2        o313(.A(ori_ori_n330_), .B(x05), .Y(ori_ori_n336_));
  AOI210     o314(.A0(ori_ori_n126_), .A1(ori_ori_n197_), .B0(ori_ori_n336_), .Y(ori_ori_n337_));
  AOI210     o315(.A0(ori_ori_n207_), .A1(ori_ori_n79_), .B0(ori_ori_n111_), .Y(ori_ori_n338_));
  OAI220     o316(.A0(ori_ori_n338_), .A1(ori_ori_n59_), .B0(ori_ori_n280_), .B1(ori_ori_n273_), .Y(ori_ori_n339_));
  OAI210     o317(.A0(ori_ori_n339_), .A1(ori_ori_n337_), .B0(ori_ori_n99_), .Y(ori_ori_n340_));
  AOI210     o318(.A0(ori_ori_n133_), .A1(ori_ori_n60_), .B0(ori_ori_n38_), .Y(ori_ori_n341_));
  NO2        o319(.A(ori_ori_n155_), .B(ori_ori_n121_), .Y(ori_ori_n342_));
  OAI220     o320(.A0(ori_ori_n342_), .A1(ori_ori_n37_), .B0(ori_ori_n136_), .B1(x13), .Y(ori_ori_n343_));
  OAI210     o321(.A0(ori_ori_n343_), .A1(ori_ori_n341_), .B0(x04), .Y(ori_ori_n344_));
  NO3        o322(.A(ori_ori_n302_), .B(ori_ori_n84_), .C(ori_ori_n59_), .Y(ori_ori_n345_));
  AOI210     o323(.A0(ori_ori_n170_), .A1(ori_ori_n99_), .B0(ori_ori_n133_), .Y(ori_ori_n346_));
  OA210      o324(.A0(ori_ori_n148_), .A1(x12), .B0(ori_ori_n121_), .Y(ori_ori_n347_));
  NO3        o325(.A(ori_ori_n347_), .B(ori_ori_n346_), .C(ori_ori_n345_), .Y(ori_ori_n348_));
  NA4        o326(.A(ori_ori_n348_), .B(ori_ori_n344_), .C(ori_ori_n340_), .D(ori_ori_n335_), .Y(ori04));
  NO2        o327(.A(ori_ori_n88_), .B(ori_ori_n39_), .Y(ori_ori_n350_));
  XO2        o328(.A(ori_ori_n350_), .B(ori_ori_n226_), .Y(ori05));
  NO2        o329(.A(ori_ori_n52_), .B(ori_ori_n194_), .Y(ori_ori_n352_));
  AOI210     o330(.A0(ori_ori_n352_), .A1(ori_ori_n279_), .B0(ori_ori_n25_), .Y(ori_ori_n353_));
  NA3        o331(.A(ori_ori_n129_), .B(ori_ori_n118_), .C(ori_ori_n31_), .Y(ori_ori_n354_));
  NO2        o332(.A(ori_ori_n354_), .B(ori_ori_n24_), .Y(ori_ori_n355_));
  OAI210     o333(.A0(ori_ori_n355_), .A1(ori_ori_n353_), .B0(ori_ori_n99_), .Y(ori_ori_n356_));
  NA2        o334(.A(x11), .B(ori_ori_n31_), .Y(ori_ori_n357_));
  NA2        o335(.A(ori_ori_n23_), .B(ori_ori_n28_), .Y(ori_ori_n358_));
  NA2        o336(.A(ori_ori_n231_), .B(x03), .Y(ori_ori_n359_));
  OAI220     o337(.A0(ori_ori_n359_), .A1(ori_ori_n358_), .B0(ori_ori_n357_), .B1(ori_ori_n80_), .Y(ori_ori_n360_));
  OAI210     o338(.A0(ori_ori_n26_), .A1(ori_ori_n99_), .B0(x07), .Y(ori_ori_n361_));
  AOI210     o339(.A0(ori_ori_n360_), .A1(x06), .B0(ori_ori_n361_), .Y(ori_ori_n362_));
  AOI210     o340(.A0(ori_ori_n80_), .A1(ori_ori_n31_), .B0(ori_ori_n52_), .Y(ori_ori_n363_));
  NO3        o341(.A(ori_ori_n363_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n364_));
  OR2        o342(.A(x03), .B(ori_ori_n216_), .Y(ori_ori_n365_));
  NA2        o343(.A(ori_ori_n219_), .B(ori_ori_n214_), .Y(ori_ori_n366_));
  NA2        o344(.A(ori_ori_n366_), .B(ori_ori_n365_), .Y(ori_ori_n367_));
  OAI210     o345(.A0(ori_ori_n367_), .A1(ori_ori_n364_), .B0(ori_ori_n99_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n33_), .B(ori_ori_n99_), .Y(ori_ori_n369_));
  AOI210     o347(.A0(ori_ori_n369_), .A1(ori_ori_n90_), .B0(x07), .Y(ori_ori_n370_));
  AOI220     o348(.A0(ori_ori_n370_), .A1(ori_ori_n368_), .B0(ori_ori_n362_), .B1(ori_ori_n356_), .Y(ori_ori_n371_));
  AOI210     o349(.A0(ori_ori_n241_), .A1(ori_ori_n47_), .B0(x02), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n372_), .B(ori_ori_n100_), .Y(ori_ori_n373_));
  AOI210     o351(.A0(ori_ori_n310_), .A1(ori_ori_n105_), .B0(ori_ori_n237_), .Y(ori_ori_n374_));
  NOi21      o352(.An(ori_ori_n292_), .B(ori_ori_n121_), .Y(ori_ori_n375_));
  NO2        o353(.A(ori_ori_n375_), .B(ori_ori_n238_), .Y(ori_ori_n376_));
  OAI210     o354(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n377_));
  AOI210     o355(.A0(ori_ori_n226_), .A1(ori_ori_n47_), .B0(ori_ori_n377_), .Y(ori_ori_n378_));
  NO4        o356(.A(ori_ori_n378_), .B(ori_ori_n376_), .C(ori_ori_n374_), .D(x08), .Y(ori_ori_n379_));
  NO2        o357(.A(ori_ori_n118_), .B(ori_ori_n28_), .Y(ori_ori_n380_));
  NO2        o358(.A(ori_ori_n380_), .B(ori_ori_n242_), .Y(ori_ori_n381_));
  OR3        o359(.A(ori_ori_n381_), .B(x12), .C(x03), .Y(ori_ori_n382_));
  NA3        o360(.A(ori_ori_n305_), .B(ori_ori_n112_), .C(x12), .Y(ori_ori_n383_));
  AO210      o361(.A0(ori_ori_n305_), .A1(ori_ori_n112_), .B0(ori_ori_n226_), .Y(ori_ori_n384_));
  NA4        o362(.A(ori_ori_n384_), .B(ori_ori_n383_), .C(ori_ori_n382_), .D(x08), .Y(ori_ori_n385_));
  INV        o363(.A(ori_ori_n385_), .Y(ori_ori_n386_));
  AOI210     o364(.A0(ori_ori_n379_), .A1(ori_ori_n373_), .B0(ori_ori_n386_), .Y(ori_ori_n387_));
  INV        o365(.A(x03), .Y(ori_ori_n388_));
  NO2        o366(.A(ori_ori_n132_), .B(ori_ori_n43_), .Y(ori_ori_n389_));
  OAI210     o367(.A0(ori_ori_n389_), .A1(ori_ori_n388_), .B0(ori_ori_n169_), .Y(ori_ori_n390_));
  NA3        o368(.A(ori_ori_n381_), .B(ori_ori_n375_), .C(ori_ori_n301_), .Y(ori_ori_n391_));
  INV        o369(.A(x14), .Y(ori_ori_n392_));
  NO3        o370(.A(ori_ori_n147_), .B(ori_ori_n73_), .C(ori_ori_n57_), .Y(ori_ori_n393_));
  NO2        o371(.A(ori_ori_n393_), .B(ori_ori_n392_), .Y(ori_ori_n394_));
  NA3        o372(.A(ori_ori_n394_), .B(ori_ori_n391_), .C(ori_ori_n390_), .Y(ori_ori_n395_));
  NA2        o373(.A(ori_ori_n369_), .B(ori_ori_n61_), .Y(ori_ori_n396_));
  NOi21      o374(.An(ori_ori_n246_), .B(ori_ori_n136_), .Y(ori_ori_n397_));
  NO2        o375(.A(ori_ori_n44_), .B(x04), .Y(ori_ori_n398_));
  OAI210     o376(.A0(ori_ori_n398_), .A1(ori_ori_n397_), .B0(ori_ori_n99_), .Y(ori_ori_n399_));
  OAI210     o377(.A0(ori_ori_n396_), .A1(ori_ori_n89_), .B0(ori_ori_n399_), .Y(ori_ori_n400_));
  NO4        o378(.A(ori_ori_n400_), .B(ori_ori_n395_), .C(ori_ori_n387_), .D(ori_ori_n371_), .Y(ori06));
  INV        o379(.A(ori_ori_n40_), .Y(ori_ori_n404_));
  INV        o380(.A(x06), .Y(ori_ori_n405_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m046(.A0(mai_mai_n68_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n70_));
  NO2        m048(.A(mai_mai_n61_), .B(mai_mai_n23_), .Y(mai_mai_n71_));
  NA2        m049(.A(x09), .B(x05), .Y(mai_mai_n72_));
  NA2        m050(.A(x10), .B(x06), .Y(mai_mai_n73_));
  NA3        m051(.A(mai_mai_n73_), .B(mai_mai_n72_), .C(mai_mai_n28_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n74_), .A1(mai_mai_n71_), .B0(x03), .Y(mai_mai_n75_));
  NOi31      m053(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n76_));
  NO2        m054(.A(x10), .B(x09), .Y(mai_mai_n77_));
  INV        m055(.A(mai_mai_n24_), .Y(mai_mai_n78_));
  NO2        m056(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n79_));
  NO2        m057(.A(mai_mai_n79_), .B(mai_mai_n36_), .Y(mai_mai_n80_));
  OAI210     m058(.A0(mai_mai_n79_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n81_));
  INV        m059(.A(mai_mai_n81_), .Y(mai_mai_n82_));
  NO2        m060(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n83_));
  NO2        m061(.A(x08), .B(x01), .Y(mai_mai_n84_));
  OAI210     m062(.A0(mai_mai_n84_), .A1(mai_mai_n83_), .B0(mai_mai_n35_), .Y(mai_mai_n85_));
  NA2        m063(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n86_));
  NO3        m064(.A(mai_mai_n85_), .B(mai_mai_n82_), .C(mai_mai_n78_), .Y(mai_mai_n87_));
  AN2        m065(.A(mai_mai_n87_), .B(mai_mai_n75_), .Y(mai_mai_n88_));
  INV        m066(.A(mai_mai_n85_), .Y(mai_mai_n89_));
  NO2        m067(.A(x06), .B(x05), .Y(mai_mai_n90_));
  NA2        m068(.A(x11), .B(x00), .Y(mai_mai_n91_));
  NO2        m069(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n92_));
  NOi21      m070(.An(mai_mai_n91_), .B(mai_mai_n92_), .Y(mai_mai_n93_));
  AOI210     m071(.A0(mai_mai_n90_), .A1(mai_mai_n89_), .B0(mai_mai_n93_), .Y(mai_mai_n94_));
  NOi21      m072(.An(x01), .B(x10), .Y(mai_mai_n95_));
  NO2        m073(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n96_));
  NO3        m074(.A(mai_mai_n96_), .B(mai_mai_n95_), .C(x06), .Y(mai_mai_n97_));
  NA2        m075(.A(mai_mai_n97_), .B(mai_mai_n27_), .Y(mai_mai_n98_));
  OAI210     m076(.A0(mai_mai_n94_), .A1(x07), .B0(mai_mai_n98_), .Y(mai_mai_n99_));
  NO3        m077(.A(mai_mai_n99_), .B(mai_mai_n88_), .C(mai_mai_n70_), .Y(mai01));
  INV        m078(.A(x12), .Y(mai_mai_n101_));
  INV        m079(.A(x13), .Y(mai_mai_n102_));
  NA2        m080(.A(x08), .B(x04), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n57_), .Y(mai_mai_n104_));
  NA2        m082(.A(mai_mai_n104_), .B(mai_mai_n90_), .Y(mai_mai_n105_));
  NA2        m083(.A(mai_mai_n95_), .B(mai_mai_n28_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n106_), .B(mai_mai_n72_), .Y(mai_mai_n107_));
  NO2        m085(.A(x10), .B(x01), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n109_), .B(mai_mai_n108_), .Y(mai_mai_n110_));
  NA2        m088(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n111_));
  NO3        m089(.A(mai_mai_n111_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n112_));
  AOI210     m090(.A0(mai_mai_n112_), .A1(mai_mai_n110_), .B0(mai_mai_n107_), .Y(mai_mai_n113_));
  AOI210     m091(.A0(mai_mai_n113_), .A1(mai_mai_n105_), .B0(mai_mai_n102_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n116_));
  NO2        m094(.A(mai_mai_n102_), .B(mai_mai_n36_), .Y(mai_mai_n117_));
  NA3        m095(.A(mai_mai_n117_), .B(mai_mai_n116_), .C(x06), .Y(mai_mai_n118_));
  INV        m096(.A(mai_mai_n118_), .Y(mai_mai_n119_));
  NO2        m097(.A(mai_mai_n84_), .B(x13), .Y(mai_mai_n120_));
  NA2        m098(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n121_));
  NA2        m099(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n122_));
  NO2        m100(.A(mai_mai_n122_), .B(x05), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n124_));
  NO2        m102(.A(mai_mai_n120_), .B(mai_mai_n73_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n126_));
  NA2        m104(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(mai_mai_n126_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n129_));
  NA2        m107(.A(mai_mai_n36_), .B(x04), .Y(mai_mai_n130_));
  NA3        m108(.A(mai_mai_n130_), .B(mai_mai_n129_), .C(x13), .Y(mai_mai_n131_));
  NO2        m109(.A(mai_mai_n124_), .B(mai_mai_n36_), .Y(mai_mai_n132_));
  NO2        m110(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n133_));
  NOi41      m111(.An(mai_mai_n131_), .B(mai_mai_n133_), .C(mai_mai_n132_), .D(mai_mai_n128_), .Y(mai_mai_n134_));
  NO3        m112(.A(mai_mai_n134_), .B(x06), .C(x03), .Y(mai_mai_n135_));
  NO4        m113(.A(mai_mai_n135_), .B(mai_mai_n125_), .C(mai_mai_n119_), .D(mai_mai_n114_), .Y(mai_mai_n136_));
  NA2        m114(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n137_));
  OAI210     m115(.A0(mai_mai_n84_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n138_));
  NA2        m116(.A(mai_mai_n138_), .B(mai_mai_n137_), .Y(mai_mai_n139_));
  NO2        m117(.A(mai_mai_n35_), .B(mai_mai_n47_), .Y(mai_mai_n140_));
  OA210      m118(.A0(x00), .A1(mai_mai_n77_), .B0(mai_mai_n140_), .Y(mai_mai_n141_));
  NO2        m119(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n143_));
  AN2        m121(.A(mai_mai_n141_), .B(mai_mai_n139_), .Y(mai_mai_n144_));
  NO2        m122(.A(x09), .B(x05), .Y(mai_mai_n145_));
  NA2        m123(.A(mai_mai_n145_), .B(mai_mai_n47_), .Y(mai_mai_n146_));
  AOI210     m124(.A0(mai_mai_n146_), .A1(mai_mai_n110_), .B0(mai_mai_n49_), .Y(mai_mai_n147_));
  NA2        m125(.A(x09), .B(x00), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n115_), .B(mai_mai_n148_), .Y(mai_mai_n149_));
  NA2        m127(.A(mai_mai_n76_), .B(mai_mai_n51_), .Y(mai_mai_n150_));
  AOI210     m128(.A0(mai_mai_n150_), .A1(mai_mai_n149_), .B0(mai_mai_n143_), .Y(mai_mai_n151_));
  NO3        m129(.A(mai_mai_n151_), .B(mai_mai_n147_), .C(mai_mai_n144_), .Y(mai_mai_n152_));
  NO2        m130(.A(x03), .B(x02), .Y(mai_mai_n153_));
  NA2        m131(.A(mai_mai_n85_), .B(mai_mai_n102_), .Y(mai_mai_n154_));
  NA2        m132(.A(mai_mai_n154_), .B(mai_mai_n153_), .Y(mai_mai_n155_));
  OA210      m133(.A0(mai_mai_n152_), .A1(x11), .B0(mai_mai_n155_), .Y(mai_mai_n156_));
  OAI210     m134(.A0(mai_mai_n136_), .A1(mai_mai_n23_), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  NA2        m135(.A(mai_mai_n110_), .B(mai_mai_n40_), .Y(mai_mai_n158_));
  NAi21      m136(.An(x06), .B(x10), .Y(mai_mai_n159_));
  NOi21      m137(.An(x01), .B(x13), .Y(mai_mai_n160_));
  NA2        m138(.A(mai_mai_n160_), .B(mai_mai_n159_), .Y(mai_mai_n161_));
  BUFFER     m139(.A(mai_mai_n161_), .Y(mai_mai_n162_));
  AOI210     m140(.A0(mai_mai_n162_), .A1(mai_mai_n158_), .B0(mai_mai_n41_), .Y(mai_mai_n163_));
  NO2        m141(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n164_));
  NA2        m142(.A(mai_mai_n102_), .B(x01), .Y(mai_mai_n165_));
  NO2        m143(.A(mai_mai_n165_), .B(x08), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n164_), .B(mai_mai_n48_), .Y(mai_mai_n167_));
  AOI210     m145(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n168_));
  OAI210     m146(.A0(mai_mai_n167_), .A1(mai_mai_n163_), .B0(mai_mai_n168_), .Y(mai_mai_n169_));
  NA2        m147(.A(x04), .B(x02), .Y(mai_mai_n170_));
  NA2        m148(.A(x10), .B(x05), .Y(mai_mai_n171_));
  INV        m149(.A(x06), .Y(mai_mai_n172_));
  NO2        m150(.A(x09), .B(x01), .Y(mai_mai_n173_));
  NO3        m151(.A(mai_mai_n173_), .B(mai_mai_n108_), .C(mai_mai_n31_), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n174_), .B(x00), .Y(mai_mai_n175_));
  NO2        m153(.A(mai_mai_n115_), .B(x08), .Y(mai_mai_n176_));
  NA3        m154(.A(mai_mai_n160_), .B(mai_mai_n159_), .C(mai_mai_n51_), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n95_), .B(x05), .Y(mai_mai_n178_));
  OAI210     m156(.A0(mai_mai_n178_), .A1(mai_mai_n117_), .B0(mai_mai_n177_), .Y(mai_mai_n179_));
  AOI210     m157(.A0(mai_mai_n176_), .A1(x06), .B0(mai_mai_n179_), .Y(mai_mai_n180_));
  OAI210     m158(.A0(mai_mai_n180_), .A1(x11), .B0(mai_mai_n175_), .Y(mai_mai_n181_));
  NAi21      m159(.An(mai_mai_n170_), .B(mai_mai_n181_), .Y(mai_mai_n182_));
  INV        m160(.A(mai_mai_n25_), .Y(mai_mai_n183_));
  NAi21      m161(.An(x13), .B(x00), .Y(mai_mai_n184_));
  BUFFER     m162(.A(mai_mai_n72_), .Y(mai_mai_n185_));
  NO2        m163(.A(mai_mai_n96_), .B(x06), .Y(mai_mai_n186_));
  NO2        m164(.A(mai_mai_n184_), .B(mai_mai_n36_), .Y(mai_mai_n187_));
  INV        m165(.A(mai_mai_n187_), .Y(mai_mai_n188_));
  OAI220     m166(.A0(mai_mai_n188_), .A1(mai_mai_n172_), .B0(mai_mai_n186_), .B1(mai_mai_n185_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n189_), .B(mai_mai_n183_), .Y(mai_mai_n190_));
  NOi21      m168(.An(x09), .B(x00), .Y(mai_mai_n191_));
  NO3        m169(.A(mai_mai_n83_), .B(mai_mai_n191_), .C(mai_mai_n47_), .Y(mai_mai_n192_));
  NA2        m170(.A(mai_mai_n192_), .B(mai_mai_n127_), .Y(mai_mai_n193_));
  NA2        m171(.A(x06), .B(x05), .Y(mai_mai_n194_));
  OAI210     m172(.A0(mai_mai_n194_), .A1(mai_mai_n35_), .B0(mai_mai_n101_), .Y(mai_mai_n195_));
  NA2        m173(.A(mai_mai_n101_), .B(mai_mai_n193_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n102_), .B(x12), .Y(mai_mai_n197_));
  AOI210     m175(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n197_), .Y(mai_mai_n198_));
  NA2        m176(.A(mai_mai_n95_), .B(mai_mai_n51_), .Y(mai_mai_n199_));
  NO2        m177(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n200_), .B(x02), .Y(mai_mai_n201_));
  NO2        m179(.A(mai_mai_n201_), .B(mai_mai_n199_), .Y(mai_mai_n202_));
  AOI210     m180(.A0(mai_mai_n198_), .A1(mai_mai_n196_), .B0(mai_mai_n202_), .Y(mai_mai_n203_));
  NA4        m181(.A(mai_mai_n203_), .B(mai_mai_n190_), .C(mai_mai_n182_), .D(mai_mai_n169_), .Y(mai_mai_n204_));
  AOI210     m182(.A0(mai_mai_n157_), .A1(mai_mai_n101_), .B0(mai_mai_n204_), .Y(mai_mai_n205_));
  INV        m183(.A(mai_mai_n74_), .Y(mai_mai_n206_));
  NA2        m184(.A(mai_mai_n206_), .B(mai_mai_n139_), .Y(mai_mai_n207_));
  NA2        m185(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n208_));
  NA2        m186(.A(mai_mai_n208_), .B(mai_mai_n138_), .Y(mai_mai_n209_));
  AOI210     m187(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n210_));
  NO2        m188(.A(mai_mai_n126_), .B(x06), .Y(mai_mai_n211_));
  AOI210     m189(.A0(mai_mai_n210_), .A1(mai_mai_n209_), .B0(mai_mai_n211_), .Y(mai_mai_n212_));
  AOI210     m190(.A0(mai_mai_n212_), .A1(mai_mai_n207_), .B0(x12), .Y(mai_mai_n213_));
  INV        m191(.A(mai_mai_n76_), .Y(mai_mai_n214_));
  NO2        m192(.A(x05), .B(mai_mai_n51_), .Y(mai_mai_n215_));
  OAI210     m193(.A0(mai_mai_n215_), .A1(mai_mai_n161_), .B0(mai_mai_n57_), .Y(mai_mai_n216_));
  NA2        m194(.A(mai_mai_n216_), .B(mai_mai_n214_), .Y(mai_mai_n217_));
  NO2        m195(.A(mai_mai_n95_), .B(x06), .Y(mai_mai_n218_));
  AOI210     m196(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n219_));
  NO3        m197(.A(mai_mai_n219_), .B(mai_mai_n218_), .C(mai_mai_n41_), .Y(mai_mai_n220_));
  NA4        m198(.A(mai_mai_n159_), .B(mai_mai_n56_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n221_));
  NA2        m199(.A(mai_mai_n221_), .B(mai_mai_n143_), .Y(mai_mai_n222_));
  OAI210     m200(.A0(mai_mai_n222_), .A1(mai_mai_n220_), .B0(x02), .Y(mai_mai_n223_));
  AOI210     m201(.A0(mai_mai_n223_), .A1(mai_mai_n217_), .B0(mai_mai_n23_), .Y(mai_mai_n224_));
  OAI210     m202(.A0(mai_mai_n213_), .A1(mai_mai_n57_), .B0(mai_mai_n224_), .Y(mai_mai_n225_));
  INV        m203(.A(mai_mai_n143_), .Y(mai_mai_n226_));
  NO2        m204(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n227_));
  OAI210     m205(.A0(mai_mai_n79_), .A1(mai_mai_n36_), .B0(mai_mai_n121_), .Y(mai_mai_n228_));
  NO2        m206(.A(mai_mai_n102_), .B(x03), .Y(mai_mai_n229_));
  AOI220     m207(.A0(mai_mai_n229_), .A1(mai_mai_n228_), .B0(mai_mai_n76_), .B1(mai_mai_n227_), .Y(mai_mai_n230_));
  NA2        m208(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n231_));
  INV        m209(.A(mai_mai_n159_), .Y(mai_mai_n232_));
  NOi21      m210(.An(x13), .B(x04), .Y(mai_mai_n233_));
  NO3        m211(.A(mai_mai_n233_), .B(mai_mai_n76_), .C(mai_mai_n191_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n234_), .B(x05), .Y(mai_mai_n235_));
  AOI220     m213(.A0(mai_mai_n235_), .A1(mai_mai_n231_), .B0(mai_mai_n232_), .B1(mai_mai_n57_), .Y(mai_mai_n236_));
  OAI210     m214(.A0(mai_mai_n230_), .A1(mai_mai_n226_), .B0(mai_mai_n236_), .Y(mai_mai_n237_));
  INV        m215(.A(mai_mai_n92_), .Y(mai_mai_n238_));
  NO2        m216(.A(mai_mai_n238_), .B(x12), .Y(mai_mai_n239_));
  NA2        m217(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n240_));
  NO2        m218(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n241_));
  AOI210     m219(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n242_));
  NO2        m220(.A(x06), .B(x00), .Y(mai_mai_n243_));
  NO3        m221(.A(mai_mai_n243_), .B(mai_mai_n242_), .C(mai_mai_n41_), .Y(mai_mai_n244_));
  INV        m222(.A(mai_mai_n73_), .Y(mai_mai_n245_));
  NO2        m223(.A(mai_mai_n245_), .B(mai_mai_n244_), .Y(mai_mai_n246_));
  NA2        m224(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n247_), .B(x03), .Y(mai_mai_n248_));
  OR2        m226(.A(mai_mai_n248_), .B(mai_mai_n246_), .Y(mai_mai_n249_));
  NA2        m227(.A(x13), .B(mai_mai_n101_), .Y(mai_mai_n250_));
  NA3        m228(.A(mai_mai_n250_), .B(mai_mai_n195_), .C(mai_mai_n93_), .Y(mai_mai_n251_));
  OAI210     m229(.A0(mai_mai_n249_), .A1(mai_mai_n240_), .B0(mai_mai_n251_), .Y(mai_mai_n252_));
  AOI210     m230(.A0(mai_mai_n239_), .A1(mai_mai_n237_), .B0(mai_mai_n252_), .Y(mai_mai_n253_));
  AOI210     m231(.A0(mai_mai_n253_), .A1(mai_mai_n225_), .B0(x07), .Y(mai_mai_n254_));
  NA2        m232(.A(mai_mai_n72_), .B(mai_mai_n29_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n233_), .B(mai_mai_n191_), .Y(mai_mai_n256_));
  AOI210     m234(.A0(mai_mai_n256_), .A1(mai_mai_n150_), .B0(mai_mai_n255_), .Y(mai_mai_n257_));
  NO2        m235(.A(mai_mai_n102_), .B(x06), .Y(mai_mai_n258_));
  INV        m236(.A(mai_mai_n258_), .Y(mai_mai_n259_));
  NO2        m237(.A(x08), .B(x05), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n260_), .B(mai_mai_n242_), .Y(mai_mai_n261_));
  OAI210     m239(.A0(mai_mai_n76_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n262_));
  OAI210     m240(.A0(mai_mai_n261_), .A1(mai_mai_n259_), .B0(mai_mai_n262_), .Y(mai_mai_n263_));
  NO2        m241(.A(x12), .B(x02), .Y(mai_mai_n264_));
  INV        m242(.A(mai_mai_n264_), .Y(mai_mai_n265_));
  NO2        m243(.A(mai_mai_n265_), .B(mai_mai_n238_), .Y(mai_mai_n266_));
  OA210      m244(.A0(mai_mai_n263_), .A1(mai_mai_n257_), .B0(mai_mai_n266_), .Y(mai_mai_n267_));
  NA2        m245(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n268_));
  NO2        m246(.A(mai_mai_n268_), .B(x01), .Y(mai_mai_n269_));
  INV        m247(.A(mai_mai_n269_), .Y(mai_mai_n270_));
  AOI210     m248(.A0(mai_mai_n270_), .A1(mai_mai_n131_), .B0(mai_mai_n29_), .Y(mai_mai_n271_));
  NA2        m249(.A(mai_mai_n258_), .B(mai_mai_n228_), .Y(mai_mai_n272_));
  NA2        m250(.A(mai_mai_n102_), .B(x04), .Y(mai_mai_n273_));
  OAI210     m251(.A0(x02), .A1(mai_mai_n120_), .B0(mai_mai_n272_), .Y(mai_mai_n274_));
  NO3        m252(.A(mai_mai_n91_), .B(x12), .C(x03), .Y(mai_mai_n275_));
  OAI210     m253(.A0(mai_mai_n274_), .A1(mai_mai_n271_), .B0(mai_mai_n275_), .Y(mai_mai_n276_));
  NOi21      m254(.An(mai_mai_n255_), .B(mai_mai_n218_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n278_));
  NA2        m256(.A(mai_mai_n277_), .B(mai_mai_n278_), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n280_));
  NO3        m258(.A(mai_mai_n280_), .B(mai_mai_n219_), .C(mai_mai_n186_), .Y(mai_mai_n281_));
  NO2        m259(.A(mai_mai_n240_), .B(mai_mai_n28_), .Y(mai_mai_n282_));
  OAI210     m260(.A0(mai_mai_n281_), .A1(mai_mai_n226_), .B0(mai_mai_n282_), .Y(mai_mai_n283_));
  NA3        m261(.A(mai_mai_n283_), .B(mai_mai_n279_), .C(mai_mai_n276_), .Y(mai_mai_n284_));
  NO3        m262(.A(mai_mai_n284_), .B(mai_mai_n267_), .C(mai_mai_n254_), .Y(mai_mai_n285_));
  OAI210     m263(.A0(mai_mai_n205_), .A1(mai_mai_n61_), .B0(mai_mai_n285_), .Y(mai02));
  AOI210     m264(.A0(mai_mai_n137_), .A1(mai_mai_n85_), .B0(mai_mai_n129_), .Y(mai_mai_n287_));
  NOi21      m265(.An(mai_mai_n234_), .B(mai_mai_n173_), .Y(mai_mai_n288_));
  NO2        m266(.A(mai_mai_n288_), .B(mai_mai_n32_), .Y(mai_mai_n289_));
  OAI210     m267(.A0(mai_mai_n289_), .A1(mai_mai_n287_), .B0(mai_mai_n171_), .Y(mai_mai_n290_));
  INV        m268(.A(mai_mai_n171_), .Y(mai_mai_n291_));
  AOI210     m269(.A0(mai_mai_n116_), .A1(mai_mai_n86_), .B0(mai_mai_n219_), .Y(mai_mai_n292_));
  NO2        m270(.A(mai_mai_n292_), .B(mai_mai_n102_), .Y(mai_mai_n293_));
  AOI220     m271(.A0(mai_mai_n293_), .A1(mai_mai_n291_), .B0(mai_mai_n154_), .B1(mai_mai_n153_), .Y(mai_mai_n294_));
  AOI210     m272(.A0(mai_mai_n294_), .A1(mai_mai_n290_), .B0(mai_mai_n48_), .Y(mai_mai_n295_));
  NO2        m273(.A(x05), .B(x02), .Y(mai_mai_n296_));
  OAI210     m274(.A0(mai_mai_n209_), .A1(mai_mai_n191_), .B0(mai_mai_n296_), .Y(mai_mai_n297_));
  AOI220     m275(.A0(mai_mai_n260_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n233_), .B(mai_mai_n79_), .Y(mai_mai_n299_));
  AOI210     m277(.A0(mai_mai_n299_), .A1(mai_mai_n297_), .B0(mai_mai_n143_), .Y(mai_mai_n300_));
  NAi21      m278(.An(mai_mai_n235_), .B(mai_mai_n230_), .Y(mai_mai_n301_));
  NO2        m279(.A(mai_mai_n247_), .B(mai_mai_n47_), .Y(mai_mai_n302_));
  NA2        m280(.A(mai_mai_n302_), .B(mai_mai_n301_), .Y(mai_mai_n303_));
  AN2        m281(.A(mai_mai_n229_), .B(mai_mai_n228_), .Y(mai_mai_n304_));
  OAI210     m282(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n305_));
  NA2        m283(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n306_));
  OA210      m284(.A0(mai_mai_n306_), .A1(x08), .B0(mai_mai_n146_), .Y(mai_mai_n307_));
  AOI210     m285(.A0(mai_mai_n307_), .A1(mai_mai_n138_), .B0(mai_mai_n305_), .Y(mai_mai_n308_));
  OAI210     m286(.A0(mai_mai_n308_), .A1(mai_mai_n304_), .B0(mai_mai_n96_), .Y(mai_mai_n309_));
  NA3        m287(.A(mai_mai_n96_), .B(mai_mai_n84_), .C(mai_mai_n227_), .Y(mai_mai_n310_));
  NA3        m288(.A(mai_mai_n95_), .B(mai_mai_n83_), .C(mai_mai_n42_), .Y(mai_mai_n311_));
  AOI210     m289(.A0(mai_mai_n311_), .A1(mai_mai_n310_), .B0(x04), .Y(mai_mai_n312_));
  INV        m290(.A(mai_mai_n153_), .Y(mai_mai_n313_));
  OAI220     m291(.A0(mai_mai_n261_), .A1(mai_mai_n106_), .B0(mai_mai_n313_), .B1(mai_mai_n128_), .Y(mai_mai_n314_));
  AOI210     m292(.A0(mai_mai_n314_), .A1(x13), .B0(mai_mai_n312_), .Y(mai_mai_n315_));
  NA3        m293(.A(mai_mai_n315_), .B(mai_mai_n309_), .C(mai_mai_n303_), .Y(mai_mai_n316_));
  NO3        m294(.A(mai_mai_n316_), .B(mai_mai_n300_), .C(mai_mai_n295_), .Y(mai_mai_n317_));
  NA2        m295(.A(mai_mai_n142_), .B(x03), .Y(mai_mai_n318_));
  OAI210     m296(.A0(mai_mai_n184_), .A1(mai_mai_n280_), .B0(mai_mai_n318_), .Y(mai_mai_n319_));
  NA2        m297(.A(mai_mai_n319_), .B(mai_mai_n108_), .Y(mai_mai_n320_));
  NA2        m298(.A(mai_mai_n170_), .B(mai_mai_n165_), .Y(mai_mai_n321_));
  AN2        m299(.A(mai_mai_n321_), .B(mai_mai_n176_), .Y(mai_mai_n322_));
  INV        m300(.A(mai_mai_n56_), .Y(mai_mai_n323_));
  OAI220     m301(.A0(mai_mai_n273_), .A1(mai_mai_n323_), .B0(mai_mai_n129_), .B1(mai_mai_n28_), .Y(mai_mai_n324_));
  OAI210     m302(.A0(mai_mai_n324_), .A1(mai_mai_n322_), .B0(mai_mai_n109_), .Y(mai_mai_n325_));
  NA2        m303(.A(mai_mai_n273_), .B(mai_mai_n101_), .Y(mai_mai_n326_));
  NA2        m304(.A(mai_mai_n101_), .B(mai_mai_n41_), .Y(mai_mai_n327_));
  NA3        m305(.A(mai_mai_n327_), .B(mai_mai_n326_), .C(mai_mai_n128_), .Y(mai_mai_n328_));
  NA4        m306(.A(mai_mai_n328_), .B(mai_mai_n325_), .C(mai_mai_n320_), .D(mai_mai_n48_), .Y(mai_mai_n329_));
  INV        m307(.A(mai_mai_n200_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n166_), .B(mai_mai_n40_), .Y(mai_mai_n331_));
  NA2        m309(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n332_));
  OAI220     m310(.A0(mai_mai_n332_), .A1(mai_mai_n331_), .B0(mai_mai_n330_), .B1(mai_mai_n59_), .Y(mai_mai_n333_));
  NA2        m311(.A(mai_mai_n333_), .B(x02), .Y(mai_mai_n334_));
  INV        m312(.A(mai_mai_n241_), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n197_), .B(x04), .Y(mai_mai_n336_));
  NO3        m314(.A(mai_mai_n197_), .B(mai_mai_n164_), .C(mai_mai_n52_), .Y(mai_mai_n337_));
  OAI210     m315(.A0(mai_mai_n148_), .A1(mai_mai_n36_), .B0(mai_mai_n101_), .Y(mai_mai_n338_));
  OAI210     m316(.A0(mai_mai_n338_), .A1(mai_mai_n192_), .B0(mai_mai_n337_), .Y(mai_mai_n339_));
  NA3        m317(.A(mai_mai_n339_), .B(mai_mai_n334_), .C(x06), .Y(mai_mai_n340_));
  NA2        m318(.A(x09), .B(x03), .Y(mai_mai_n341_));
  OAI220     m319(.A0(mai_mai_n341_), .A1(mai_mai_n127_), .B0(mai_mai_n208_), .B1(mai_mai_n64_), .Y(mai_mai_n342_));
  OAI220     m320(.A0(mai_mai_n165_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n343_));
  NO3        m321(.A(mai_mai_n280_), .B(mai_mai_n126_), .C(x08), .Y(mai_mai_n344_));
  AOI210     m322(.A0(mai_mai_n343_), .A1(mai_mai_n226_), .B0(mai_mai_n344_), .Y(mai_mai_n345_));
  NO2        m323(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n346_));
  NO3        m324(.A(mai_mai_n115_), .B(mai_mai_n127_), .C(mai_mai_n38_), .Y(mai_mai_n347_));
  AOI210     m325(.A0(mai_mai_n337_), .A1(mai_mai_n346_), .B0(mai_mai_n347_), .Y(mai_mai_n348_));
  OAI210     m326(.A0(mai_mai_n345_), .A1(mai_mai_n28_), .B0(mai_mai_n348_), .Y(mai_mai_n349_));
  AO220      m327(.A0(mai_mai_n349_), .A1(x04), .B0(mai_mai_n342_), .B1(x05), .Y(mai_mai_n350_));
  AOI210     m328(.A0(mai_mai_n340_), .A1(mai_mai_n329_), .B0(mai_mai_n350_), .Y(mai_mai_n351_));
  OAI210     m329(.A0(mai_mai_n317_), .A1(x12), .B0(mai_mai_n351_), .Y(mai03));
  OR2        m330(.A(mai_mai_n42_), .B(mai_mai_n227_), .Y(mai_mai_n353_));
  AOI210     m331(.A0(mai_mai_n154_), .A1(mai_mai_n101_), .B0(mai_mai_n353_), .Y(mai_mai_n354_));
  AO210      m332(.A0(mai_mai_n335_), .A1(mai_mai_n86_), .B0(mai_mai_n336_), .Y(mai_mai_n355_));
  NA2        m333(.A(mai_mai_n197_), .B(mai_mai_n153_), .Y(mai_mai_n356_));
  NA3        m334(.A(mai_mai_n356_), .B(mai_mai_n355_), .C(mai_mai_n201_), .Y(mai_mai_n357_));
  OAI210     m335(.A0(mai_mai_n357_), .A1(mai_mai_n354_), .B0(x05), .Y(mai_mai_n358_));
  NA2        m336(.A(mai_mai_n353_), .B(x05), .Y(mai_mai_n359_));
  AOI210     m337(.A0(mai_mai_n138_), .A1(mai_mai_n214_), .B0(mai_mai_n359_), .Y(mai_mai_n360_));
  AOI210     m338(.A0(mai_mai_n229_), .A1(mai_mai_n80_), .B0(mai_mai_n123_), .Y(mai_mai_n361_));
  OAI220     m339(.A0(mai_mai_n361_), .A1(mai_mai_n59_), .B0(mai_mai_n306_), .B1(mai_mai_n298_), .Y(mai_mai_n362_));
  OAI210     m340(.A0(mai_mai_n362_), .A1(mai_mai_n360_), .B0(mai_mai_n101_), .Y(mai_mai_n363_));
  AOI210     m341(.A0(mai_mai_n146_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n364_));
  NO2        m342(.A(mai_mai_n173_), .B(mai_mai_n133_), .Y(mai_mai_n365_));
  OAI220     m343(.A0(mai_mai_n365_), .A1(mai_mai_n37_), .B0(mai_mai_n149_), .B1(x13), .Y(mai_mai_n366_));
  OAI210     m344(.A0(mai_mai_n366_), .A1(mai_mai_n364_), .B0(x04), .Y(mai_mai_n367_));
  NO3        m345(.A(mai_mai_n327_), .B(mai_mai_n85_), .C(mai_mai_n59_), .Y(mai_mai_n368_));
  AOI210     m346(.A0(mai_mai_n188_), .A1(mai_mai_n101_), .B0(mai_mai_n146_), .Y(mai_mai_n369_));
  OA210      m347(.A0(mai_mai_n166_), .A1(x12), .B0(mai_mai_n133_), .Y(mai_mai_n370_));
  NO3        m348(.A(mai_mai_n370_), .B(mai_mai_n369_), .C(mai_mai_n368_), .Y(mai_mai_n371_));
  NA4        m349(.A(mai_mai_n371_), .B(mai_mai_n367_), .C(mai_mai_n363_), .D(mai_mai_n358_), .Y(mai04));
  NO2        m350(.A(mai_mai_n89_), .B(mai_mai_n39_), .Y(mai_mai_n373_));
  XO2        m351(.A(mai_mai_n373_), .B(mai_mai_n250_), .Y(mai05));
  AOI210     m352(.A0(mai_mai_n72_), .A1(mai_mai_n52_), .B0(mai_mai_n211_), .Y(mai_mai_n375_));
  AOI210     m353(.A0(mai_mai_n375_), .A1(mai_mai_n305_), .B0(mai_mai_n25_), .Y(mai_mai_n376_));
  NO2        m354(.A(x06), .B(mai_mai_n24_), .Y(mai_mai_n377_));
  OAI210     m355(.A0(mai_mai_n377_), .A1(mai_mai_n376_), .B0(mai_mai_n101_), .Y(mai_mai_n378_));
  OAI210     m356(.A0(mai_mai_n26_), .A1(mai_mai_n101_), .B0(x07), .Y(mai_mai_n379_));
  INV        m357(.A(mai_mai_n379_), .Y(mai_mai_n380_));
  NO2        m358(.A(mai_mai_n435_), .B(mai_mai_n258_), .Y(mai_mai_n381_));
  OR2        m359(.A(mai_mai_n381_), .B(mai_mai_n240_), .Y(mai_mai_n382_));
  NA2        m360(.A(mai_mai_n160_), .B(x05), .Y(mai_mai_n383_));
  NA3        m361(.A(mai_mai_n383_), .B(mai_mai_n243_), .C(mai_mai_n238_), .Y(mai_mai_n384_));
  NO2        m362(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n385_));
  OAI210     m363(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n386_));
  OR3        m364(.A(mai_mai_n386_), .B(mai_mai_n385_), .C(mai_mai_n44_), .Y(mai_mai_n387_));
  NA3        m365(.A(mai_mai_n387_), .B(mai_mai_n384_), .C(mai_mai_n382_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n388_), .B(mai_mai_n101_), .Y(mai_mai_n389_));
  NA2        m367(.A(mai_mai_n33_), .B(mai_mai_n101_), .Y(mai_mai_n390_));
  AOI210     m368(.A0(mai_mai_n390_), .A1(mai_mai_n92_), .B0(x07), .Y(mai_mai_n391_));
  AOI220     m369(.A0(mai_mai_n391_), .A1(mai_mai_n389_), .B0(mai_mai_n380_), .B1(mai_mai_n378_), .Y(mai_mai_n392_));
  NA3        m370(.A(mai_mai_n23_), .B(mai_mai_n61_), .C(mai_mai_n48_), .Y(mai_mai_n393_));
  NO2        m371(.A(x07), .B(mai_mai_n142_), .Y(mai_mai_n394_));
  OR2        m372(.A(mai_mai_n394_), .B(x03), .Y(mai_mai_n395_));
  NA2        m373(.A(mai_mai_n346_), .B(mai_mai_n61_), .Y(mai_mai_n396_));
  NO2        m374(.A(mai_mai_n396_), .B(x11), .Y(mai_mai_n397_));
  NO3        m375(.A(mai_mai_n397_), .B(mai_mai_n145_), .C(mai_mai_n28_), .Y(mai_mai_n398_));
  AOI210     m376(.A0(mai_mai_n398_), .A1(mai_mai_n395_), .B0(mai_mai_n47_), .Y(mai_mai_n399_));
  NO4        m377(.A(mai_mai_n327_), .B(mai_mai_n32_), .C(x11), .D(x09), .Y(mai_mai_n400_));
  OAI210     m378(.A0(mai_mai_n400_), .A1(mai_mai_n399_), .B0(mai_mai_n102_), .Y(mai_mai_n401_));
  AOI210     m379(.A0(mai_mai_n336_), .A1(mai_mai_n111_), .B0(mai_mai_n264_), .Y(mai_mai_n402_));
  NOi21      m380(.An(mai_mai_n318_), .B(mai_mai_n133_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n403_), .B(mai_mai_n265_), .Y(mai_mai_n404_));
  OAI210     m382(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n405_));
  AOI210     m383(.A0(mai_mai_n250_), .A1(mai_mai_n47_), .B0(mai_mai_n405_), .Y(mai_mai_n406_));
  NO4        m384(.A(mai_mai_n406_), .B(mai_mai_n404_), .C(mai_mai_n402_), .D(x08), .Y(mai_mai_n407_));
  NO2        m385(.A(x05), .B(x03), .Y(mai_mai_n408_));
  NO2        m386(.A(x13), .B(x12), .Y(mai_mai_n409_));
  NO2        m387(.A(mai_mai_n129_), .B(mai_mai_n28_), .Y(mai_mai_n410_));
  NO2        m388(.A(mai_mai_n410_), .B(mai_mai_n269_), .Y(mai_mai_n411_));
  NA3        m389(.A(mai_mai_n330_), .B(mai_mai_n124_), .C(x12), .Y(mai_mai_n412_));
  AO210      m390(.A0(mai_mai_n330_), .A1(mai_mai_n124_), .B0(mai_mai_n250_), .Y(mai_mai_n413_));
  NA3        m391(.A(mai_mai_n413_), .B(mai_mai_n412_), .C(x08), .Y(mai_mai_n414_));
  AOI210     m392(.A0(mai_mai_n409_), .A1(mai_mai_n408_), .B0(mai_mai_n414_), .Y(mai_mai_n415_));
  AOI210     m393(.A0(mai_mai_n407_), .A1(mai_mai_n401_), .B0(mai_mai_n415_), .Y(mai_mai_n416_));
  OAI210     m394(.A0(mai_mai_n396_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n417_));
  OAI220     m395(.A0(mai_mai_n171_), .A1(x02), .B0(mai_mai_n145_), .B1(mai_mai_n43_), .Y(mai_mai_n418_));
  OAI210     m396(.A0(mai_mai_n418_), .A1(mai_mai_n417_), .B0(mai_mai_n187_), .Y(mai_mai_n419_));
  NA3        m397(.A(mai_mai_n411_), .B(mai_mai_n403_), .C(mai_mai_n326_), .Y(mai_mai_n420_));
  INV        m398(.A(x14), .Y(mai_mai_n421_));
  NO3        m399(.A(mai_mai_n318_), .B(mai_mai_n106_), .C(x11), .Y(mai_mai_n422_));
  NO3        m400(.A(mai_mai_n393_), .B(mai_mai_n327_), .C(mai_mai_n184_), .Y(mai_mai_n423_));
  NO3        m401(.A(mai_mai_n423_), .B(mai_mai_n422_), .C(mai_mai_n421_), .Y(mai_mai_n424_));
  NA3        m402(.A(mai_mai_n424_), .B(mai_mai_n420_), .C(mai_mai_n419_), .Y(mai_mai_n425_));
  AOI220     m403(.A0(mai_mai_n390_), .A1(mai_mai_n61_), .B0(mai_mai_n410_), .B1(mai_mai_n164_), .Y(mai_mai_n426_));
  NOi21      m404(.An(mai_mai_n273_), .B(mai_mai_n149_), .Y(mai_mai_n427_));
  NA2        m405(.A(mai_mai_n278_), .B(mai_mai_n232_), .Y(mai_mai_n428_));
  OAI210     m406(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n428_), .Y(mai_mai_n429_));
  OAI210     m407(.A0(mai_mai_n429_), .A1(mai_mai_n427_), .B0(mai_mai_n101_), .Y(mai_mai_n430_));
  OAI210     m408(.A0(mai_mai_n426_), .A1(mai_mai_n91_), .B0(mai_mai_n430_), .Y(mai_mai_n431_));
  NO4        m409(.A(mai_mai_n431_), .B(mai_mai_n425_), .C(mai_mai_n416_), .D(mai_mai_n392_), .Y(mai06));
  INV        m410(.A(x02), .Y(mai_mai_n435_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  INV        u027(.A(x09), .Y(men_men_n50_));
  NO2        u028(.A(x10), .B(x02), .Y(men_men_n51_));
  NOi21      u029(.An(x01), .B(x09), .Y(men_men_n52_));
  INV        u030(.A(x00), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n54_));
  NO2        u032(.A(men_men_n54_), .B(men_men_n52_), .Y(men_men_n55_));
  NA2        u033(.A(x09), .B(men_men_n53_), .Y(men_men_n56_));
  INV        u034(.A(x07), .Y(men_men_n57_));
  AOI220     u035(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n57_), .Y(men_men_n58_));
  INV        u036(.A(men_men_n55_), .Y(men_men_n59_));
  NA2        u037(.A(men_men_n29_), .B(x02), .Y(men_men_n60_));
  NA2        u038(.A(men_men_n60_), .B(men_men_n24_), .Y(men_men_n61_));
  OAI220     u039(.A0(men_men_n61_), .A1(men_men_n59_), .B0(men_men_n58_), .B1(men_men_n56_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n57_), .B(men_men_n48_), .Y(men_men_n63_));
  OAI210     u041(.A0(men_men_n30_), .A1(x11), .B0(men_men_n63_), .Y(men_men_n64_));
  AOI220     u042(.A0(men_men_n64_), .A1(men_men_n55_), .B0(men_men_n62_), .B1(men_men_n31_), .Y(men_men_n65_));
  NO2        u043(.A(men_men_n65_), .B(x05), .Y(men_men_n66_));
  NA2        u044(.A(x10), .B(x09), .Y(men_men_n67_));
  NO2        u045(.A(men_men_n57_), .B(men_men_n23_), .Y(men_men_n68_));
  NA2        u046(.A(x09), .B(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x06), .Y(men_men_n70_));
  NA2        u048(.A(men_men_n70_), .B(men_men_n69_), .Y(men_men_n71_));
  NO2        u049(.A(men_men_n57_), .B(men_men_n41_), .Y(men_men_n72_));
  OAI210     u050(.A0(men_men_n71_), .A1(men_men_n68_), .B0(x03), .Y(men_men_n73_));
  NOi31      u051(.An(x08), .B(x04), .C(x00), .Y(men_men_n74_));
  NO2        u052(.A(men_men_n436_), .B(men_men_n24_), .Y(men_men_n75_));
  NO2        u053(.A(x09), .B(men_men_n41_), .Y(men_men_n76_));
  NO2        u054(.A(men_men_n76_), .B(men_men_n36_), .Y(men_men_n77_));
  OAI210     u055(.A0(men_men_n76_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n78_));
  AOI210     u056(.A0(men_men_n77_), .A1(men_men_n48_), .B0(men_men_n78_), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n36_), .B(x00), .Y(men_men_n80_));
  NO2        u058(.A(x08), .B(x01), .Y(men_men_n81_));
  OAI210     u059(.A0(men_men_n81_), .A1(men_men_n80_), .B0(men_men_n35_), .Y(men_men_n82_));
  NA2        u060(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n83_));
  NO3        u061(.A(men_men_n82_), .B(men_men_n79_), .C(men_men_n75_), .Y(men_men_n84_));
  AN2        u062(.A(men_men_n84_), .B(men_men_n73_), .Y(men_men_n85_));
  INV        u063(.A(men_men_n82_), .Y(men_men_n86_));
  NO2        u064(.A(x06), .B(x05), .Y(men_men_n87_));
  NA2        u065(.A(x11), .B(x00), .Y(men_men_n88_));
  NO2        u066(.A(x11), .B(men_men_n47_), .Y(men_men_n89_));
  NOi21      u067(.An(men_men_n88_), .B(men_men_n89_), .Y(men_men_n90_));
  NOi21      u068(.An(x01), .B(x10), .Y(men_men_n91_));
  NO2        u069(.A(men_men_n29_), .B(men_men_n53_), .Y(men_men_n92_));
  NO3        u070(.A(men_men_n92_), .B(men_men_n91_), .C(x06), .Y(men_men_n93_));
  NA2        u071(.A(men_men_n93_), .B(men_men_n27_), .Y(men_men_n94_));
  OAI210     u072(.A0(men_men_n438_), .A1(x07), .B0(men_men_n94_), .Y(men_men_n95_));
  NO3        u073(.A(men_men_n95_), .B(men_men_n85_), .C(men_men_n66_), .Y(men01));
  INV        u074(.A(x12), .Y(men_men_n97_));
  INV        u075(.A(x13), .Y(men_men_n98_));
  NA2        u076(.A(men_men_n87_), .B(x01), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n99_), .B(men_men_n67_), .Y(men_men_n100_));
  NA2        u078(.A(x08), .B(x04), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n101_), .B(men_men_n53_), .Y(men_men_n102_));
  NA2        u080(.A(men_men_n102_), .B(men_men_n100_), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n91_), .B(men_men_n28_), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n104_), .B(men_men_n69_), .Y(men_men_n105_));
  NO2        u083(.A(x10), .B(x01), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n29_), .B(x00), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NA2        u086(.A(x04), .B(men_men_n28_), .Y(men_men_n109_));
  NO3        u087(.A(men_men_n109_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n110_));
  AOI210     u088(.A0(men_men_n110_), .A1(men_men_n108_), .B0(men_men_n105_), .Y(men_men_n111_));
  AOI210     u089(.A0(men_men_n111_), .A1(men_men_n103_), .B0(men_men_n98_), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n52_), .B(x05), .Y(men_men_n113_));
  NOi21      u091(.An(men_men_n113_), .B(men_men_n54_), .Y(men_men_n114_));
  NO2        u092(.A(men_men_n35_), .B(x02), .Y(men_men_n115_));
  NA3        u093(.A(x13), .B(men_men_n115_), .C(x06), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n116_), .B(men_men_n114_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n81_), .B(x13), .Y(men_men_n118_));
  NA2        u096(.A(x09), .B(men_men_n35_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NA2        u098(.A(x13), .B(men_men_n35_), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n121_), .B(x05), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n122_), .B(men_men_n120_), .Y(men_men_n123_));
  NA2        u101(.A(men_men_n35_), .B(men_men_n53_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n124_), .B(men_men_n98_), .Y(men_men_n125_));
  AOI210     u103(.A0(men_men_n125_), .A1(men_men_n77_), .B0(men_men_n114_), .Y(men_men_n126_));
  AOI210     u104(.A0(men_men_n126_), .A1(men_men_n123_), .B0(men_men_n70_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n128_));
  NA2        u106(.A(x10), .B(men_men_n53_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n129_), .B(men_men_n128_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n50_), .B(x05), .Y(men_men_n131_));
  NO3        u109(.A(men_men_n124_), .B(men_men_n76_), .C(men_men_n36_), .Y(men_men_n132_));
  NO2        u110(.A(men_men_n56_), .B(x05), .Y(men_men_n133_));
  NO3        u111(.A(men_men_n133_), .B(men_men_n132_), .C(men_men_n130_), .Y(men_men_n134_));
  NO3        u112(.A(men_men_n134_), .B(x06), .C(x03), .Y(men_men_n135_));
  NO4        u113(.A(men_men_n135_), .B(men_men_n127_), .C(men_men_n117_), .D(men_men_n112_), .Y(men_men_n136_));
  NA2        u114(.A(x13), .B(men_men_n36_), .Y(men_men_n137_));
  OAI210     u115(.A0(men_men_n81_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n138_));
  NA2        u116(.A(men_men_n138_), .B(men_men_n137_), .Y(men_men_n139_));
  NO2        u117(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n140_));
  NA2        u118(.A(men_men_n29_), .B(x06), .Y(men_men_n141_));
  AOI210     u119(.A0(men_men_n141_), .A1(men_men_n49_), .B0(men_men_n140_), .Y(men_men_n142_));
  AN2        u120(.A(men_men_n142_), .B(men_men_n139_), .Y(men_men_n143_));
  NO2        u121(.A(x09), .B(x05), .Y(men_men_n144_));
  NA2        u122(.A(men_men_n144_), .B(men_men_n47_), .Y(men_men_n145_));
  NO2        u123(.A(men_men_n108_), .B(men_men_n49_), .Y(men_men_n146_));
  NA2        u124(.A(x09), .B(x00), .Y(men_men_n147_));
  NA2        u125(.A(men_men_n113_), .B(men_men_n147_), .Y(men_men_n148_));
  NA2        u126(.A(men_men_n74_), .B(men_men_n50_), .Y(men_men_n149_));
  AOI210     u127(.A0(men_men_n149_), .A1(men_men_n148_), .B0(men_men_n141_), .Y(men_men_n150_));
  NO3        u128(.A(men_men_n150_), .B(men_men_n146_), .C(men_men_n143_), .Y(men_men_n151_));
  NO2        u129(.A(x03), .B(x02), .Y(men_men_n152_));
  NA2        u130(.A(men_men_n82_), .B(men_men_n98_), .Y(men_men_n153_));
  OAI210     u131(.A0(men_men_n153_), .A1(men_men_n114_), .B0(men_men_n152_), .Y(men_men_n154_));
  OA210      u132(.A0(men_men_n151_), .A1(x11), .B0(men_men_n154_), .Y(men_men_n155_));
  OAI210     u133(.A0(men_men_n136_), .A1(men_men_n23_), .B0(men_men_n155_), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n108_), .B(men_men_n40_), .Y(men_men_n157_));
  NAi21      u135(.An(x06), .B(x10), .Y(men_men_n158_));
  NOi21      u136(.An(x01), .B(x13), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  OR2        u138(.A(men_men_n160_), .B(x08), .Y(men_men_n161_));
  AOI210     u139(.A0(men_men_n161_), .A1(men_men_n157_), .B0(men_men_n41_), .Y(men_men_n162_));
  NO2        u140(.A(men_men_n29_), .B(x03), .Y(men_men_n163_));
  NA2        u141(.A(men_men_n98_), .B(x01), .Y(men_men_n164_));
  NO2        u142(.A(men_men_n164_), .B(x08), .Y(men_men_n165_));
  OAI210     u143(.A0(x05), .A1(men_men_n165_), .B0(men_men_n50_), .Y(men_men_n166_));
  AOI210     u144(.A0(men_men_n166_), .A1(men_men_n163_), .B0(men_men_n48_), .Y(men_men_n167_));
  AOI210     u145(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n168_));
  OAI210     u146(.A0(men_men_n167_), .A1(men_men_n162_), .B0(men_men_n168_), .Y(men_men_n169_));
  NA2        u147(.A(x04), .B(x02), .Y(men_men_n170_));
  NA2        u148(.A(x10), .B(x05), .Y(men_men_n171_));
  NA2        u149(.A(x09), .B(x06), .Y(men_men_n172_));
  NO2        u150(.A(x09), .B(x01), .Y(men_men_n173_));
  NO2        u151(.A(men_men_n439_), .B(x11), .Y(men_men_n174_));
  NAi21      u152(.An(men_men_n170_), .B(men_men_n174_), .Y(men_men_n175_));
  INV        u153(.A(men_men_n25_), .Y(men_men_n176_));
  NAi21      u154(.An(x13), .B(x00), .Y(men_men_n177_));
  AOI210     u155(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n177_), .Y(men_men_n178_));
  AOI220     u156(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n179_));
  OAI210     u157(.A0(men_men_n171_), .A1(men_men_n35_), .B0(men_men_n179_), .Y(men_men_n180_));
  AN2        u158(.A(men_men_n180_), .B(men_men_n178_), .Y(men_men_n181_));
  NO2        u159(.A(men_men_n177_), .B(men_men_n36_), .Y(men_men_n182_));
  INV        u160(.A(men_men_n182_), .Y(men_men_n183_));
  OAI210     u161(.A0(men_men_n183_), .A1(men_men_n172_), .B0(men_men_n70_), .Y(men_men_n184_));
  OAI210     u162(.A0(men_men_n184_), .A1(men_men_n181_), .B0(men_men_n176_), .Y(men_men_n185_));
  NOi21      u163(.An(x09), .B(x00), .Y(men_men_n186_));
  NO3        u164(.A(men_men_n80_), .B(men_men_n186_), .C(men_men_n47_), .Y(men_men_n187_));
  NA2        u165(.A(men_men_n187_), .B(men_men_n129_), .Y(men_men_n188_));
  NA2        u166(.A(x10), .B(x08), .Y(men_men_n189_));
  INV        u167(.A(men_men_n189_), .Y(men_men_n190_));
  NA2        u168(.A(x06), .B(x05), .Y(men_men_n191_));
  OAI210     u169(.A0(men_men_n191_), .A1(men_men_n35_), .B0(men_men_n97_), .Y(men_men_n192_));
  AOI210     u170(.A0(men_men_n190_), .A1(men_men_n54_), .B0(men_men_n192_), .Y(men_men_n193_));
  NA2        u171(.A(men_men_n193_), .B(men_men_n188_), .Y(men_men_n194_));
  NO2        u172(.A(men_men_n98_), .B(x12), .Y(men_men_n195_));
  AOI210     u173(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n195_), .Y(men_men_n196_));
  NA2        u174(.A(men_men_n91_), .B(men_men_n50_), .Y(men_men_n197_));
  NO2        u175(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n198_));
  NA2        u176(.A(men_men_n198_), .B(x02), .Y(men_men_n199_));
  NO2        u177(.A(men_men_n199_), .B(men_men_n197_), .Y(men_men_n200_));
  AOI210     u178(.A0(men_men_n196_), .A1(men_men_n194_), .B0(men_men_n200_), .Y(men_men_n201_));
  NA4        u179(.A(men_men_n201_), .B(men_men_n185_), .C(men_men_n175_), .D(men_men_n169_), .Y(men_men_n202_));
  AOI210     u180(.A0(men_men_n156_), .A1(men_men_n97_), .B0(men_men_n202_), .Y(men_men_n203_));
  NA2        u181(.A(men_men_n50_), .B(men_men_n47_), .Y(men_men_n204_));
  NA2        u182(.A(men_men_n204_), .B(men_men_n138_), .Y(men_men_n205_));
  AOI210     u183(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n206_));
  NO2        u184(.A(men_men_n128_), .B(x06), .Y(men_men_n207_));
  AOI210     u185(.A0(men_men_n206_), .A1(men_men_n205_), .B0(men_men_n207_), .Y(men_men_n208_));
  NO2        u186(.A(men_men_n208_), .B(x12), .Y(men_men_n209_));
  INV        u187(.A(men_men_n74_), .Y(men_men_n210_));
  NO2        u188(.A(x05), .B(men_men_n50_), .Y(men_men_n211_));
  OAI210     u189(.A0(men_men_n211_), .A1(men_men_n160_), .B0(men_men_n53_), .Y(men_men_n212_));
  NA2        u190(.A(men_men_n212_), .B(men_men_n210_), .Y(men_men_n213_));
  NO2        u191(.A(men_men_n91_), .B(x06), .Y(men_men_n214_));
  NA3        u192(.A(men_men_n52_), .B(men_men_n36_), .C(x04), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n215_), .B(men_men_n141_), .Y(men_men_n216_));
  NA2        u194(.A(men_men_n216_), .B(x02), .Y(men_men_n217_));
  AOI210     u195(.A0(men_men_n217_), .A1(men_men_n213_), .B0(men_men_n23_), .Y(men_men_n218_));
  OAI210     u196(.A0(men_men_n209_), .A1(men_men_n53_), .B0(men_men_n218_), .Y(men_men_n219_));
  INV        u197(.A(men_men_n141_), .Y(men_men_n220_));
  NO2        u198(.A(men_men_n50_), .B(x03), .Y(men_men_n221_));
  OAI210     u199(.A0(men_men_n76_), .A1(men_men_n36_), .B0(men_men_n119_), .Y(men_men_n222_));
  NO2        u200(.A(men_men_n98_), .B(x03), .Y(men_men_n223_));
  AOI220     u201(.A0(men_men_n223_), .A1(men_men_n222_), .B0(men_men_n74_), .B1(men_men_n221_), .Y(men_men_n224_));
  NA2        u202(.A(men_men_n32_), .B(x06), .Y(men_men_n225_));
  INV        u203(.A(men_men_n158_), .Y(men_men_n226_));
  NOi21      u204(.An(x13), .B(x04), .Y(men_men_n227_));
  NO3        u205(.A(men_men_n227_), .B(men_men_n74_), .C(men_men_n186_), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n228_), .B(x05), .Y(men_men_n229_));
  AOI220     u207(.A0(men_men_n229_), .A1(men_men_n225_), .B0(men_men_n226_), .B1(men_men_n53_), .Y(men_men_n230_));
  OAI210     u208(.A0(men_men_n224_), .A1(men_men_n220_), .B0(men_men_n230_), .Y(men_men_n231_));
  INV        u209(.A(men_men_n89_), .Y(men_men_n232_));
  NO2        u210(.A(men_men_n232_), .B(x12), .Y(men_men_n233_));
  NA2        u211(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n234_));
  NO2        u212(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n235_));
  OAI210     u213(.A0(men_men_n235_), .A1(men_men_n180_), .B0(men_men_n178_), .Y(men_men_n236_));
  AOI210     u214(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n237_));
  NA2        u215(.A(men_men_n147_), .B(men_men_n70_), .Y(men_men_n238_));
  INV        u216(.A(men_men_n238_), .Y(men_men_n239_));
  NA2        u217(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n240_));
  NA2        u218(.A(men_men_n240_), .B(x03), .Y(men_men_n241_));
  OA210      u219(.A0(men_men_n241_), .A1(men_men_n239_), .B0(men_men_n236_), .Y(men_men_n242_));
  NA2        u220(.A(x13), .B(men_men_n97_), .Y(men_men_n243_));
  NA3        u221(.A(men_men_n243_), .B(men_men_n192_), .C(men_men_n90_), .Y(men_men_n244_));
  OAI210     u222(.A0(men_men_n242_), .A1(men_men_n234_), .B0(men_men_n244_), .Y(men_men_n245_));
  AOI210     u223(.A0(men_men_n233_), .A1(men_men_n231_), .B0(men_men_n245_), .Y(men_men_n246_));
  AOI210     u224(.A0(men_men_n246_), .A1(men_men_n219_), .B0(x07), .Y(men_men_n247_));
  NA2        u225(.A(men_men_n69_), .B(men_men_n29_), .Y(men_men_n248_));
  BUFFER     u226(.A(men_men_n137_), .Y(men_men_n249_));
  AOI210     u227(.A0(men_men_n249_), .A1(men_men_n149_), .B0(men_men_n248_), .Y(men_men_n250_));
  NO2        u228(.A(men_men_n98_), .B(x06), .Y(men_men_n251_));
  INV        u229(.A(men_men_n251_), .Y(men_men_n252_));
  NO2        u230(.A(x08), .B(x05), .Y(men_men_n253_));
  NO2        u231(.A(men_men_n253_), .B(men_men_n237_), .Y(men_men_n254_));
  NA2        u232(.A(x13), .B(men_men_n31_), .Y(men_men_n255_));
  OAI210     u233(.A0(men_men_n254_), .A1(men_men_n252_), .B0(men_men_n255_), .Y(men_men_n256_));
  NO2        u234(.A(x12), .B(x02), .Y(men_men_n257_));
  INV        u235(.A(men_men_n257_), .Y(men_men_n258_));
  NO2        u236(.A(men_men_n258_), .B(men_men_n232_), .Y(men_men_n259_));
  OA210      u237(.A0(men_men_n256_), .A1(men_men_n250_), .B0(men_men_n259_), .Y(men_men_n260_));
  NA2        u238(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n261_));
  NO2        u239(.A(men_men_n261_), .B(x01), .Y(men_men_n262_));
  NOi21      u240(.An(men_men_n81_), .B(men_men_n119_), .Y(men_men_n263_));
  NA2        u241(.A(men_men_n251_), .B(men_men_n222_), .Y(men_men_n264_));
  NA2        u242(.A(men_men_n98_), .B(x04), .Y(men_men_n265_));
  NA2        u243(.A(men_men_n265_), .B(men_men_n28_), .Y(men_men_n266_));
  OAI210     u244(.A0(men_men_n266_), .A1(men_men_n118_), .B0(men_men_n264_), .Y(men_men_n267_));
  NO3        u245(.A(men_men_n88_), .B(x12), .C(x03), .Y(men_men_n268_));
  OAI210     u246(.A0(men_men_n267_), .A1(men_men_n263_), .B0(men_men_n268_), .Y(men_men_n269_));
  AOI210     u247(.A0(men_men_n197_), .A1(men_men_n191_), .B0(men_men_n101_), .Y(men_men_n270_));
  NOi21      u248(.An(men_men_n248_), .B(men_men_n214_), .Y(men_men_n271_));
  NO2        u249(.A(men_men_n25_), .B(x00), .Y(men_men_n272_));
  OAI210     u250(.A0(men_men_n271_), .A1(men_men_n270_), .B0(men_men_n272_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n54_), .B(x05), .Y(men_men_n274_));
  NO2        u252(.A(men_men_n234_), .B(men_men_n28_), .Y(men_men_n275_));
  NA2        u253(.A(men_men_n220_), .B(men_men_n275_), .Y(men_men_n276_));
  NA3        u254(.A(men_men_n276_), .B(men_men_n273_), .C(men_men_n269_), .Y(men_men_n277_));
  NO3        u255(.A(men_men_n277_), .B(men_men_n260_), .C(men_men_n247_), .Y(men_men_n278_));
  OAI210     u256(.A0(men_men_n203_), .A1(men_men_n57_), .B0(men_men_n278_), .Y(men02));
  AOI210     u257(.A0(men_men_n137_), .A1(men_men_n82_), .B0(men_men_n131_), .Y(men_men_n280_));
  NOi21      u258(.An(men_men_n228_), .B(men_men_n173_), .Y(men_men_n281_));
  NO2        u259(.A(men_men_n98_), .B(men_men_n35_), .Y(men_men_n282_));
  NA3        u260(.A(men_men_n282_), .B(men_men_n190_), .C(men_men_n52_), .Y(men_men_n283_));
  OAI210     u261(.A0(men_men_n281_), .A1(men_men_n32_), .B0(men_men_n283_), .Y(men_men_n284_));
  OAI210     u262(.A0(men_men_n284_), .A1(men_men_n280_), .B0(men_men_n171_), .Y(men_men_n285_));
  INV        u263(.A(men_men_n171_), .Y(men_men_n286_));
  AOI210     u264(.A0(men_men_n115_), .A1(men_men_n83_), .B0(x09), .Y(men_men_n287_));
  OAI220     u265(.A0(men_men_n287_), .A1(men_men_n98_), .B0(men_men_n82_), .B1(men_men_n50_), .Y(men_men_n288_));
  AOI220     u266(.A0(men_men_n288_), .A1(men_men_n286_), .B0(men_men_n153_), .B1(men_men_n152_), .Y(men_men_n289_));
  AOI210     u267(.A0(men_men_n289_), .A1(men_men_n285_), .B0(men_men_n48_), .Y(men_men_n290_));
  NO2        u268(.A(x05), .B(x02), .Y(men_men_n291_));
  OAI210     u269(.A0(men_men_n205_), .A1(men_men_n186_), .B0(men_men_n291_), .Y(men_men_n292_));
  AOI220     u270(.A0(men_men_n253_), .A1(men_men_n54_), .B0(men_men_n52_), .B1(men_men_n36_), .Y(men_men_n293_));
  NOi21      u271(.An(men_men_n282_), .B(men_men_n293_), .Y(men_men_n294_));
  INV        u272(.A(men_men_n294_), .Y(men_men_n295_));
  AOI210     u273(.A0(men_men_n295_), .A1(men_men_n292_), .B0(men_men_n141_), .Y(men_men_n296_));
  NAi21      u274(.An(men_men_n229_), .B(men_men_n224_), .Y(men_men_n297_));
  NO2        u275(.A(men_men_n240_), .B(men_men_n47_), .Y(men_men_n298_));
  NA2        u276(.A(men_men_n298_), .B(men_men_n297_), .Y(men_men_n299_));
  AN2        u277(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n300_));
  OAI210     u278(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n301_));
  NA2        u279(.A(x13), .B(men_men_n28_), .Y(men_men_n302_));
  BUFFER     u280(.A(men_men_n145_), .Y(men_men_n303_));
  AOI210     u281(.A0(men_men_n303_), .A1(men_men_n138_), .B0(men_men_n301_), .Y(men_men_n304_));
  OAI210     u282(.A0(men_men_n304_), .A1(men_men_n300_), .B0(men_men_n92_), .Y(men_men_n305_));
  INV        u283(.A(men_men_n152_), .Y(men_men_n306_));
  OAI220     u284(.A0(men_men_n254_), .A1(men_men_n104_), .B0(men_men_n306_), .B1(men_men_n130_), .Y(men_men_n307_));
  NA2        u285(.A(men_men_n307_), .B(x13), .Y(men_men_n308_));
  NA3        u286(.A(men_men_n308_), .B(men_men_n305_), .C(men_men_n299_), .Y(men_men_n309_));
  NO3        u287(.A(men_men_n309_), .B(men_men_n296_), .C(men_men_n290_), .Y(men_men_n310_));
  NA2        u288(.A(men_men_n140_), .B(x03), .Y(men_men_n311_));
  INV        u289(.A(men_men_n177_), .Y(men_men_n312_));
  OAI210     u290(.A0(men_men_n50_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n313_));
  AOI220     u291(.A0(men_men_n313_), .A1(men_men_n312_), .B0(men_men_n198_), .B1(x08), .Y(men_men_n314_));
  OAI210     u292(.A0(men_men_n314_), .A1(men_men_n274_), .B0(men_men_n311_), .Y(men_men_n315_));
  NA2        u293(.A(men_men_n315_), .B(men_men_n106_), .Y(men_men_n316_));
  INV        u294(.A(men_men_n52_), .Y(men_men_n317_));
  OAI220     u295(.A0(men_men_n265_), .A1(men_men_n317_), .B0(men_men_n131_), .B1(men_men_n28_), .Y(men_men_n318_));
  NA2        u296(.A(men_men_n318_), .B(men_men_n107_), .Y(men_men_n319_));
  NA2        u297(.A(men_men_n265_), .B(men_men_n97_), .Y(men_men_n320_));
  NA2        u298(.A(men_men_n97_), .B(men_men_n41_), .Y(men_men_n321_));
  NA3        u299(.A(men_men_n321_), .B(men_men_n320_), .C(men_men_n130_), .Y(men_men_n322_));
  NA4        u300(.A(men_men_n322_), .B(men_men_n319_), .C(men_men_n316_), .D(men_men_n48_), .Y(men_men_n323_));
  INV        u301(.A(men_men_n198_), .Y(men_men_n324_));
  NO2        u302(.A(men_men_n165_), .B(men_men_n40_), .Y(men_men_n325_));
  NA2        u303(.A(men_men_n32_), .B(x05), .Y(men_men_n326_));
  OAI220     u304(.A0(men_men_n326_), .A1(men_men_n325_), .B0(men_men_n324_), .B1(men_men_n55_), .Y(men_men_n327_));
  NA2        u305(.A(men_men_n327_), .B(x02), .Y(men_men_n328_));
  INV        u306(.A(men_men_n235_), .Y(men_men_n329_));
  NA2        u307(.A(men_men_n195_), .B(x04), .Y(men_men_n330_));
  NO2        u308(.A(men_men_n330_), .B(men_men_n329_), .Y(men_men_n331_));
  NO3        u309(.A(men_men_n179_), .B(x13), .C(men_men_n31_), .Y(men_men_n332_));
  OAI210     u310(.A0(men_men_n332_), .A1(men_men_n331_), .B0(men_men_n92_), .Y(men_men_n333_));
  NO3        u311(.A(men_men_n195_), .B(men_men_n163_), .C(men_men_n51_), .Y(men_men_n334_));
  OAI210     u312(.A0(men_men_n147_), .A1(men_men_n36_), .B0(men_men_n97_), .Y(men_men_n335_));
  OAI210     u313(.A0(men_men_n335_), .A1(men_men_n187_), .B0(men_men_n334_), .Y(men_men_n336_));
  NA4        u314(.A(men_men_n336_), .B(men_men_n333_), .C(men_men_n328_), .D(x06), .Y(men_men_n337_));
  NA2        u315(.A(x09), .B(x03), .Y(men_men_n338_));
  OAI220     u316(.A0(men_men_n338_), .A1(men_men_n129_), .B0(men_men_n204_), .B1(men_men_n60_), .Y(men_men_n339_));
  AN2        u317(.A(men_men_n339_), .B(x05), .Y(men_men_n340_));
  AOI210     u318(.A0(men_men_n337_), .A1(men_men_n323_), .B0(men_men_n340_), .Y(men_men_n341_));
  OAI210     u319(.A0(men_men_n310_), .A1(x12), .B0(men_men_n341_), .Y(men03));
  OR2        u320(.A(men_men_n42_), .B(men_men_n221_), .Y(men_men_n343_));
  AOI210     u321(.A0(men_men_n153_), .A1(men_men_n97_), .B0(men_men_n343_), .Y(men_men_n344_));
  AO210      u322(.A0(men_men_n329_), .A1(men_men_n83_), .B0(men_men_n330_), .Y(men_men_n345_));
  NA2        u323(.A(men_men_n195_), .B(men_men_n152_), .Y(men_men_n346_));
  NA3        u324(.A(men_men_n346_), .B(men_men_n345_), .C(men_men_n199_), .Y(men_men_n347_));
  OAI210     u325(.A0(men_men_n347_), .A1(men_men_n344_), .B0(x05), .Y(men_men_n348_));
  NA2        u326(.A(men_men_n343_), .B(x05), .Y(men_men_n349_));
  AOI210     u327(.A0(men_men_n138_), .A1(men_men_n210_), .B0(men_men_n349_), .Y(men_men_n350_));
  AOI210     u328(.A0(men_men_n223_), .A1(men_men_n77_), .B0(men_men_n122_), .Y(men_men_n351_));
  OAI220     u329(.A0(men_men_n351_), .A1(men_men_n55_), .B0(men_men_n302_), .B1(men_men_n293_), .Y(men_men_n352_));
  OAI210     u330(.A0(men_men_n352_), .A1(men_men_n350_), .B0(men_men_n97_), .Y(men_men_n353_));
  AOI210     u331(.A0(men_men_n145_), .A1(men_men_n56_), .B0(men_men_n38_), .Y(men_men_n354_));
  NO2        u332(.A(men_men_n173_), .B(men_men_n133_), .Y(men_men_n355_));
  OAI220     u333(.A0(men_men_n355_), .A1(men_men_n37_), .B0(men_men_n148_), .B1(x13), .Y(men_men_n356_));
  OAI210     u334(.A0(men_men_n356_), .A1(men_men_n354_), .B0(x04), .Y(men_men_n357_));
  NO3        u335(.A(men_men_n321_), .B(men_men_n82_), .C(men_men_n55_), .Y(men_men_n358_));
  AOI210     u336(.A0(men_men_n183_), .A1(men_men_n97_), .B0(men_men_n145_), .Y(men_men_n359_));
  OA210      u337(.A0(men_men_n165_), .A1(x12), .B0(men_men_n133_), .Y(men_men_n360_));
  NO3        u338(.A(men_men_n360_), .B(men_men_n359_), .C(men_men_n358_), .Y(men_men_n361_));
  NA4        u339(.A(men_men_n361_), .B(men_men_n357_), .C(men_men_n353_), .D(men_men_n348_), .Y(men04));
  NO2        u340(.A(men_men_n86_), .B(men_men_n39_), .Y(men_men_n363_));
  XO2        u341(.A(men_men_n363_), .B(men_men_n243_), .Y(men05));
  NO2        u342(.A(men_men_n301_), .B(men_men_n25_), .Y(men_men_n365_));
  NA3        u343(.A(men_men_n141_), .B(men_men_n131_), .C(men_men_n31_), .Y(men_men_n366_));
  AOI210     u344(.A0(men_men_n226_), .A1(men_men_n53_), .B0(men_men_n87_), .Y(men_men_n367_));
  AOI210     u345(.A0(men_men_n367_), .A1(men_men_n366_), .B0(men_men_n24_), .Y(men_men_n368_));
  OAI210     u346(.A0(men_men_n368_), .A1(men_men_n365_), .B0(men_men_n97_), .Y(men_men_n369_));
  NA2        u347(.A(x11), .B(men_men_n31_), .Y(men_men_n370_));
  NA2        u348(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n371_));
  NA2        u349(.A(men_men_n248_), .B(x03), .Y(men_men_n372_));
  OAI220     u350(.A0(men_men_n372_), .A1(men_men_n371_), .B0(men_men_n370_), .B1(men_men_n78_), .Y(men_men_n373_));
  OAI210     u351(.A0(men_men_n26_), .A1(men_men_n97_), .B0(x07), .Y(men_men_n374_));
  AOI210     u352(.A0(men_men_n373_), .A1(x06), .B0(men_men_n374_), .Y(men_men_n375_));
  AOI220     u353(.A0(men_men_n78_), .A1(men_men_n31_), .B0(men_men_n51_), .B1(men_men_n50_), .Y(men_men_n376_));
  NO3        u354(.A(men_men_n376_), .B(men_men_n23_), .C(x00), .Y(men_men_n377_));
  NA2        u355(.A(men_men_n67_), .B(x02), .Y(men_men_n378_));
  AOI210     u356(.A0(men_men_n378_), .A1(men_men_n372_), .B0(men_men_n251_), .Y(men_men_n379_));
  OR2        u357(.A(men_men_n379_), .B(men_men_n234_), .Y(men_men_n380_));
  NO2        u358(.A(men_men_n23_), .B(x10), .Y(men_men_n381_));
  OAI210     u359(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n382_));
  OR3        u360(.A(men_men_n382_), .B(men_men_n381_), .C(men_men_n44_), .Y(men_men_n383_));
  NA2        u361(.A(men_men_n383_), .B(men_men_n380_), .Y(men_men_n384_));
  OAI210     u362(.A0(men_men_n384_), .A1(men_men_n377_), .B0(men_men_n97_), .Y(men_men_n385_));
  NA2        u363(.A(men_men_n33_), .B(men_men_n97_), .Y(men_men_n386_));
  AOI210     u364(.A0(men_men_n386_), .A1(men_men_n89_), .B0(x07), .Y(men_men_n387_));
  AOI220     u365(.A0(men_men_n387_), .A1(men_men_n385_), .B0(men_men_n375_), .B1(men_men_n369_), .Y(men_men_n388_));
  NA3        u366(.A(men_men_n23_), .B(men_men_n57_), .C(men_men_n48_), .Y(men_men_n389_));
  AO210      u367(.A0(men_men_n389_), .A1(men_men_n261_), .B0(men_men_n258_), .Y(men_men_n390_));
  AOI210     u368(.A0(men_men_n381_), .A1(men_men_n72_), .B0(men_men_n140_), .Y(men_men_n391_));
  OR2        u369(.A(men_men_n391_), .B(x03), .Y(men_men_n392_));
  NO2        u370(.A(x07), .B(x11), .Y(men_men_n393_));
  NO3        u371(.A(men_men_n393_), .B(men_men_n144_), .C(men_men_n28_), .Y(men_men_n394_));
  AOI220     u372(.A0(men_men_n394_), .A1(men_men_n392_), .B0(men_men_n390_), .B1(men_men_n47_), .Y(men_men_n395_));
  NO3        u373(.A(men_men_n321_), .B(men_men_n32_), .C(x11), .Y(men_men_n396_));
  OAI210     u374(.A0(men_men_n396_), .A1(men_men_n395_), .B0(men_men_n98_), .Y(men_men_n397_));
  AOI210     u375(.A0(men_men_n330_), .A1(men_men_n109_), .B0(men_men_n257_), .Y(men_men_n398_));
  NOi21      u376(.An(men_men_n311_), .B(men_men_n133_), .Y(men_men_n399_));
  NO2        u377(.A(men_men_n399_), .B(men_men_n258_), .Y(men_men_n400_));
  OAI210     u378(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n401_));
  AOI210     u379(.A0(men_men_n243_), .A1(men_men_n47_), .B0(men_men_n401_), .Y(men_men_n402_));
  NO4        u380(.A(men_men_n402_), .B(men_men_n400_), .C(men_men_n398_), .D(x08), .Y(men_men_n403_));
  NO2        u381(.A(men_men_n381_), .B(men_men_n31_), .Y(men_men_n404_));
  NA2        u382(.A(x09), .B(men_men_n41_), .Y(men_men_n405_));
  OAI220     u383(.A0(men_men_n405_), .A1(men_men_n404_), .B0(men_men_n370_), .B1(men_men_n63_), .Y(men_men_n406_));
  NO2        u384(.A(x13), .B(x12), .Y(men_men_n407_));
  NO2        u385(.A(men_men_n131_), .B(men_men_n28_), .Y(men_men_n408_));
  NO2        u386(.A(men_men_n408_), .B(men_men_n262_), .Y(men_men_n409_));
  OR3        u387(.A(men_men_n409_), .B(x12), .C(x03), .Y(men_men_n410_));
  NA3        u388(.A(men_men_n324_), .B(men_men_n124_), .C(x12), .Y(men_men_n411_));
  AO210      u389(.A0(men_men_n324_), .A1(men_men_n124_), .B0(men_men_n243_), .Y(men_men_n412_));
  NA4        u390(.A(men_men_n412_), .B(men_men_n411_), .C(men_men_n410_), .D(x08), .Y(men_men_n413_));
  AOI210     u391(.A0(men_men_n407_), .A1(men_men_n406_), .B0(men_men_n413_), .Y(men_men_n414_));
  AOI210     u392(.A0(men_men_n403_), .A1(men_men_n397_), .B0(men_men_n414_), .Y(men_men_n415_));
  OAI210     u393(.A0(x07), .A1(men_men_n23_), .B0(x03), .Y(men_men_n416_));
  NO2        u394(.A(men_men_n437_), .B(men_men_n371_), .Y(men_men_n417_));
  OAI210     u395(.A0(men_men_n417_), .A1(men_men_n416_), .B0(men_men_n182_), .Y(men_men_n418_));
  NA3        u396(.A(men_men_n409_), .B(men_men_n399_), .C(men_men_n320_), .Y(men_men_n419_));
  INV        u397(.A(x14), .Y(men_men_n420_));
  NO3        u398(.A(men_men_n311_), .B(men_men_n104_), .C(x11), .Y(men_men_n421_));
  NO3        u399(.A(men_men_n164_), .B(men_men_n72_), .C(men_men_n53_), .Y(men_men_n422_));
  NO3        u400(.A(men_men_n389_), .B(men_men_n321_), .C(men_men_n177_), .Y(men_men_n423_));
  NO4        u401(.A(men_men_n423_), .B(men_men_n422_), .C(men_men_n421_), .D(men_men_n420_), .Y(men_men_n424_));
  NA3        u402(.A(men_men_n424_), .B(men_men_n419_), .C(men_men_n418_), .Y(men_men_n425_));
  AOI220     u403(.A0(men_men_n386_), .A1(men_men_n57_), .B0(men_men_n408_), .B1(men_men_n163_), .Y(men_men_n426_));
  NOi21      u404(.An(men_men_n265_), .B(men_men_n148_), .Y(men_men_n427_));
  NO3        u405(.A(men_men_n128_), .B(men_men_n24_), .C(x06), .Y(men_men_n428_));
  AOI210     u406(.A0(men_men_n272_), .A1(men_men_n226_), .B0(men_men_n428_), .Y(men_men_n429_));
  OAI210     u407(.A0(men_men_n44_), .A1(x04), .B0(men_men_n429_), .Y(men_men_n430_));
  OAI210     u408(.A0(men_men_n430_), .A1(men_men_n427_), .B0(men_men_n97_), .Y(men_men_n431_));
  OAI210     u409(.A0(men_men_n426_), .A1(men_men_n88_), .B0(men_men_n431_), .Y(men_men_n432_));
  NO4        u410(.A(men_men_n432_), .B(men_men_n425_), .C(men_men_n415_), .D(men_men_n388_), .Y(men06));
  INV        u411(.A(x07), .Y(men_men_n436_));
  INV        u412(.A(x07), .Y(men_men_n437_));
  INV        u413(.A(men_men_n90_), .Y(men_men_n438_));
  INV        u414(.A(x01), .Y(men_men_n439_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule