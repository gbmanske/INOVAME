// Benchmark "top" written by ABC on Fri Jun 21 17:49:22 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n139_,
    new_new_n140_, new_new_n141_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1071_,
    new_new_n1072_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(mai1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  NO2        g0037(.A(new_new_n59_), .B(new_new_n58_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n51_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g0062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g0063(.A(i_6_), .Y(new_new_n86_));
  OR4        g0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g0065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g0066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  NO2        g0067(.A(new_new_n88_), .B(new_new_n89_), .Y(new_new_n90_));
  OAI210     g0068(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n90_), .Y(new_new_n91_));
  NAi21      g0069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g0070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g0071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n63_), .Y(new_new_n94_));
  NA2        g0072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  INV        g0073(.A(new_new_n94_), .Y(new_new_n96_));
  AOI210     g0074(.A0(new_new_n96_), .A1(new_new_n91_), .B0(new_new_n80_), .Y(new_new_n97_));
  AN3        g0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n98_));
  NAi21      g0076(.An(i_6_), .B(i_11_), .Y(new_new_n99_));
  NO2        g0077(.A(i_5_), .B(i_8_), .Y(new_new_n100_));
  NOi21      g0078(.An(new_new_n100_), .B(new_new_n99_), .Y(new_new_n101_));
  AOI220     g0079(.A0(new_new_n101_), .A1(new_new_n62_), .B0(new_new_n98_), .B1(new_new_n32_), .Y(new_new_n102_));
  INV        g0080(.A(i_7_), .Y(new_new_n103_));
  NA2        g0081(.A(new_new_n47_), .B(new_new_n103_), .Y(new_new_n104_));
  NO2        g0082(.A(i_0_), .B(i_5_), .Y(new_new_n105_));
  NO2        g0083(.A(new_new_n105_), .B(new_new_n86_), .Y(new_new_n106_));
  NA2        g0084(.A(i_12_), .B(i_3_), .Y(new_new_n107_));
  INV        g0085(.A(new_new_n107_), .Y(new_new_n108_));
  NA3        g0086(.A(new_new_n108_), .B(new_new_n106_), .C(new_new_n104_), .Y(new_new_n109_));
  NAi21      g0087(.An(i_7_), .B(i_11_), .Y(new_new_n110_));
  AN2        g0088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g0089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g0090(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n113_));
  NO2        g0091(.A(i_8_), .B(new_new_n103_), .Y(new_new_n114_));
  NO3        g0092(.A(new_new_n114_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n115_));
  NA2        g0093(.A(i_12_), .B(i_7_), .Y(new_new_n116_));
  NO2        g0094(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n117_));
  NA2        g0095(.A(i_11_), .B(i_12_), .Y(new_new_n118_));
  INV        g0096(.A(new_new_n118_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n119_), .B(new_new_n115_), .Y(new_new_n120_));
  NA3        g0098(.A(new_new_n120_), .B(new_new_n109_), .C(new_new_n102_), .Y(new_new_n121_));
  NOi21      g0099(.An(i_1_), .B(i_5_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(i_11_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n124_));
  NA2        g0102(.A(i_7_), .B(new_new_n25_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n125_), .B(new_new_n124_), .Y(new_new_n126_));
  NO2        g0104(.A(new_new_n126_), .B(new_new_n47_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n128_));
  NAi21      g0106(.An(i_3_), .B(i_8_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n129_), .B(new_new_n62_), .Y(new_new_n130_));
  NOi31      g0108(.An(new_new_n130_), .B(new_new_n128_), .C(new_new_n127_), .Y(new_new_n131_));
  NO2        g0109(.A(i_1_), .B(new_new_n86_), .Y(new_new_n132_));
  NO2        g0110(.A(i_6_), .B(i_5_), .Y(new_new_n133_));
  NA2        g0111(.A(new_new_n133_), .B(i_3_), .Y(new_new_n134_));
  AO210      g0112(.A0(new_new_n134_), .A1(new_new_n48_), .B0(new_new_n132_), .Y(new_new_n135_));
  OAI220     g0113(.A0(new_new_n135_), .A1(new_new_n110_), .B0(new_new_n131_), .B1(new_new_n123_), .Y(new_new_n136_));
  NO3        g0114(.A(new_new_n136_), .B(new_new_n121_), .C(new_new_n97_), .Y(new_new_n137_));
  NA3        g0115(.A(new_new_n137_), .B(new_new_n79_), .C(new_new_n57_), .Y(mai2));
  NO2        g0116(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n139_));
  NA2        g0117(.A(i_6_), .B(new_new_n25_), .Y(new_new_n140_));
  NA2        g0118(.A(new_new_n140_), .B(new_new_n139_), .Y(new_new_n141_));
  NA4        g0119(.A(new_new_n141_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(mai0));
  AN2        g0120(.A(i_8_), .B(i_7_), .Y(new_new_n143_));
  NA2        g0121(.A(new_new_n143_), .B(i_6_), .Y(new_new_n144_));
  NO2        g0122(.A(i_12_), .B(i_13_), .Y(new_new_n145_));
  NAi21      g0123(.An(i_5_), .B(i_11_), .Y(new_new_n146_));
  NOi21      g0124(.An(new_new_n145_), .B(new_new_n146_), .Y(new_new_n147_));
  NO2        g0125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NA2        g0126(.A(i_2_), .B(i_3_), .Y(new_new_n149_));
  NO2        g0127(.A(new_new_n149_), .B(i_4_), .Y(new_new_n150_));
  NA3        g0128(.A(new_new_n150_), .B(new_new_n148_), .C(new_new_n147_), .Y(new_new_n151_));
  AN2        g0129(.A(new_new_n145_), .B(new_new_n83_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n152_), .B(new_new_n27_), .Y(new_new_n153_));
  NA2        g0131(.A(i_1_), .B(i_5_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n73_), .B(new_new_n47_), .Y(new_new_n155_));
  NA2        g0133(.A(new_new_n155_), .B(new_new_n36_), .Y(new_new_n156_));
  NO3        g0134(.A(new_new_n156_), .B(new_new_n154_), .C(new_new_n153_), .Y(new_new_n157_));
  OR2        g0135(.A(i_0_), .B(i_1_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n159_));
  NAi32      g0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n160_));
  NAi21      g0138(.An(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  NOi21      g0139(.An(i_4_), .B(i_10_), .Y(new_new_n162_));
  NA2        g0140(.A(new_new_n162_), .B(new_new_n40_), .Y(new_new_n163_));
  NO2        g0141(.A(i_3_), .B(i_5_), .Y(new_new_n164_));
  NO3        g0142(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n165_));
  NA2        g0143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OAI210     g0144(.A0(new_new_n166_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n167_));
  NO2        g0145(.A(new_new_n167_), .B(new_new_n157_), .Y(new_new_n168_));
  AOI210     g0146(.A0(new_new_n168_), .A1(new_new_n151_), .B0(new_new_n144_), .Y(new_new_n169_));
  NA3        g0147(.A(new_new_n73_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n170_));
  NA2        g0148(.A(i_3_), .B(new_new_n49_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_4_), .B(i_9_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_11_), .B(i_13_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n173_), .B(new_new_n172_), .Y(new_new_n174_));
  OR2        g0152(.A(new_new_n174_), .B(new_new_n171_), .Y(new_new_n175_));
  NO2        g0153(.A(i_4_), .B(i_5_), .Y(new_new_n176_));
  NAi21      g0154(.An(i_12_), .B(i_11_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n177_), .B(i_13_), .Y(new_new_n178_));
  NA3        g0156(.A(new_new_n178_), .B(new_new_n176_), .C(new_new_n83_), .Y(new_new_n179_));
  AOI210     g0157(.A0(new_new_n179_), .A1(new_new_n175_), .B0(new_new_n170_), .Y(new_new_n180_));
  NO2        g0158(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n181_), .B(new_new_n47_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n36_), .B(i_5_), .Y(new_new_n183_));
  NAi31      g0161(.An(new_new_n183_), .B(new_new_n152_), .C(i_11_), .Y(new_new_n184_));
  NA2        g0162(.A(i_3_), .B(i_5_), .Y(new_new_n185_));
  OR2        g0163(.A(new_new_n185_), .B(new_new_n174_), .Y(new_new_n186_));
  AOI210     g0164(.A0(new_new_n186_), .A1(new_new_n184_), .B0(new_new_n182_), .Y(new_new_n187_));
  NO2        g0165(.A(new_new_n73_), .B(i_5_), .Y(new_new_n188_));
  NO2        g0166(.A(i_13_), .B(i_10_), .Y(new_new_n189_));
  NA3        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n45_), .Y(new_new_n190_));
  NO2        g0168(.A(i_2_), .B(i_1_), .Y(new_new_n191_));
  NA2        g0169(.A(new_new_n191_), .B(i_3_), .Y(new_new_n192_));
  NAi21      g0170(.An(i_4_), .B(i_12_), .Y(new_new_n193_));
  NO4        g0171(.A(new_new_n193_), .B(new_new_n192_), .C(new_new_n190_), .D(new_new_n25_), .Y(new_new_n194_));
  NO3        g0172(.A(new_new_n194_), .B(new_new_n187_), .C(new_new_n180_), .Y(new_new_n195_));
  INV        g0173(.A(i_8_), .Y(new_new_n196_));
  NO2        g0174(.A(new_new_n196_), .B(i_7_), .Y(new_new_n197_));
  NA2        g0175(.A(new_new_n197_), .B(i_6_), .Y(new_new_n198_));
  NO3        g0176(.A(i_3_), .B(new_new_n86_), .C(new_new_n49_), .Y(new_new_n199_));
  NA2        g0177(.A(new_new_n199_), .B(new_new_n114_), .Y(new_new_n200_));
  NO3        g0178(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n201_));
  NA3        g0179(.A(new_new_n201_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n202_));
  NO3        g0180(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n203_));
  OAI210     g0181(.A0(new_new_n98_), .A1(i_12_), .B0(new_new_n203_), .Y(new_new_n204_));
  AOI210     g0182(.A0(new_new_n204_), .A1(new_new_n202_), .B0(new_new_n200_), .Y(new_new_n205_));
  NO2        g0183(.A(i_3_), .B(i_8_), .Y(new_new_n206_));
  NO3        g0184(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n207_));
  NO2        g0185(.A(new_new_n105_), .B(new_new_n58_), .Y(new_new_n208_));
  NO2        g0186(.A(i_13_), .B(i_9_), .Y(new_new_n209_));
  NA3        g0187(.A(new_new_n209_), .B(i_6_), .C(new_new_n196_), .Y(new_new_n210_));
  NAi21      g0188(.An(i_12_), .B(i_3_), .Y(new_new_n211_));
  NO2        g0189(.A(new_new_n45_), .B(i_5_), .Y(new_new_n212_));
  NO3        g0190(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n213_));
  NA3        g0191(.A(new_new_n213_), .B(new_new_n212_), .C(i_10_), .Y(new_new_n214_));
  NO2        g0192(.A(new_new_n214_), .B(new_new_n210_), .Y(new_new_n215_));
  AOI210     g0193(.A0(new_new_n215_), .A1(i_7_), .B0(new_new_n205_), .Y(new_new_n216_));
  OAI220     g0194(.A0(new_new_n216_), .A1(i_4_), .B0(new_new_n198_), .B1(new_new_n195_), .Y(new_new_n217_));
  NAi21      g0195(.An(i_12_), .B(i_7_), .Y(new_new_n218_));
  NA3        g0196(.A(i_13_), .B(new_new_n196_), .C(i_10_), .Y(new_new_n219_));
  NO2        g0197(.A(new_new_n219_), .B(new_new_n218_), .Y(new_new_n220_));
  NA2        g0198(.A(i_0_), .B(i_5_), .Y(new_new_n221_));
  NA2        g0199(.A(new_new_n221_), .B(new_new_n106_), .Y(new_new_n222_));
  OAI220     g0200(.A0(new_new_n222_), .A1(new_new_n192_), .B0(new_new_n182_), .B1(new_new_n134_), .Y(new_new_n223_));
  NAi31      g0201(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n36_), .B(i_13_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n226_));
  NO2        g0204(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n227_));
  NA3        g0205(.A(new_new_n227_), .B(new_new_n226_), .C(new_new_n225_), .Y(new_new_n228_));
  INV        g0206(.A(i_13_), .Y(new_new_n229_));
  NO2        g0207(.A(i_12_), .B(new_new_n229_), .Y(new_new_n230_));
  NA3        g0208(.A(new_new_n230_), .B(new_new_n201_), .C(new_new_n199_), .Y(new_new_n231_));
  OAI210     g0209(.A0(new_new_n228_), .A1(new_new_n224_), .B0(new_new_n231_), .Y(new_new_n232_));
  AOI220     g0210(.A0(new_new_n232_), .A1(new_new_n143_), .B0(new_new_n223_), .B1(new_new_n220_), .Y(new_new_n233_));
  NO2        g0211(.A(i_12_), .B(new_new_n37_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n185_), .B(i_4_), .Y(new_new_n235_));
  NA2        g0213(.A(new_new_n235_), .B(new_new_n234_), .Y(new_new_n236_));
  OR2        g0214(.A(i_8_), .B(i_7_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n237_), .B(new_new_n86_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n54_), .B(i_1_), .Y(new_new_n239_));
  NA2        g0217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  INV        g0218(.A(i_12_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n45_), .B(new_new_n241_), .Y(new_new_n242_));
  NO3        g0220(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n243_));
  NA2        g0221(.A(i_2_), .B(i_1_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n240_), .B(new_new_n236_), .Y(new_new_n245_));
  NO3        g0223(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n246_));
  NAi21      g0224(.An(i_4_), .B(i_3_), .Y(new_new_n247_));
  NO2        g0225(.A(new_new_n247_), .B(new_new_n75_), .Y(new_new_n248_));
  NO2        g0226(.A(i_0_), .B(i_6_), .Y(new_new_n249_));
  NOi41      g0227(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n250_));
  NA2        g0228(.A(new_new_n250_), .B(new_new_n249_), .Y(new_new_n251_));
  NO2        g0229(.A(new_new_n244_), .B(new_new_n185_), .Y(new_new_n252_));
  NAi21      g0230(.An(new_new_n251_), .B(new_new_n252_), .Y(new_new_n253_));
  INV        g0231(.A(new_new_n253_), .Y(new_new_n254_));
  AOI210     g0232(.A0(new_new_n254_), .A1(new_new_n40_), .B0(new_new_n245_), .Y(new_new_n255_));
  NO2        g0233(.A(i_11_), .B(new_new_n229_), .Y(new_new_n256_));
  NOi21      g0234(.An(i_1_), .B(i_6_), .Y(new_new_n257_));
  NAi21      g0235(.An(i_3_), .B(i_7_), .Y(new_new_n258_));
  NA2        g0236(.A(new_new_n241_), .B(i_9_), .Y(new_new_n259_));
  OR4        g0237(.A(new_new_n259_), .B(new_new_n258_), .C(new_new_n257_), .D(new_new_n188_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n261_));
  NO2        g0239(.A(i_12_), .B(i_3_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n73_), .B(i_5_), .Y(new_new_n263_));
  NA2        g0241(.A(i_3_), .B(i_9_), .Y(new_new_n264_));
  NAi21      g0242(.An(i_7_), .B(i_10_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n266_));
  NA3        g0244(.A(new_new_n266_), .B(new_new_n263_), .C(new_new_n64_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n267_), .B(new_new_n260_), .Y(new_new_n268_));
  NA3        g0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n269_));
  INV        g0247(.A(new_new_n144_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n241_), .B(i_13_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n271_), .B(new_new_n75_), .Y(new_new_n272_));
  AOI220     g0250(.A0(new_new_n272_), .A1(new_new_n270_), .B0(new_new_n268_), .B1(new_new_n256_), .Y(new_new_n273_));
  NO2        g0251(.A(new_new_n237_), .B(new_new_n37_), .Y(new_new_n274_));
  NA2        g0252(.A(i_12_), .B(i_6_), .Y(new_new_n275_));
  OR2        g0253(.A(i_13_), .B(i_9_), .Y(new_new_n276_));
  NO2        g0254(.A(new_new_n247_), .B(i_2_), .Y(new_new_n277_));
  NA2        g0255(.A(new_new_n256_), .B(i_9_), .Y(new_new_n278_));
  NA2        g0256(.A(new_new_n155_), .B(new_new_n63_), .Y(new_new_n279_));
  NO3        g0257(.A(i_11_), .B(new_new_n229_), .C(new_new_n25_), .Y(new_new_n280_));
  NO2        g0258(.A(new_new_n258_), .B(i_8_), .Y(new_new_n281_));
  NO2        g0259(.A(i_6_), .B(new_new_n49_), .Y(new_new_n282_));
  NA3        g0260(.A(new_new_n282_), .B(new_new_n281_), .C(new_new_n280_), .Y(new_new_n283_));
  NO3        g0261(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n284_));
  NA3        g0262(.A(new_new_n284_), .B(new_new_n274_), .C(new_new_n230_), .Y(new_new_n285_));
  AOI210     g0263(.A0(new_new_n285_), .A1(new_new_n283_), .B0(new_new_n279_), .Y(new_new_n286_));
  INV        g0264(.A(new_new_n286_), .Y(new_new_n287_));
  NA4        g0265(.A(new_new_n287_), .B(new_new_n273_), .C(new_new_n255_), .D(new_new_n233_), .Y(new_new_n288_));
  NO3        g0266(.A(i_12_), .B(new_new_n229_), .C(new_new_n37_), .Y(new_new_n289_));
  INV        g0267(.A(new_new_n289_), .Y(new_new_n290_));
  NA2        g0268(.A(i_8_), .B(new_new_n103_), .Y(new_new_n291_));
  NOi21      g0269(.An(new_new_n164_), .B(new_new_n86_), .Y(new_new_n292_));
  NO3        g0270(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n293_));
  AOI220     g0271(.A0(new_new_n293_), .A1(new_new_n199_), .B0(new_new_n292_), .B1(new_new_n239_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n294_), .B(new_new_n291_), .Y(new_new_n295_));
  NO3        g0273(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n296_));
  NO2        g0274(.A(new_new_n244_), .B(i_0_), .Y(new_new_n297_));
  AOI220     g0275(.A0(new_new_n297_), .A1(new_new_n197_), .B0(new_new_n296_), .B1(new_new_n143_), .Y(new_new_n298_));
  NA2        g0276(.A(new_new_n282_), .B(new_new_n26_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n299_), .B(new_new_n298_), .Y(new_new_n300_));
  NA2        g0278(.A(i_0_), .B(i_1_), .Y(new_new_n301_));
  NO2        g0279(.A(new_new_n301_), .B(i_2_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n59_), .B(i_6_), .Y(new_new_n303_));
  NA3        g0281(.A(new_new_n303_), .B(new_new_n302_), .C(new_new_n164_), .Y(new_new_n304_));
  OAI210     g0282(.A0(new_new_n166_), .A1(new_new_n144_), .B0(new_new_n304_), .Y(new_new_n305_));
  NO3        g0283(.A(new_new_n305_), .B(new_new_n300_), .C(new_new_n295_), .Y(new_new_n306_));
  NO2        g0284(.A(i_3_), .B(i_10_), .Y(new_new_n307_));
  NA3        g0285(.A(new_new_n307_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n308_));
  NO2        g0286(.A(i_2_), .B(new_new_n103_), .Y(new_new_n309_));
  NA2        g0287(.A(i_1_), .B(new_new_n36_), .Y(new_new_n310_));
  NO2        g0288(.A(new_new_n310_), .B(i_8_), .Y(new_new_n311_));
  NA2        g0289(.A(new_new_n311_), .B(new_new_n309_), .Y(new_new_n312_));
  AN2        g0290(.A(i_3_), .B(i_10_), .Y(new_new_n313_));
  NA4        g0291(.A(new_new_n313_), .B(new_new_n201_), .C(new_new_n178_), .D(new_new_n176_), .Y(new_new_n314_));
  NO2        g0292(.A(i_5_), .B(new_new_n37_), .Y(new_new_n315_));
  NO2        g0293(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n316_));
  OR2        g0294(.A(new_new_n312_), .B(new_new_n308_), .Y(new_new_n317_));
  OAI220     g0295(.A0(new_new_n317_), .A1(i_6_), .B0(new_new_n306_), .B1(new_new_n290_), .Y(new_new_n318_));
  NO4        g0296(.A(new_new_n318_), .B(new_new_n288_), .C(new_new_n217_), .D(new_new_n169_), .Y(new_new_n319_));
  NO3        g0297(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n320_));
  NO2        g0298(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n321_));
  NA2        g0299(.A(new_new_n297_), .B(new_new_n321_), .Y(new_new_n322_));
  NO3        g0300(.A(i_6_), .B(new_new_n196_), .C(i_7_), .Y(new_new_n323_));
  NA2        g0301(.A(new_new_n323_), .B(new_new_n201_), .Y(new_new_n324_));
  AOI210     g0302(.A0(new_new_n324_), .A1(new_new_n322_), .B0(new_new_n171_), .Y(new_new_n325_));
  NO2        g0303(.A(i_2_), .B(i_3_), .Y(new_new_n326_));
  OR2        g0304(.A(i_0_), .B(i_5_), .Y(new_new_n327_));
  NA2        g0305(.A(new_new_n221_), .B(new_new_n327_), .Y(new_new_n328_));
  NA4        g0306(.A(new_new_n328_), .B(new_new_n238_), .C(new_new_n326_), .D(i_1_), .Y(new_new_n329_));
  NA3        g0307(.A(new_new_n297_), .B(new_new_n292_), .C(new_new_n114_), .Y(new_new_n330_));
  NAi21      g0308(.An(i_8_), .B(i_7_), .Y(new_new_n331_));
  NO2        g0309(.A(new_new_n331_), .B(i_6_), .Y(new_new_n332_));
  NO2        g0310(.A(new_new_n158_), .B(new_new_n47_), .Y(new_new_n333_));
  NA3        g0311(.A(new_new_n333_), .B(new_new_n332_), .C(new_new_n164_), .Y(new_new_n334_));
  NA3        g0312(.A(new_new_n334_), .B(new_new_n330_), .C(new_new_n329_), .Y(new_new_n335_));
  OAI210     g0313(.A0(new_new_n335_), .A1(new_new_n325_), .B0(i_4_), .Y(new_new_n336_));
  NO2        g0314(.A(i_12_), .B(i_10_), .Y(new_new_n337_));
  NOi21      g0315(.An(i_5_), .B(i_0_), .Y(new_new_n338_));
  NO3        g0316(.A(new_new_n310_), .B(new_new_n338_), .C(new_new_n129_), .Y(new_new_n339_));
  NA4        g0317(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n340_));
  NA2        g0318(.A(new_new_n339_), .B(new_new_n337_), .Y(new_new_n341_));
  NO2        g0319(.A(i_6_), .B(i_8_), .Y(new_new_n342_));
  NOi21      g0320(.An(i_0_), .B(i_2_), .Y(new_new_n343_));
  AN2        g0321(.A(new_new_n343_), .B(new_new_n342_), .Y(new_new_n344_));
  NO2        g0322(.A(i_1_), .B(i_7_), .Y(new_new_n345_));
  AO220      g0323(.A0(new_new_n345_), .A1(new_new_n344_), .B0(new_new_n332_), .B1(new_new_n239_), .Y(new_new_n346_));
  NA3        g0324(.A(new_new_n346_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n347_));
  NA3        g0325(.A(new_new_n347_), .B(new_new_n341_), .C(new_new_n336_), .Y(new_new_n348_));
  NO3        g0326(.A(new_new_n237_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n349_));
  NO3        g0327(.A(new_new_n331_), .B(i_2_), .C(i_1_), .Y(new_new_n350_));
  OAI210     g0328(.A0(new_new_n350_), .A1(new_new_n349_), .B0(i_6_), .Y(new_new_n351_));
  NA3        g0329(.A(new_new_n257_), .B(new_new_n309_), .C(new_new_n196_), .Y(new_new_n352_));
  AOI210     g0330(.A0(new_new_n352_), .A1(new_new_n351_), .B0(new_new_n328_), .Y(new_new_n353_));
  INV        g0331(.A(new_new_n106_), .Y(new_new_n354_));
  NA2        g0332(.A(new_new_n353_), .B(i_3_), .Y(new_new_n355_));
  INV        g0333(.A(new_new_n84_), .Y(new_new_n356_));
  NO2        g0334(.A(new_new_n301_), .B(new_new_n81_), .Y(new_new_n357_));
  NA2        g0335(.A(new_new_n357_), .B(new_new_n133_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n95_), .B(new_new_n196_), .Y(new_new_n359_));
  NA2        g0337(.A(new_new_n359_), .B(new_new_n63_), .Y(new_new_n360_));
  AOI210     g0338(.A0(new_new_n360_), .A1(new_new_n358_), .B0(new_new_n356_), .Y(new_new_n361_));
  NO2        g0339(.A(new_new_n196_), .B(i_9_), .Y(new_new_n362_));
  NA2        g0340(.A(new_new_n362_), .B(new_new_n208_), .Y(new_new_n363_));
  NO2        g0341(.A(new_new_n361_), .B(new_new_n300_), .Y(new_new_n364_));
  AOI210     g0342(.A0(new_new_n364_), .A1(new_new_n355_), .B0(new_new_n163_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n348_), .A1(new_new_n320_), .B0(new_new_n365_), .Y(new_new_n366_));
  NOi32      g0344(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n367_));
  INV        g0345(.A(new_new_n367_), .Y(new_new_n368_));
  NAi21      g0346(.An(i_0_), .B(i_6_), .Y(new_new_n369_));
  NAi21      g0347(.An(i_1_), .B(i_5_), .Y(new_new_n370_));
  NA2        g0348(.A(new_new_n370_), .B(new_new_n369_), .Y(new_new_n371_));
  NA2        g0349(.A(new_new_n371_), .B(new_new_n25_), .Y(new_new_n372_));
  OAI210     g0350(.A0(new_new_n372_), .A1(new_new_n160_), .B0(new_new_n251_), .Y(new_new_n373_));
  NAi41      g0351(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n374_));
  OAI220     g0352(.A0(new_new_n374_), .A1(new_new_n370_), .B0(new_new_n224_), .B1(new_new_n160_), .Y(new_new_n375_));
  AOI210     g0353(.A0(new_new_n374_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n376_));
  NOi32      g0354(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n377_));
  OR2        g0355(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n378_));
  NO2        g0356(.A(i_1_), .B(new_new_n103_), .Y(new_new_n379_));
  NAi21      g0357(.An(i_3_), .B(i_4_), .Y(new_new_n380_));
  NO2        g0358(.A(new_new_n380_), .B(i_9_), .Y(new_new_n381_));
  AN2        g0359(.A(i_6_), .B(i_7_), .Y(new_new_n382_));
  OAI210     g0360(.A0(new_new_n382_), .A1(new_new_n379_), .B0(new_new_n381_), .Y(new_new_n383_));
  NA2        g0361(.A(i_2_), .B(i_7_), .Y(new_new_n384_));
  NO2        g0362(.A(new_new_n380_), .B(i_10_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n383_), .B(new_new_n188_), .Y(new_new_n386_));
  AOI210     g0364(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n387_));
  OAI210     g0365(.A0(new_new_n387_), .A1(new_new_n191_), .B0(new_new_n385_), .Y(new_new_n388_));
  AOI220     g0366(.A0(new_new_n385_), .A1(new_new_n345_), .B0(new_new_n243_), .B1(new_new_n191_), .Y(new_new_n389_));
  AOI210     g0367(.A0(new_new_n389_), .A1(new_new_n388_), .B0(i_5_), .Y(new_new_n390_));
  NO4        g0368(.A(new_new_n390_), .B(new_new_n386_), .C(new_new_n378_), .D(new_new_n373_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n391_), .B(new_new_n368_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n393_));
  AN2        g0371(.A(i_12_), .B(i_5_), .Y(new_new_n394_));
  NO2        g0372(.A(i_4_), .B(new_new_n26_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n395_), .B(new_new_n394_), .Y(new_new_n396_));
  NO2        g0374(.A(i_11_), .B(i_6_), .Y(new_new_n397_));
  NA3        g0375(.A(new_new_n397_), .B(new_new_n333_), .C(new_new_n229_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n398_), .B(new_new_n396_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n247_), .B(i_5_), .Y(new_new_n400_));
  NO2        g0378(.A(i_5_), .B(i_10_), .Y(new_new_n401_));
  AOI220     g0379(.A0(new_new_n401_), .A1(new_new_n277_), .B0(new_new_n400_), .B1(new_new_n201_), .Y(new_new_n402_));
  NA2        g0380(.A(new_new_n145_), .B(new_new_n46_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n403_), .B(new_new_n402_), .Y(new_new_n404_));
  OAI210     g0382(.A0(new_new_n404_), .A1(new_new_n399_), .B0(new_new_n393_), .Y(new_new_n405_));
  NO2        g0383(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n406_));
  NO2        g0384(.A(new_new_n151_), .B(new_new_n86_), .Y(new_new_n407_));
  OAI210     g0385(.A0(new_new_n407_), .A1(new_new_n399_), .B0(new_new_n406_), .Y(new_new_n408_));
  NO3        g0386(.A(new_new_n86_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n409_));
  NO2        g0387(.A(i_3_), .B(new_new_n103_), .Y(new_new_n410_));
  NA3        g0388(.A(new_new_n307_), .B(new_new_n93_), .C(new_new_n55_), .Y(new_new_n411_));
  NO2        g0389(.A(i_11_), .B(i_12_), .Y(new_new_n412_));
  NA2        g0390(.A(new_new_n412_), .B(new_new_n36_), .Y(new_new_n413_));
  NO2        g0391(.A(new_new_n411_), .B(new_new_n413_), .Y(new_new_n414_));
  NA2        g0392(.A(new_new_n401_), .B(new_new_n241_), .Y(new_new_n415_));
  NA3        g0393(.A(new_new_n114_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n416_), .B(new_new_n224_), .Y(new_new_n417_));
  NAi21      g0395(.An(i_13_), .B(i_0_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n418_), .B(new_new_n244_), .Y(new_new_n419_));
  OAI210     g0397(.A0(new_new_n417_), .A1(new_new_n414_), .B0(new_new_n419_), .Y(new_new_n420_));
  NA3        g0398(.A(new_new_n420_), .B(new_new_n408_), .C(new_new_n405_), .Y(new_new_n421_));
  NA2        g0399(.A(new_new_n45_), .B(new_new_n229_), .Y(new_new_n422_));
  NO3        g0400(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n423_));
  NO2        g0401(.A(i_0_), .B(i_11_), .Y(new_new_n424_));
  INV        g0402(.A(i_5_), .Y(new_new_n425_));
  AN2        g0403(.A(i_1_), .B(i_6_), .Y(new_new_n426_));
  NOi21      g0404(.An(i_2_), .B(i_12_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n427_), .B(new_new_n426_), .Y(new_new_n428_));
  NO2        g0406(.A(new_new_n428_), .B(new_new_n425_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n143_), .B(i_9_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n430_), .B(i_4_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n429_), .B(new_new_n431_), .Y(new_new_n432_));
  NAi21      g0410(.An(i_9_), .B(i_4_), .Y(new_new_n433_));
  OR2        g0411(.A(i_13_), .B(i_10_), .Y(new_new_n434_));
  NO3        g0412(.A(new_new_n434_), .B(new_new_n118_), .C(new_new_n433_), .Y(new_new_n435_));
  OR2        g0413(.A(new_new_n219_), .B(new_new_n218_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n103_), .B(new_new_n25_), .Y(new_new_n437_));
  NA2        g0415(.A(new_new_n289_), .B(new_new_n437_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n282_), .B(new_new_n213_), .Y(new_new_n439_));
  OAI220     g0417(.A0(new_new_n439_), .A1(new_new_n436_), .B0(new_new_n438_), .B1(new_new_n354_), .Y(new_new_n440_));
  INV        g0418(.A(new_new_n440_), .Y(new_new_n441_));
  AOI210     g0419(.A0(new_new_n441_), .A1(new_new_n432_), .B0(new_new_n26_), .Y(new_new_n442_));
  NA2        g0420(.A(new_new_n330_), .B(new_new_n329_), .Y(new_new_n443_));
  AOI220     g0421(.A0(new_new_n303_), .A1(new_new_n293_), .B0(new_new_n297_), .B1(new_new_n321_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n444_), .B(new_new_n171_), .Y(new_new_n445_));
  NO2        g0423(.A(new_new_n185_), .B(new_new_n86_), .Y(new_new_n446_));
  AOI220     g0424(.A0(new_new_n446_), .A1(new_new_n302_), .B0(new_new_n284_), .B1(new_new_n213_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n447_), .B(new_new_n291_), .Y(new_new_n448_));
  NO3        g0426(.A(new_new_n448_), .B(new_new_n445_), .C(new_new_n443_), .Y(new_new_n449_));
  NA2        g0427(.A(new_new_n199_), .B(new_new_n98_), .Y(new_new_n450_));
  NA3        g0428(.A(new_new_n333_), .B(new_new_n164_), .C(new_new_n86_), .Y(new_new_n451_));
  AOI210     g0429(.A0(new_new_n451_), .A1(new_new_n450_), .B0(new_new_n331_), .Y(new_new_n452_));
  NA2        g0430(.A(new_new_n196_), .B(i_10_), .Y(new_new_n453_));
  NA3        g0431(.A(new_new_n263_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n454_));
  NA2        g0432(.A(new_new_n303_), .B(new_new_n239_), .Y(new_new_n455_));
  OAI220     g0433(.A0(new_new_n455_), .A1(new_new_n185_), .B0(new_new_n454_), .B1(new_new_n453_), .Y(new_new_n456_));
  NO2        g0434(.A(i_3_), .B(new_new_n49_), .Y(new_new_n457_));
  NA3        g0435(.A(new_new_n345_), .B(new_new_n344_), .C(new_new_n457_), .Y(new_new_n458_));
  NA2        g0436(.A(new_new_n323_), .B(new_new_n328_), .Y(new_new_n459_));
  OAI210     g0437(.A0(new_new_n459_), .A1(new_new_n192_), .B0(new_new_n458_), .Y(new_new_n460_));
  NO3        g0438(.A(new_new_n460_), .B(new_new_n456_), .C(new_new_n452_), .Y(new_new_n461_));
  AOI210     g0439(.A0(new_new_n461_), .A1(new_new_n449_), .B0(new_new_n278_), .Y(new_new_n462_));
  NO4        g0440(.A(new_new_n462_), .B(new_new_n442_), .C(new_new_n421_), .D(new_new_n392_), .Y(new_new_n463_));
  NO2        g0441(.A(new_new_n63_), .B(i_4_), .Y(new_new_n464_));
  NO2        g0442(.A(new_new_n73_), .B(i_13_), .Y(new_new_n465_));
  NO2        g0443(.A(i_10_), .B(i_9_), .Y(new_new_n466_));
  NAi21      g0444(.An(i_12_), .B(i_8_), .Y(new_new_n467_));
  NO2        g0445(.A(new_new_n467_), .B(i_3_), .Y(new_new_n468_));
  NO2        g0446(.A(new_new_n47_), .B(i_4_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n316_), .B(i_0_), .Y(new_new_n470_));
  NO3        g0448(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n275_), .B(new_new_n99_), .Y(new_new_n472_));
  NA2        g0450(.A(new_new_n472_), .B(new_new_n471_), .Y(new_new_n473_));
  NA2        g0451(.A(i_8_), .B(i_9_), .Y(new_new_n474_));
  AOI210     g0452(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n475_));
  OR2        g0453(.A(new_new_n475_), .B(new_new_n474_), .Y(new_new_n476_));
  NA2        g0454(.A(new_new_n289_), .B(new_new_n208_), .Y(new_new_n477_));
  NO2        g0455(.A(new_new_n477_), .B(new_new_n476_), .Y(new_new_n478_));
  NA2        g0456(.A(new_new_n256_), .B(new_new_n315_), .Y(new_new_n479_));
  NO3        g0457(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n480_));
  AOI210     g0458(.A0(new_new_n262_), .A1(new_new_n191_), .B0(new_new_n480_), .Y(new_new_n481_));
  NA3        g0459(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n482_));
  NA4        g0460(.A(new_new_n146_), .B(new_new_n117_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n483_));
  OAI220     g0461(.A0(new_new_n483_), .A1(new_new_n482_), .B0(new_new_n481_), .B1(new_new_n479_), .Y(new_new_n484_));
  NO2        g0462(.A(new_new_n484_), .B(new_new_n478_), .Y(new_new_n485_));
  INV        g0463(.A(new_new_n302_), .Y(new_new_n486_));
  OR2        g0464(.A(new_new_n486_), .B(new_new_n210_), .Y(new_new_n487_));
  OA210      g0465(.A0(new_new_n363_), .A1(new_new_n103_), .B0(new_new_n304_), .Y(new_new_n488_));
  OA220      g0466(.A0(new_new_n488_), .A1(new_new_n163_), .B0(new_new_n487_), .B1(new_new_n236_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n98_), .B(i_13_), .Y(new_new_n490_));
  NA2        g0468(.A(new_new_n446_), .B(new_new_n393_), .Y(new_new_n491_));
  NO2        g0469(.A(i_2_), .B(i_13_), .Y(new_new_n492_));
  NO2        g0470(.A(new_new_n491_), .B(new_new_n490_), .Y(new_new_n493_));
  NO3        g0471(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n494_));
  NO2        g0472(.A(i_6_), .B(i_7_), .Y(new_new_n495_));
  NA2        g0473(.A(new_new_n495_), .B(new_new_n494_), .Y(new_new_n496_));
  NO2        g0474(.A(i_11_), .B(i_1_), .Y(new_new_n497_));
  NO2        g0475(.A(new_new_n73_), .B(i_3_), .Y(new_new_n498_));
  OR2        g0476(.A(i_11_), .B(i_8_), .Y(new_new_n499_));
  NOi21      g0477(.An(i_2_), .B(i_7_), .Y(new_new_n500_));
  NAi31      g0478(.An(new_new_n499_), .B(new_new_n500_), .C(new_new_n498_), .Y(new_new_n501_));
  NO2        g0479(.A(new_new_n434_), .B(i_6_), .Y(new_new_n502_));
  NA2        g0480(.A(new_new_n502_), .B(new_new_n464_), .Y(new_new_n503_));
  NO2        g0481(.A(new_new_n503_), .B(new_new_n501_), .Y(new_new_n504_));
  NO2        g0482(.A(i_3_), .B(new_new_n196_), .Y(new_new_n505_));
  NO2        g0483(.A(i_6_), .B(i_10_), .Y(new_new_n506_));
  NA4        g0484(.A(new_new_n506_), .B(new_new_n320_), .C(new_new_n505_), .D(new_new_n241_), .Y(new_new_n507_));
  NO2        g0485(.A(new_new_n507_), .B(new_new_n156_), .Y(new_new_n508_));
  NA3        g0486(.A(new_new_n250_), .B(new_new_n173_), .C(new_new_n133_), .Y(new_new_n509_));
  NA2        g0487(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n510_));
  NO2        g0488(.A(new_new_n158_), .B(i_3_), .Y(new_new_n511_));
  NAi31      g0489(.An(new_new_n510_), .B(new_new_n511_), .C(new_new_n230_), .Y(new_new_n512_));
  NA3        g0490(.A(new_new_n406_), .B(new_new_n181_), .C(new_new_n150_), .Y(new_new_n513_));
  NA3        g0491(.A(new_new_n513_), .B(new_new_n512_), .C(new_new_n509_), .Y(new_new_n514_));
  NO4        g0492(.A(new_new_n514_), .B(new_new_n508_), .C(new_new_n504_), .D(new_new_n493_), .Y(new_new_n515_));
  NA2        g0493(.A(new_new_n471_), .B(new_new_n394_), .Y(new_new_n516_));
  NA2        g0494(.A(new_new_n480_), .B(new_new_n401_), .Y(new_new_n517_));
  NO2        g0495(.A(new_new_n517_), .B(new_new_n228_), .Y(new_new_n518_));
  NAi21      g0496(.An(new_new_n219_), .B(new_new_n412_), .Y(new_new_n519_));
  NO2        g0497(.A(new_new_n26_), .B(i_5_), .Y(new_new_n520_));
  NO2        g0498(.A(i_0_), .B(new_new_n86_), .Y(new_new_n521_));
  NA3        g0499(.A(new_new_n521_), .B(new_new_n520_), .C(new_new_n143_), .Y(new_new_n522_));
  OR3        g0500(.A(new_new_n310_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n523_));
  NO2        g0501(.A(new_new_n523_), .B(new_new_n522_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n27_), .B(i_10_), .Y(new_new_n525_));
  NA2        g0503(.A(new_new_n320_), .B(new_new_n243_), .Y(new_new_n526_));
  OAI220     g0504(.A0(new_new_n526_), .A1(new_new_n454_), .B0(new_new_n525_), .B1(new_new_n490_), .Y(new_new_n527_));
  NA4        g0505(.A(new_new_n313_), .B(new_new_n227_), .C(new_new_n73_), .D(new_new_n241_), .Y(new_new_n528_));
  NO2        g0506(.A(new_new_n528_), .B(new_new_n496_), .Y(new_new_n529_));
  NO4        g0507(.A(new_new_n529_), .B(new_new_n527_), .C(new_new_n524_), .D(new_new_n518_), .Y(new_new_n530_));
  NA4        g0508(.A(new_new_n530_), .B(new_new_n515_), .C(new_new_n489_), .D(new_new_n485_), .Y(new_new_n531_));
  NA3        g0509(.A(new_new_n313_), .B(new_new_n178_), .C(new_new_n176_), .Y(new_new_n532_));
  INV        g0510(.A(new_new_n532_), .Y(new_new_n533_));
  AN2        g0511(.A(new_new_n293_), .B(new_new_n238_), .Y(new_new_n534_));
  NA2        g0512(.A(new_new_n534_), .B(new_new_n533_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n123_), .B(new_new_n113_), .Y(new_new_n536_));
  AN2        g0514(.A(new_new_n536_), .B(new_new_n471_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n320_), .B(new_new_n165_), .Y(new_new_n538_));
  OAI210     g0516(.A0(new_new_n538_), .A1(new_new_n236_), .B0(new_new_n314_), .Y(new_new_n539_));
  AOI220     g0517(.A0(new_new_n539_), .A1(new_new_n332_), .B0(new_new_n537_), .B1(new_new_n316_), .Y(new_new_n540_));
  NA2        g0518(.A(new_new_n394_), .B(new_new_n229_), .Y(new_new_n541_));
  NA2        g0519(.A(new_new_n367_), .B(new_new_n73_), .Y(new_new_n542_));
  NA2        g0520(.A(new_new_n382_), .B(new_new_n377_), .Y(new_new_n543_));
  OR2        g0521(.A(new_new_n541_), .B(new_new_n543_), .Y(new_new_n544_));
  NO2        g0522(.A(new_new_n36_), .B(i_8_), .Y(new_new_n545_));
  NAi41      g0523(.An(new_new_n542_), .B(new_new_n506_), .C(new_new_n545_), .D(new_new_n47_), .Y(new_new_n546_));
  AOI210     g0524(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n435_), .Y(new_new_n547_));
  NA3        g0525(.A(new_new_n547_), .B(new_new_n546_), .C(new_new_n544_), .Y(new_new_n548_));
  INV        g0526(.A(new_new_n548_), .Y(new_new_n549_));
  NO2        g0527(.A(i_7_), .B(new_new_n202_), .Y(new_new_n550_));
  OR2        g0528(.A(new_new_n185_), .B(i_4_), .Y(new_new_n551_));
  NO2        g0529(.A(new_new_n551_), .B(new_new_n86_), .Y(new_new_n552_));
  NA2        g0530(.A(new_new_n552_), .B(new_new_n550_), .Y(new_new_n553_));
  NA4        g0531(.A(new_new_n553_), .B(new_new_n549_), .C(new_new_n540_), .D(new_new_n535_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n400_), .B(new_new_n302_), .Y(new_new_n555_));
  OAI210     g0533(.A0(new_new_n396_), .A1(new_new_n170_), .B0(new_new_n555_), .Y(new_new_n556_));
  NO2        g0534(.A(i_12_), .B(new_new_n196_), .Y(new_new_n557_));
  NA2        g0535(.A(new_new_n557_), .B(new_new_n229_), .Y(new_new_n558_));
  NA2        g0536(.A(new_new_n506_), .B(new_new_n27_), .Y(new_new_n559_));
  NO2        g0537(.A(new_new_n559_), .B(new_new_n558_), .Y(new_new_n560_));
  NOi31      g0538(.An(new_new_n323_), .B(new_new_n434_), .C(new_new_n38_), .Y(new_new_n561_));
  OAI210     g0539(.A0(new_new_n561_), .A1(new_new_n560_), .B0(new_new_n556_), .Y(new_new_n562_));
  NO2        g0540(.A(i_8_), .B(i_7_), .Y(new_new_n563_));
  OAI210     g0541(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n564_));
  NA2        g0542(.A(new_new_n564_), .B(new_new_n227_), .Y(new_new_n565_));
  AOI220     g0543(.A0(new_new_n333_), .A1(new_new_n40_), .B0(new_new_n239_), .B1(new_new_n209_), .Y(new_new_n566_));
  OAI220     g0544(.A0(new_new_n566_), .A1(new_new_n551_), .B0(new_new_n565_), .B1(new_new_n247_), .Y(new_new_n567_));
  NA2        g0545(.A(new_new_n45_), .B(i_10_), .Y(new_new_n568_));
  NO2        g0546(.A(new_new_n568_), .B(i_6_), .Y(new_new_n569_));
  NA3        g0547(.A(new_new_n569_), .B(new_new_n567_), .C(new_new_n563_), .Y(new_new_n570_));
  AOI220     g0548(.A0(new_new_n446_), .A1(new_new_n333_), .B0(new_new_n252_), .B1(new_new_n249_), .Y(new_new_n571_));
  OAI220     g0549(.A0(new_new_n571_), .A1(new_new_n271_), .B0(new_new_n490_), .B1(new_new_n134_), .Y(new_new_n572_));
  NA2        g0550(.A(new_new_n572_), .B(new_new_n274_), .Y(new_new_n573_));
  NOi31      g0551(.An(new_new_n297_), .B(new_new_n308_), .C(new_new_n183_), .Y(new_new_n574_));
  NA3        g0552(.A(new_new_n313_), .B(new_new_n176_), .C(new_new_n98_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n225_), .B(new_new_n45_), .Y(new_new_n576_));
  NO2        g0554(.A(new_new_n158_), .B(i_5_), .Y(new_new_n577_));
  NA3        g0555(.A(new_new_n577_), .B(new_new_n422_), .C(new_new_n326_), .Y(new_new_n578_));
  OAI210     g0556(.A0(new_new_n578_), .A1(new_new_n576_), .B0(new_new_n575_), .Y(new_new_n579_));
  OAI210     g0557(.A0(new_new_n579_), .A1(new_new_n574_), .B0(new_new_n480_), .Y(new_new_n580_));
  NA4        g0558(.A(new_new_n580_), .B(new_new_n573_), .C(new_new_n570_), .D(new_new_n562_), .Y(new_new_n581_));
  NA3        g0559(.A(new_new_n221_), .B(new_new_n71_), .C(new_new_n45_), .Y(new_new_n582_));
  NA2        g0560(.A(new_new_n289_), .B(new_new_n84_), .Y(new_new_n583_));
  AOI210     g0561(.A0(new_new_n582_), .A1(new_new_n358_), .B0(new_new_n583_), .Y(new_new_n584_));
  NA2        g0562(.A(new_new_n303_), .B(new_new_n293_), .Y(new_new_n585_));
  NO2        g0563(.A(new_new_n585_), .B(new_new_n175_), .Y(new_new_n586_));
  NA2        g0564(.A(new_new_n227_), .B(new_new_n226_), .Y(new_new_n587_));
  NA2        g0565(.A(new_new_n466_), .B(new_new_n225_), .Y(new_new_n588_));
  NO2        g0566(.A(new_new_n587_), .B(new_new_n588_), .Y(new_new_n589_));
  AOI210     g0567(.A0(i_6_), .A1(new_new_n47_), .B0(new_new_n379_), .Y(new_new_n590_));
  NA2        g0568(.A(i_0_), .B(new_new_n49_), .Y(new_new_n591_));
  NA3        g0569(.A(new_new_n557_), .B(new_new_n280_), .C(new_new_n591_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n590_), .B(new_new_n592_), .Y(new_new_n593_));
  NO4        g0571(.A(new_new_n593_), .B(new_new_n589_), .C(new_new_n586_), .D(new_new_n584_), .Y(new_new_n594_));
  NO4        g0572(.A(new_new_n257_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n595_));
  NO3        g0573(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n237_), .B(new_new_n36_), .Y(new_new_n597_));
  AN2        g0575(.A(new_new_n597_), .B(new_new_n596_), .Y(new_new_n598_));
  OA210      g0576(.A0(new_new_n598_), .A1(new_new_n595_), .B0(new_new_n367_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n434_), .B(i_1_), .Y(new_new_n600_));
  NOi31      g0578(.An(new_new_n600_), .B(new_new_n472_), .C(new_new_n73_), .Y(new_new_n601_));
  AN4        g0579(.A(new_new_n601_), .B(new_new_n431_), .C(new_new_n520_), .D(i_2_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n444_), .B(new_new_n179_), .Y(new_new_n603_));
  NO3        g0581(.A(new_new_n603_), .B(new_new_n602_), .C(new_new_n599_), .Y(new_new_n604_));
  NOi21      g0582(.An(i_10_), .B(i_6_), .Y(new_new_n605_));
  NO2        g0583(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n606_));
  NO2        g0584(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n607_));
  NA2        g0585(.A(new_new_n323_), .B(new_new_n165_), .Y(new_new_n608_));
  AOI220     g0586(.A0(new_new_n608_), .A1(new_new_n455_), .B0(new_new_n186_), .B1(new_new_n184_), .Y(new_new_n609_));
  NOi31      g0587(.An(new_new_n147_), .B(i_1_), .C(new_new_n340_), .Y(new_new_n610_));
  NO2        g0588(.A(new_new_n610_), .B(new_new_n609_), .Y(new_new_n611_));
  NO2        g0589(.A(new_new_n542_), .B(new_new_n389_), .Y(new_new_n612_));
  INV        g0590(.A(new_new_n326_), .Y(new_new_n613_));
  NO2        g0591(.A(i_12_), .B(new_new_n86_), .Y(new_new_n614_));
  NO3        g0592(.A(i_4_), .B(new_new_n351_), .C(new_new_n308_), .Y(new_new_n615_));
  OR2        g0593(.A(i_2_), .B(i_5_), .Y(new_new_n616_));
  OR2        g0594(.A(new_new_n616_), .B(new_new_n426_), .Y(new_new_n617_));
  AOI210     g0595(.A0(new_new_n384_), .A1(new_new_n249_), .B0(new_new_n201_), .Y(new_new_n618_));
  AOI210     g0596(.A0(new_new_n618_), .A1(new_new_n617_), .B0(new_new_n519_), .Y(new_new_n619_));
  NO3        g0597(.A(new_new_n619_), .B(new_new_n615_), .C(new_new_n612_), .Y(new_new_n620_));
  NA4        g0598(.A(new_new_n620_), .B(new_new_n611_), .C(new_new_n604_), .D(new_new_n594_), .Y(new_new_n621_));
  NO4        g0599(.A(new_new_n621_), .B(new_new_n581_), .C(new_new_n554_), .D(new_new_n531_), .Y(new_new_n622_));
  NA4        g0600(.A(new_new_n622_), .B(new_new_n463_), .C(new_new_n366_), .D(new_new_n319_), .Y(mai7));
  NO2        g0601(.A(new_new_n95_), .B(new_new_n55_), .Y(new_new_n624_));
  NO2        g0602(.A(new_new_n110_), .B(new_new_n92_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n506_), .B(new_new_n84_), .Y(new_new_n626_));
  NA2        g0604(.A(i_11_), .B(new_new_n196_), .Y(new_new_n627_));
  NA3        g0605(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n628_));
  NO2        g0606(.A(new_new_n241_), .B(i_4_), .Y(new_new_n629_));
  NA2        g0607(.A(new_new_n629_), .B(i_8_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n107_), .B(new_new_n628_), .Y(new_new_n631_));
  NA2        g0609(.A(i_2_), .B(new_new_n86_), .Y(new_new_n632_));
  OAI210     g0610(.A0(new_new_n89_), .A1(new_new_n206_), .B0(new_new_n207_), .Y(new_new_n633_));
  NO2        g0611(.A(i_7_), .B(new_new_n37_), .Y(new_new_n634_));
  NA2        g0612(.A(i_4_), .B(i_8_), .Y(new_new_n635_));
  AOI210     g0613(.A0(new_new_n635_), .A1(new_new_n313_), .B0(new_new_n634_), .Y(new_new_n636_));
  OAI220     g0614(.A0(new_new_n636_), .A1(new_new_n632_), .B0(new_new_n633_), .B1(i_13_), .Y(new_new_n637_));
  NO3        g0615(.A(new_new_n637_), .B(new_new_n631_), .C(new_new_n624_), .Y(new_new_n638_));
  AOI210     g0616(.A0(new_new_n129_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n639_));
  AOI210     g0617(.A0(new_new_n639_), .A1(new_new_n241_), .B0(new_new_n162_), .Y(new_new_n640_));
  OR2        g0618(.A(i_6_), .B(i_10_), .Y(new_new_n641_));
  NO2        g0619(.A(new_new_n641_), .B(new_new_n23_), .Y(new_new_n642_));
  OR3        g0620(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n643_));
  NO3        g0621(.A(new_new_n643_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n644_));
  INV        g0622(.A(new_new_n203_), .Y(new_new_n645_));
  NO2        g0623(.A(new_new_n644_), .B(new_new_n642_), .Y(new_new_n646_));
  OA220      g0624(.A0(new_new_n646_), .A1(new_new_n613_), .B0(new_new_n640_), .B1(new_new_n276_), .Y(new_new_n647_));
  AOI210     g0625(.A0(new_new_n647_), .A1(new_new_n638_), .B0(new_new_n63_), .Y(new_new_n648_));
  NOi21      g0626(.An(i_11_), .B(i_7_), .Y(new_new_n649_));
  AO210      g0627(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n650_));
  NO2        g0628(.A(new_new_n650_), .B(new_new_n649_), .Y(new_new_n651_));
  NA2        g0629(.A(new_new_n651_), .B(new_new_n209_), .Y(new_new_n652_));
  NA3        g0630(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n653_));
  NAi31      g0631(.An(new_new_n653_), .B(new_new_n218_), .C(i_11_), .Y(new_new_n654_));
  AOI210     g0632(.A0(new_new_n654_), .A1(new_new_n652_), .B0(new_new_n63_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n88_), .B(new_new_n63_), .Y(new_new_n656_));
  AO210      g0634(.A0(new_new_n656_), .A1(new_new_n389_), .B0(new_new_n41_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n230_), .B(new_new_n63_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n63_), .B(i_9_), .Y(new_new_n659_));
  NO2        g0637(.A(i_1_), .B(i_12_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n658_), .B(new_new_n657_), .Y(new_new_n661_));
  OAI210     g0639(.A0(new_new_n661_), .A1(new_new_n655_), .B0(i_6_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n653_), .B(new_new_n110_), .Y(new_new_n663_));
  NA2        g0641(.A(new_new_n663_), .B(new_new_n614_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n241_), .B(new_new_n86_), .Y(new_new_n665_));
  NO2        g0643(.A(new_new_n665_), .B(i_11_), .Y(new_new_n666_));
  NA2        g0644(.A(new_new_n664_), .B(new_new_n473_), .Y(new_new_n667_));
  NO4        g0645(.A(new_new_n218_), .B(new_new_n129_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n668_));
  NA2        g0646(.A(new_new_n668_), .B(new_new_n659_), .Y(new_new_n669_));
  NA2        g0647(.A(new_new_n241_), .B(i_6_), .Y(new_new_n670_));
  NO3        g0648(.A(new_new_n641_), .B(new_new_n237_), .C(new_new_n23_), .Y(new_new_n671_));
  AOI210     g0649(.A0(i_1_), .A1(new_new_n266_), .B0(new_new_n671_), .Y(new_new_n672_));
  OAI210     g0650(.A0(new_new_n672_), .A1(new_new_n45_), .B0(new_new_n669_), .Y(new_new_n673_));
  NA3        g0651(.A(new_new_n563_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n674_));
  NA2        g0652(.A(new_new_n139_), .B(i_9_), .Y(new_new_n675_));
  NA3        g0653(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n676_));
  NO2        g0654(.A(new_new_n47_), .B(i_1_), .Y(new_new_n677_));
  NO2        g0655(.A(new_new_n675_), .B(new_new_n1072_), .Y(new_new_n678_));
  NA3        g0656(.A(new_new_n659_), .B(new_new_n326_), .C(i_6_), .Y(new_new_n679_));
  NO2        g0657(.A(new_new_n679_), .B(new_new_n23_), .Y(new_new_n680_));
  AOI210     g0658(.A0(new_new_n497_), .A1(new_new_n437_), .B0(new_new_n246_), .Y(new_new_n681_));
  NO2        g0659(.A(new_new_n681_), .B(new_new_n632_), .Y(new_new_n682_));
  NAi21      g0660(.An(new_new_n674_), .B(new_new_n94_), .Y(new_new_n683_));
  NA2        g0661(.A(new_new_n677_), .B(new_new_n275_), .Y(new_new_n684_));
  NO2        g0662(.A(i_11_), .B(new_new_n37_), .Y(new_new_n685_));
  NA2        g0663(.A(new_new_n685_), .B(new_new_n24_), .Y(new_new_n686_));
  OAI210     g0664(.A0(new_new_n686_), .A1(new_new_n684_), .B0(new_new_n683_), .Y(new_new_n687_));
  OR4        g0665(.A(new_new_n687_), .B(new_new_n682_), .C(new_new_n680_), .D(new_new_n678_), .Y(new_new_n688_));
  NO3        g0666(.A(new_new_n688_), .B(new_new_n673_), .C(new_new_n667_), .Y(new_new_n689_));
  NO2        g0667(.A(new_new_n241_), .B(new_new_n103_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n690_), .B(new_new_n649_), .Y(new_new_n691_));
  NA2        g0669(.A(new_new_n691_), .B(i_1_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n692_), .B(new_new_n643_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n433_), .B(new_new_n86_), .Y(new_new_n694_));
  NA2        g0672(.A(new_new_n693_), .B(new_new_n47_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n237_), .B(new_new_n45_), .Y(new_new_n696_));
  NO3        g0674(.A(new_new_n696_), .B(new_new_n316_), .C(new_new_n242_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n118_), .B(new_new_n37_), .Y(new_new_n698_));
  NO2        g0676(.A(new_new_n698_), .B(i_6_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n86_), .B(i_9_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n700_), .B(new_new_n63_), .Y(new_new_n701_));
  NO2        g0679(.A(new_new_n701_), .B(new_new_n660_), .Y(new_new_n702_));
  NO4        g0680(.A(new_new_n702_), .B(new_new_n699_), .C(new_new_n697_), .D(i_4_), .Y(new_new_n703_));
  NA2        g0681(.A(i_1_), .B(i_3_), .Y(new_new_n704_));
  INV        g0682(.A(new_new_n703_), .Y(new_new_n705_));
  NA4        g0683(.A(new_new_n705_), .B(new_new_n695_), .C(new_new_n689_), .D(new_new_n662_), .Y(new_new_n706_));
  NO3        g0684(.A(new_new_n499_), .B(i_3_), .C(i_7_), .Y(new_new_n707_));
  NOi21      g0685(.An(new_new_n707_), .B(i_10_), .Y(new_new_n708_));
  OA210      g0686(.A0(new_new_n708_), .A1(new_new_n250_), .B0(new_new_n86_), .Y(new_new_n709_));
  NA3        g0687(.A(new_new_n506_), .B(new_new_n545_), .C(new_new_n47_), .Y(new_new_n710_));
  NA3        g0688(.A(new_new_n162_), .B(new_new_n84_), .C(new_new_n86_), .Y(new_new_n711_));
  NA2        g0689(.A(new_new_n711_), .B(new_new_n710_), .Y(new_new_n712_));
  OAI210     g0690(.A0(new_new_n712_), .A1(new_new_n709_), .B0(i_1_), .Y(new_new_n713_));
  AOI210     g0691(.A0(new_new_n275_), .A1(new_new_n99_), .B0(i_1_), .Y(new_new_n714_));
  NO2        g0692(.A(new_new_n380_), .B(i_2_), .Y(new_new_n715_));
  NA2        g0693(.A(new_new_n715_), .B(new_new_n714_), .Y(new_new_n716_));
  OAI210     g0694(.A0(new_new_n679_), .A1(new_new_n467_), .B0(new_new_n716_), .Y(new_new_n717_));
  INV        g0695(.A(new_new_n717_), .Y(new_new_n718_));
  AOI210     g0696(.A0(new_new_n718_), .A1(new_new_n713_), .B0(i_13_), .Y(new_new_n719_));
  OR2        g0697(.A(i_11_), .B(i_7_), .Y(new_new_n720_));
  NA3        g0698(.A(new_new_n720_), .B(new_new_n108_), .C(new_new_n139_), .Y(new_new_n721_));
  AOI220     g0699(.A0(new_new_n492_), .A1(new_new_n162_), .B0(new_new_n469_), .B1(new_new_n139_), .Y(new_new_n722_));
  OAI210     g0700(.A0(new_new_n722_), .A1(new_new_n45_), .B0(new_new_n721_), .Y(new_new_n723_));
  NO2        g0701(.A(new_new_n55_), .B(i_12_), .Y(new_new_n724_));
  NO2        g0702(.A(new_new_n500_), .B(new_new_n24_), .Y(new_new_n725_));
  AOI220     g0703(.A0(new_new_n725_), .A1(new_new_n694_), .B0(new_new_n250_), .B1(new_new_n132_), .Y(new_new_n726_));
  OAI220     g0704(.A0(new_new_n726_), .A1(new_new_n41_), .B0(new_new_n1071_), .B1(new_new_n95_), .Y(new_new_n727_));
  AOI210     g0705(.A0(new_new_n723_), .A1(new_new_n342_), .B0(new_new_n727_), .Y(new_new_n728_));
  NA2        g0706(.A(new_new_n397_), .B(new_new_n677_), .Y(new_new_n729_));
  NO2        g0707(.A(new_new_n729_), .B(new_new_n247_), .Y(new_new_n730_));
  AOI210     g0708(.A0(new_new_n467_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n731_));
  NOi31      g0709(.An(new_new_n731_), .B(new_new_n626_), .C(new_new_n45_), .Y(new_new_n732_));
  NA2        g0710(.A(new_new_n128_), .B(i_13_), .Y(new_new_n733_));
  NO2        g0711(.A(new_new_n676_), .B(new_new_n116_), .Y(new_new_n734_));
  INV        g0712(.A(new_new_n734_), .Y(new_new_n735_));
  NO2        g0713(.A(new_new_n733_), .B(new_new_n714_), .Y(new_new_n736_));
  NA2        g0714(.A(new_new_n26_), .B(new_new_n196_), .Y(new_new_n737_));
  INV        g0715(.A(i_7_), .Y(new_new_n738_));
  AOI220     g0716(.A0(new_new_n397_), .A1(new_new_n677_), .B0(new_new_n94_), .B1(new_new_n104_), .Y(new_new_n739_));
  NO2        g0717(.A(new_new_n739_), .B(new_new_n630_), .Y(new_new_n740_));
  NO4        g0718(.A(new_new_n740_), .B(new_new_n736_), .C(new_new_n732_), .D(new_new_n730_), .Y(new_new_n741_));
  OR2        g0719(.A(i_11_), .B(i_6_), .Y(new_new_n742_));
  NA3        g0720(.A(new_new_n629_), .B(new_new_n737_), .C(i_7_), .Y(new_new_n743_));
  AOI210     g0721(.A0(new_new_n743_), .A1(new_new_n735_), .B0(new_new_n742_), .Y(new_new_n744_));
  NA3        g0722(.A(new_new_n427_), .B(new_new_n634_), .C(new_new_n99_), .Y(new_new_n745_));
  NA2        g0723(.A(new_new_n666_), .B(i_13_), .Y(new_new_n746_));
  NAi21      g0724(.An(i_11_), .B(i_12_), .Y(new_new_n747_));
  NOi41      g0725(.An(new_new_n112_), .B(new_new_n747_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n748_));
  NA2        g0726(.A(new_new_n748_), .B(new_new_n47_), .Y(new_new_n749_));
  NA3        g0727(.A(new_new_n749_), .B(new_new_n746_), .C(new_new_n745_), .Y(new_new_n750_));
  OAI210     g0728(.A0(new_new_n750_), .A1(new_new_n744_), .B0(new_new_n63_), .Y(new_new_n751_));
  NO2        g0729(.A(i_2_), .B(i_12_), .Y(new_new_n752_));
  NA2        g0730(.A(new_new_n379_), .B(new_new_n752_), .Y(new_new_n753_));
  NA2        g0731(.A(i_8_), .B(new_new_n25_), .Y(new_new_n754_));
  NO3        g0732(.A(new_new_n754_), .B(new_new_n395_), .C(new_new_n629_), .Y(new_new_n755_));
  OAI210     g0733(.A0(new_new_n755_), .A1(new_new_n381_), .B0(new_new_n379_), .Y(new_new_n756_));
  NO2        g0734(.A(new_new_n129_), .B(i_2_), .Y(new_new_n757_));
  NA2        g0735(.A(new_new_n756_), .B(new_new_n753_), .Y(new_new_n758_));
  NA3        g0736(.A(new_new_n758_), .B(new_new_n46_), .C(new_new_n229_), .Y(new_new_n759_));
  NA4        g0737(.A(new_new_n759_), .B(new_new_n751_), .C(new_new_n741_), .D(new_new_n728_), .Y(new_new_n760_));
  OR4        g0738(.A(new_new_n760_), .B(new_new_n719_), .C(new_new_n706_), .D(new_new_n648_), .Y(mai5));
  NA2        g0739(.A(new_new_n691_), .B(new_new_n277_), .Y(new_new_n762_));
  AN2        g0740(.A(new_new_n24_), .B(i_10_), .Y(new_new_n763_));
  NA3        g0741(.A(new_new_n763_), .B(new_new_n752_), .C(new_new_n110_), .Y(new_new_n764_));
  NO2        g0742(.A(new_new_n630_), .B(i_11_), .Y(new_new_n765_));
  NA2        g0743(.A(new_new_n89_), .B(new_new_n765_), .Y(new_new_n766_));
  NA3        g0744(.A(new_new_n766_), .B(new_new_n764_), .C(new_new_n762_), .Y(new_new_n767_));
  NO3        g0745(.A(i_11_), .B(new_new_n241_), .C(i_13_), .Y(new_new_n768_));
  NO2        g0746(.A(new_new_n125_), .B(new_new_n23_), .Y(new_new_n769_));
  NA2        g0747(.A(i_12_), .B(i_8_), .Y(new_new_n770_));
  OAI210     g0748(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n770_), .Y(new_new_n771_));
  INV        g0749(.A(new_new_n466_), .Y(new_new_n772_));
  AOI220     g0750(.A0(new_new_n326_), .A1(new_new_n607_), .B0(new_new_n771_), .B1(new_new_n769_), .Y(new_new_n773_));
  INV        g0751(.A(new_new_n773_), .Y(new_new_n774_));
  NO2        g0752(.A(new_new_n774_), .B(new_new_n767_), .Y(new_new_n775_));
  INV        g0753(.A(new_new_n173_), .Y(new_new_n776_));
  INV        g0754(.A(new_new_n250_), .Y(new_new_n777_));
  OAI210     g0755(.A0(new_new_n715_), .A1(new_new_n468_), .B0(new_new_n112_), .Y(new_new_n778_));
  AOI210     g0756(.A0(new_new_n778_), .A1(new_new_n777_), .B0(new_new_n776_), .Y(new_new_n779_));
  NO2        g0757(.A(new_new_n474_), .B(new_new_n26_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n780_), .B(new_new_n437_), .Y(new_new_n781_));
  NA2        g0759(.A(new_new_n781_), .B(i_2_), .Y(new_new_n782_));
  INV        g0760(.A(new_new_n782_), .Y(new_new_n783_));
  AOI210     g0761(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n434_), .Y(new_new_n784_));
  AOI210     g0762(.A0(new_new_n784_), .A1(new_new_n783_), .B0(new_new_n779_), .Y(new_new_n785_));
  NO2        g0763(.A(new_new_n193_), .B(new_new_n126_), .Y(new_new_n786_));
  OAI210     g0764(.A0(new_new_n786_), .A1(new_new_n769_), .B0(i_2_), .Y(new_new_n787_));
  INV        g0765(.A(new_new_n174_), .Y(new_new_n788_));
  NO3        g0766(.A(new_new_n650_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n789_));
  AOI210     g0767(.A0(new_new_n788_), .A1(new_new_n89_), .B0(new_new_n789_), .Y(new_new_n790_));
  AOI210     g0768(.A0(new_new_n790_), .A1(new_new_n787_), .B0(new_new_n196_), .Y(new_new_n791_));
  OA210      g0769(.A0(new_new_n651_), .A1(new_new_n127_), .B0(i_13_), .Y(new_new_n792_));
  NA2        g0770(.A(new_new_n152_), .B(new_new_n627_), .Y(new_new_n793_));
  NO2        g0771(.A(new_new_n793_), .B(new_new_n384_), .Y(new_new_n794_));
  AOI210     g0772(.A0(new_new_n211_), .A1(new_new_n149_), .B0(new_new_n545_), .Y(new_new_n795_));
  NA2        g0773(.A(new_new_n795_), .B(new_new_n437_), .Y(new_new_n796_));
  NO2        g0774(.A(new_new_n104_), .B(new_new_n45_), .Y(new_new_n797_));
  INV        g0775(.A(new_new_n309_), .Y(new_new_n798_));
  NA4        g0776(.A(new_new_n798_), .B(new_new_n313_), .C(new_new_n125_), .D(new_new_n43_), .Y(new_new_n799_));
  OAI210     g0777(.A0(new_new_n799_), .A1(new_new_n797_), .B0(new_new_n796_), .Y(new_new_n800_));
  NO4        g0778(.A(new_new_n800_), .B(new_new_n794_), .C(new_new_n792_), .D(new_new_n791_), .Y(new_new_n801_));
  NA2        g0779(.A(new_new_n607_), .B(new_new_n28_), .Y(new_new_n802_));
  NA2        g0780(.A(new_new_n768_), .B(new_new_n281_), .Y(new_new_n803_));
  NA2        g0781(.A(new_new_n803_), .B(new_new_n802_), .Y(new_new_n804_));
  NO2        g0782(.A(new_new_n62_), .B(i_12_), .Y(new_new_n805_));
  NO2        g0783(.A(new_new_n805_), .B(new_new_n127_), .Y(new_new_n806_));
  NO2        g0784(.A(new_new_n806_), .B(new_new_n627_), .Y(new_new_n807_));
  AOI220     g0785(.A0(new_new_n807_), .A1(new_new_n36_), .B0(new_new_n804_), .B1(new_new_n47_), .Y(new_new_n808_));
  NA4        g0786(.A(new_new_n808_), .B(new_new_n801_), .C(new_new_n785_), .D(new_new_n775_), .Y(mai6));
  NO3        g0787(.A(new_new_n261_), .B(new_new_n315_), .C(i_1_), .Y(new_new_n810_));
  NO2        g0788(.A(new_new_n188_), .B(new_new_n140_), .Y(new_new_n811_));
  OAI210     g0789(.A0(new_new_n811_), .A1(new_new_n810_), .B0(new_new_n757_), .Y(new_new_n812_));
  NO2        g0790(.A(new_new_n224_), .B(new_new_n510_), .Y(new_new_n813_));
  NO2        g0791(.A(i_11_), .B(i_9_), .Y(new_new_n814_));
  INV        g0792(.A(new_new_n338_), .Y(new_new_n815_));
  AO210      g0793(.A0(new_new_n815_), .A1(new_new_n812_), .B0(i_12_), .Y(new_new_n816_));
  NA2        g0794(.A(new_new_n385_), .B(new_new_n345_), .Y(new_new_n817_));
  NA2        g0795(.A(new_new_n614_), .B(new_new_n63_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n708_), .B(new_new_n71_), .Y(new_new_n819_));
  BUFFER     g0797(.A(new_new_n656_), .Y(new_new_n820_));
  NA4        g0798(.A(new_new_n820_), .B(new_new_n819_), .C(new_new_n818_), .D(new_new_n817_), .Y(new_new_n821_));
  INV        g0799(.A(new_new_n200_), .Y(new_new_n822_));
  AOI220     g0800(.A0(new_new_n822_), .A1(new_new_n814_), .B0(new_new_n821_), .B1(new_new_n73_), .Y(new_new_n823_));
  INV        g0801(.A(new_new_n337_), .Y(new_new_n824_));
  NA2        g0802(.A(new_new_n75_), .B(new_new_n132_), .Y(new_new_n825_));
  INV        g0803(.A(new_new_n125_), .Y(new_new_n826_));
  NA2        g0804(.A(new_new_n826_), .B(new_new_n47_), .Y(new_new_n827_));
  AOI210     g0805(.A0(new_new_n827_), .A1(new_new_n825_), .B0(new_new_n824_), .Y(new_new_n828_));
  NO2        g0806(.A(new_new_n257_), .B(i_9_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n829_), .B(new_new_n805_), .Y(new_new_n830_));
  AOI210     g0808(.A0(new_new_n830_), .A1(new_new_n543_), .B0(new_new_n188_), .Y(new_new_n831_));
  NO2        g0809(.A(new_new_n32_), .B(i_11_), .Y(new_new_n832_));
  NA3        g0810(.A(new_new_n832_), .B(new_new_n495_), .C(new_new_n401_), .Y(new_new_n833_));
  NAi32      g0811(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n834_));
  AOI210     g0812(.A0(new_new_n742_), .A1(new_new_n87_), .B0(new_new_n834_), .Y(new_new_n835_));
  OAI210     g0813(.A0(new_new_n707_), .A1(new_new_n597_), .B0(new_new_n596_), .Y(new_new_n836_));
  NAi31      g0814(.An(new_new_n835_), .B(new_new_n836_), .C(new_new_n833_), .Y(new_new_n837_));
  OR3        g0815(.A(new_new_n837_), .B(new_new_n831_), .C(new_new_n828_), .Y(new_new_n838_));
  NO2        g0816(.A(new_new_n720_), .B(i_2_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n840_));
  OAI210     g0818(.A0(new_new_n840_), .A1(new_new_n426_), .B0(new_new_n372_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n841_), .B(new_new_n839_), .Y(new_new_n842_));
  AO220      g0820(.A0(new_new_n371_), .A1(new_new_n362_), .B0(new_new_n409_), .B1(new_new_n627_), .Y(new_new_n843_));
  NA3        g0821(.A(new_new_n843_), .B(new_new_n262_), .C(i_7_), .Y(new_new_n844_));
  BUFFER     g0822(.A(new_new_n651_), .Y(new_new_n845_));
  NA3        g0823(.A(new_new_n845_), .B(new_new_n148_), .C(new_new_n69_), .Y(new_new_n846_));
  AO210      g0824(.A0(new_new_n517_), .A1(new_new_n772_), .B0(new_new_n36_), .Y(new_new_n847_));
  NA4        g0825(.A(new_new_n847_), .B(new_new_n846_), .C(new_new_n844_), .D(new_new_n842_), .Y(new_new_n848_));
  OAI210     g0826(.A0(new_new_n665_), .A1(i_11_), .B0(new_new_n87_), .Y(new_new_n849_));
  AOI220     g0827(.A0(new_new_n849_), .A1(new_new_n596_), .B0(new_new_n813_), .B1(new_new_n738_), .Y(new_new_n850_));
  NA2        g0828(.A(new_new_n409_), .B(new_new_n70_), .Y(new_new_n851_));
  NA3        g0829(.A(new_new_n851_), .B(new_new_n850_), .C(new_new_n633_), .Y(new_new_n852_));
  AO210      g0830(.A0(new_new_n545_), .A1(new_new_n47_), .B0(new_new_n88_), .Y(new_new_n853_));
  NA3        g0831(.A(new_new_n853_), .B(new_new_n506_), .C(new_new_n221_), .Y(new_new_n854_));
  AOI210     g0832(.A0(new_new_n468_), .A1(new_new_n466_), .B0(new_new_n595_), .Y(new_new_n855_));
  NO2        g0833(.A(new_new_n641_), .B(new_new_n104_), .Y(new_new_n856_));
  OAI210     g0834(.A0(new_new_n856_), .A1(new_new_n113_), .B0(new_new_n424_), .Y(new_new_n857_));
  NA2        g0835(.A(new_new_n249_), .B(new_new_n47_), .Y(new_new_n858_));
  INV        g0836(.A(new_new_n617_), .Y(new_new_n859_));
  NA3        g0837(.A(new_new_n859_), .B(new_new_n337_), .C(i_7_), .Y(new_new_n860_));
  NA4        g0838(.A(new_new_n860_), .B(new_new_n857_), .C(new_new_n855_), .D(new_new_n854_), .Y(new_new_n861_));
  NO4        g0839(.A(new_new_n861_), .B(new_new_n852_), .C(new_new_n848_), .D(new_new_n838_), .Y(new_new_n862_));
  NA4        g0840(.A(new_new_n862_), .B(new_new_n823_), .C(new_new_n816_), .D(new_new_n391_), .Y(mai3));
  NA2        g0841(.A(i_6_), .B(i_7_), .Y(new_new_n864_));
  NO2        g0842(.A(new_new_n864_), .B(i_0_), .Y(new_new_n865_));
  NO2        g0843(.A(i_11_), .B(new_new_n241_), .Y(new_new_n866_));
  OAI210     g0844(.A0(new_new_n865_), .A1(new_new_n297_), .B0(new_new_n866_), .Y(new_new_n867_));
  NO2        g0845(.A(new_new_n867_), .B(new_new_n196_), .Y(new_new_n868_));
  NO3        g0846(.A(new_new_n470_), .B(new_new_n92_), .C(new_new_n45_), .Y(new_new_n869_));
  OA210      g0847(.A0(new_new_n869_), .A1(new_new_n868_), .B0(new_new_n176_), .Y(new_new_n870_));
  NOi21      g0848(.An(new_new_n98_), .B(new_new_n781_), .Y(new_new_n871_));
  AN2        g0849(.A(new_new_n472_), .B(new_new_n56_), .Y(new_new_n872_));
  NO2        g0850(.A(new_new_n872_), .B(new_new_n871_), .Y(new_new_n873_));
  NO2        g0851(.A(new_new_n873_), .B(new_new_n49_), .Y(new_new_n874_));
  NO4        g0852(.A(new_new_n387_), .B(new_new_n394_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n875_));
  NA2        g0853(.A(new_new_n188_), .B(new_new_n605_), .Y(new_new_n876_));
  NOi21      g0854(.An(new_new_n876_), .B(new_new_n875_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n731_), .B(new_new_n700_), .Y(new_new_n878_));
  NA2        g0856(.A(new_new_n343_), .B(new_new_n457_), .Y(new_new_n879_));
  OAI220     g0857(.A0(new_new_n879_), .A1(new_new_n878_), .B0(new_new_n877_), .B1(new_new_n63_), .Y(new_new_n880_));
  NOi21      g0858(.An(i_5_), .B(i_9_), .Y(new_new_n881_));
  NA2        g0859(.A(new_new_n881_), .B(new_new_n465_), .Y(new_new_n882_));
  BUFFER     g0860(.A(new_new_n275_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n883_), .B(new_new_n497_), .Y(new_new_n884_));
  NO2        g0862(.A(new_new_n177_), .B(new_new_n149_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n885_), .B(new_new_n249_), .Y(new_new_n886_));
  OAI220     g0864(.A0(new_new_n886_), .A1(new_new_n183_), .B0(new_new_n884_), .B1(new_new_n882_), .Y(new_new_n887_));
  NO4        g0865(.A(new_new_n887_), .B(new_new_n880_), .C(new_new_n874_), .D(new_new_n870_), .Y(new_new_n888_));
  NA2        g0866(.A(new_new_n188_), .B(new_new_n24_), .Y(new_new_n889_));
  NA2        g0867(.A(new_new_n320_), .B(new_new_n130_), .Y(new_new_n890_));
  NAi21      g0868(.An(new_new_n163_), .B(new_new_n457_), .Y(new_new_n891_));
  OAI220     g0869(.A0(new_new_n891_), .A1(new_new_n858_), .B0(new_new_n890_), .B1(new_new_n415_), .Y(new_new_n892_));
  INV        g0870(.A(new_new_n892_), .Y(new_new_n893_));
  NO2        g0871(.A(new_new_n401_), .B(new_new_n301_), .Y(new_new_n894_));
  NA2        g0872(.A(new_new_n894_), .B(new_new_n734_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n606_), .B(i_0_), .Y(new_new_n896_));
  INV        g0874(.A(new_new_n495_), .Y(new_new_n897_));
  AN2        g0875(.A(new_new_n98_), .B(new_new_n248_), .Y(new_new_n898_));
  NA2        g0876(.A(new_new_n768_), .B(new_new_n338_), .Y(new_new_n899_));
  AOI210     g0877(.A0(new_new_n506_), .A1(new_new_n89_), .B0(new_new_n58_), .Y(new_new_n900_));
  OAI220     g0878(.A0(new_new_n900_), .A1(new_new_n899_), .B0(new_new_n686_), .B1(new_new_n565_), .Y(new_new_n901_));
  NO2        g0879(.A(new_new_n259_), .B(new_new_n154_), .Y(new_new_n902_));
  NA2        g0880(.A(i_0_), .B(i_10_), .Y(new_new_n903_));
  AN2        g0881(.A(new_new_n902_), .B(i_6_), .Y(new_new_n904_));
  AOI220     g0882(.A0(new_new_n343_), .A1(new_new_n100_), .B0(new_new_n188_), .B1(new_new_n84_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n600_), .B(i_4_), .Y(new_new_n906_));
  NA2        g0884(.A(new_new_n191_), .B(new_new_n206_), .Y(new_new_n907_));
  OAI220     g0885(.A0(new_new_n907_), .A1(new_new_n899_), .B0(new_new_n906_), .B1(new_new_n905_), .Y(new_new_n908_));
  NO4        g0886(.A(new_new_n908_), .B(new_new_n904_), .C(new_new_n901_), .D(new_new_n898_), .Y(new_new_n909_));
  NA3        g0887(.A(new_new_n909_), .B(new_new_n895_), .C(new_new_n893_), .Y(new_new_n910_));
  NA2        g0888(.A(i_11_), .B(i_9_), .Y(new_new_n911_));
  NO2        g0889(.A(new_new_n49_), .B(i_7_), .Y(new_new_n912_));
  NA2        g0890(.A(new_new_n406_), .B(new_new_n181_), .Y(new_new_n913_));
  NA2        g0891(.A(new_new_n913_), .B(new_new_n161_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n177_), .B(i_0_), .Y(new_new_n915_));
  INV        g0893(.A(new_new_n915_), .Y(new_new_n916_));
  NA2        g0894(.A(new_new_n495_), .B(new_new_n235_), .Y(new_new_n917_));
  AOI210     g0895(.A0(new_new_n382_), .A1(new_new_n42_), .B0(new_new_n423_), .Y(new_new_n918_));
  OAI220     g0896(.A0(new_new_n918_), .A1(new_new_n882_), .B0(new_new_n917_), .B1(new_new_n916_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n919_), .B(new_new_n914_), .Y(new_new_n920_));
  NA2        g0898(.A(new_new_n685_), .B(new_new_n122_), .Y(new_new_n921_));
  NO2        g0899(.A(i_6_), .B(new_new_n921_), .Y(new_new_n922_));
  AOI210     g0900(.A0(new_new_n467_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n923_));
  NA2        g0901(.A(new_new_n173_), .B(new_new_n105_), .Y(new_new_n924_));
  INV        g0902(.A(new_new_n922_), .Y(new_new_n925_));
  NOi21      g0903(.An(i_7_), .B(i_5_), .Y(new_new_n926_));
  NOi31      g0904(.An(new_new_n926_), .B(i_0_), .C(new_new_n747_), .Y(new_new_n927_));
  NA3        g0905(.A(new_new_n927_), .B(new_new_n395_), .C(i_6_), .Y(new_new_n928_));
  OA210      g0906(.A0(new_new_n924_), .A1(new_new_n543_), .B0(new_new_n928_), .Y(new_new_n929_));
  NO3        g0907(.A(new_new_n418_), .B(new_new_n374_), .C(new_new_n370_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n269_), .B(new_new_n327_), .Y(new_new_n931_));
  NO2        g0909(.A(new_new_n747_), .B(new_new_n264_), .Y(new_new_n932_));
  AOI210     g0910(.A0(new_new_n932_), .A1(new_new_n931_), .B0(new_new_n930_), .Y(new_new_n933_));
  NA4        g0911(.A(new_new_n933_), .B(new_new_n929_), .C(new_new_n925_), .D(new_new_n920_), .Y(new_new_n934_));
  NO2        g0912(.A(new_new_n889_), .B(new_new_n244_), .Y(new_new_n935_));
  AN2        g0913(.A(new_new_n342_), .B(new_new_n338_), .Y(new_new_n936_));
  AN2        g0914(.A(new_new_n936_), .B(new_new_n885_), .Y(new_new_n937_));
  OAI210     g0915(.A0(new_new_n937_), .A1(new_new_n935_), .B0(i_10_), .Y(new_new_n938_));
  NA3        g0916(.A(new_new_n494_), .B(new_new_n427_), .C(new_new_n46_), .Y(new_new_n939_));
  OAI210     g0917(.A0(new_new_n891_), .A1(new_new_n897_), .B0(new_new_n939_), .Y(new_new_n940_));
  NO2        g0918(.A(new_new_n262_), .B(new_new_n47_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n941_), .B(new_new_n190_), .Y(new_new_n942_));
  AOI220     g0920(.A0(new_new_n942_), .A1(new_new_n495_), .B0(new_new_n940_), .B1(new_new_n73_), .Y(new_new_n943_));
  NA3        g0921(.A(new_new_n840_), .B(new_new_n393_), .C(new_new_n665_), .Y(new_new_n944_));
  NA2        g0922(.A(new_new_n95_), .B(new_new_n45_), .Y(new_new_n945_));
  NO2        g0923(.A(new_new_n75_), .B(new_new_n770_), .Y(new_new_n946_));
  AOI220     g0924(.A0(new_new_n946_), .A1(new_new_n945_), .B0(new_new_n176_), .B1(new_new_n625_), .Y(new_new_n947_));
  AOI210     g0925(.A0(new_new_n947_), .A1(new_new_n944_), .B0(new_new_n48_), .Y(new_new_n948_));
  NO3        g0926(.A(new_new_n616_), .B(new_new_n369_), .C(new_new_n24_), .Y(new_new_n949_));
  AOI210     g0927(.A0(new_new_n725_), .A1(new_new_n577_), .B0(new_new_n949_), .Y(new_new_n950_));
  NAi21      g0928(.An(i_9_), .B(i_5_), .Y(new_new_n951_));
  NO2        g0929(.A(new_new_n951_), .B(new_new_n418_), .Y(new_new_n952_));
  NO2        g0930(.A(new_new_n628_), .B(new_new_n107_), .Y(new_new_n953_));
  AOI220     g0931(.A0(new_new_n953_), .A1(i_0_), .B0(new_new_n952_), .B1(new_new_n651_), .Y(new_new_n954_));
  OAI220     g0932(.A0(new_new_n954_), .A1(new_new_n86_), .B0(new_new_n950_), .B1(new_new_n174_), .Y(new_new_n955_));
  NO3        g0933(.A(new_new_n955_), .B(new_new_n948_), .C(new_new_n548_), .Y(new_new_n956_));
  NA3        g0934(.A(new_new_n956_), .B(new_new_n943_), .C(new_new_n938_), .Y(new_new_n957_));
  NO3        g0935(.A(new_new_n957_), .B(new_new_n934_), .C(new_new_n910_), .Y(new_new_n958_));
  NO2        g0936(.A(i_0_), .B(new_new_n747_), .Y(new_new_n959_));
  NA2        g0937(.A(new_new_n73_), .B(new_new_n45_), .Y(new_new_n960_));
  NA2        g0938(.A(new_new_n903_), .B(new_new_n960_), .Y(new_new_n961_));
  NO3        g0939(.A(new_new_n107_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n962_));
  AO220      g0940(.A0(new_new_n962_), .A1(new_new_n961_), .B0(new_new_n959_), .B1(new_new_n176_), .Y(new_new_n963_));
  NO2        g0941(.A(new_new_n818_), .B(new_new_n924_), .Y(new_new_n964_));
  AOI210     g0942(.A0(new_new_n963_), .A1(new_new_n359_), .B0(new_new_n964_), .Y(new_new_n965_));
  NA2        g0943(.A(new_new_n757_), .B(new_new_n147_), .Y(new_new_n966_));
  INV        g0944(.A(new_new_n966_), .Y(new_new_n967_));
  NA3        g0945(.A(new_new_n967_), .B(new_new_n700_), .C(new_new_n73_), .Y(new_new_n968_));
  NO2        g0946(.A(new_new_n836_), .B(new_new_n418_), .Y(new_new_n969_));
  NA3        g0947(.A(new_new_n865_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n970_));
  NA2        g0948(.A(new_new_n866_), .B(i_9_), .Y(new_new_n971_));
  AOI210     g0949(.A0(new_new_n970_), .A1(new_new_n522_), .B0(new_new_n971_), .Y(new_new_n972_));
  NA2        g0950(.A(new_new_n249_), .B(new_new_n234_), .Y(new_new_n973_));
  AOI210     g0951(.A0(new_new_n973_), .A1(new_new_n896_), .B0(new_new_n154_), .Y(new_new_n974_));
  NO3        g0952(.A(new_new_n974_), .B(new_new_n972_), .C(new_new_n969_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n975_), .B(new_new_n968_), .C(new_new_n965_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n936_), .B(new_new_n384_), .Y(new_new_n977_));
  AOI210     g0955(.A0(new_new_n308_), .A1(new_new_n163_), .B0(new_new_n977_), .Y(new_new_n978_));
  NA3        g0956(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n912_), .B(new_new_n511_), .Y(new_new_n980_));
  AOI210     g0958(.A0(new_new_n979_), .A1(new_new_n163_), .B0(new_new_n980_), .Y(new_new_n981_));
  NO2        g0959(.A(new_new_n981_), .B(new_new_n978_), .Y(new_new_n982_));
  NO3        g0960(.A(new_new_n903_), .B(new_new_n881_), .C(new_new_n193_), .Y(new_new_n983_));
  AOI220     g0961(.A0(new_new_n983_), .A1(i_11_), .B0(new_new_n601_), .B1(new_new_n75_), .Y(new_new_n984_));
  NO3        g0962(.A(new_new_n212_), .B(new_new_n394_), .C(i_0_), .Y(new_new_n985_));
  OAI210     g0963(.A0(new_new_n985_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n986_));
  INV        g0964(.A(new_new_n221_), .Y(new_new_n987_));
  OAI220     g0965(.A0(new_new_n558_), .A1(new_new_n140_), .B0(new_new_n670_), .B1(new_new_n645_), .Y(new_new_n988_));
  NA3        g0966(.A(new_new_n988_), .B(new_new_n410_), .C(new_new_n987_), .Y(new_new_n989_));
  NA4        g0967(.A(new_new_n989_), .B(new_new_n986_), .C(new_new_n984_), .D(new_new_n982_), .Y(new_new_n990_));
  AOI220     g0968(.A0(new_new_n926_), .A1(new_new_n511_), .B0(new_new_n865_), .B1(new_new_n164_), .Y(new_new_n991_));
  NA2        g0969(.A(new_new_n362_), .B(new_new_n178_), .Y(new_new_n992_));
  OR2        g0970(.A(new_new_n992_), .B(new_new_n991_), .Y(new_new_n993_));
  AOI210     g0971(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n177_), .Y(new_new_n994_));
  NA3        g0972(.A(new_new_n642_), .B(new_new_n188_), .C(new_new_n84_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n995_), .B(new_new_n575_), .Y(new_new_n996_));
  NA2        g0974(.A(new_new_n516_), .B(new_new_n509_), .Y(new_new_n997_));
  NO2        g0975(.A(new_new_n997_), .B(new_new_n996_), .Y(new_new_n998_));
  NA3        g0976(.A(new_new_n912_), .B(new_new_n297_), .C(new_new_n234_), .Y(new_new_n999_));
  INV        g0977(.A(new_new_n999_), .Y(new_new_n1000_));
  NA3        g0978(.A(new_new_n401_), .B(new_new_n344_), .C(new_new_n225_), .Y(new_new_n1001_));
  INV        g0979(.A(new_new_n1001_), .Y(new_new_n1002_));
  NOi31      g0980(.An(new_new_n400_), .B(new_new_n960_), .C(new_new_n244_), .Y(new_new_n1003_));
  NO3        g0981(.A(new_new_n911_), .B(new_new_n221_), .C(new_new_n193_), .Y(new_new_n1004_));
  NO4        g0982(.A(new_new_n1004_), .B(new_new_n1003_), .C(new_new_n1002_), .D(new_new_n1000_), .Y(new_new_n1005_));
  NA3        g0983(.A(new_new_n1005_), .B(new_new_n998_), .C(new_new_n993_), .Y(new_new_n1006_));
  INV        g0984(.A(new_new_n644_), .Y(new_new_n1007_));
  NO3        g0985(.A(new_new_n1007_), .B(new_new_n591_), .C(new_new_n356_), .Y(new_new_n1008_));
  INV        g0986(.A(new_new_n1008_), .Y(new_new_n1009_));
  NA3        g0987(.A(new_new_n313_), .B(i_5_), .C(new_new_n196_), .Y(new_new_n1010_));
  NA2        g0988(.A(new_new_n1010_), .B(new_new_n247_), .Y(new_new_n1011_));
  NO4        g0989(.A(new_new_n244_), .B(new_new_n212_), .C(i_0_), .D(i_12_), .Y(new_new_n1012_));
  NA2        g0990(.A(new_new_n1012_), .B(new_new_n1011_), .Y(new_new_n1013_));
  AN2        g0991(.A(new_new_n903_), .B(new_new_n154_), .Y(new_new_n1014_));
  NO4        g0992(.A(new_new_n1014_), .B(i_12_), .C(new_new_n674_), .D(new_new_n132_), .Y(new_new_n1015_));
  NA2        g0993(.A(new_new_n1015_), .B(new_new_n221_), .Y(new_new_n1016_));
  NA3        g0994(.A(new_new_n100_), .B(new_new_n605_), .C(i_11_), .Y(new_new_n1017_));
  NO2        g0995(.A(new_new_n1017_), .B(new_new_n156_), .Y(new_new_n1018_));
  NA2        g0996(.A(new_new_n926_), .B(new_new_n492_), .Y(new_new_n1019_));
  NA2        g0997(.A(new_new_n64_), .B(new_new_n103_), .Y(new_new_n1020_));
  OAI220     g0998(.A0(new_new_n1020_), .A1(new_new_n1010_), .B0(new_new_n1019_), .B1(new_new_n701_), .Y(new_new_n1021_));
  AOI210     g0999(.A0(new_new_n1021_), .A1(new_new_n915_), .B0(new_new_n1018_), .Y(new_new_n1022_));
  NA4        g1000(.A(new_new_n1022_), .B(new_new_n1016_), .C(new_new_n1013_), .D(new_new_n1009_), .Y(new_new_n1023_));
  NO4        g1001(.A(new_new_n1023_), .B(new_new_n1006_), .C(new_new_n990_), .D(new_new_n976_), .Y(new_new_n1024_));
  OAI210     g1002(.A0(new_new_n839_), .A1(new_new_n832_), .B0(new_new_n37_), .Y(new_new_n1025_));
  NA3        g1003(.A(new_new_n923_), .B(new_new_n379_), .C(i_5_), .Y(new_new_n1026_));
  NA3        g1004(.A(new_new_n1026_), .B(new_new_n1025_), .C(new_new_n640_), .Y(new_new_n1027_));
  NA2        g1005(.A(new_new_n1027_), .B(new_new_n209_), .Y(new_new_n1028_));
  NA2        g1006(.A(new_new_n189_), .B(new_new_n191_), .Y(new_new_n1029_));
  AO210      g1007(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n1029_), .Y(new_new_n1030_));
  OAI210     g1008(.A0(new_new_n644_), .A1(new_new_n642_), .B0(new_new_n326_), .Y(new_new_n1031_));
  NAi31      g1009(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1032_));
  AOI210     g1010(.A0(new_new_n118_), .A1(new_new_n70_), .B0(new_new_n1032_), .Y(new_new_n1033_));
  NO2        g1011(.A(new_new_n1033_), .B(new_new_n671_), .Y(new_new_n1034_));
  NA3        g1012(.A(new_new_n1034_), .B(new_new_n1031_), .C(new_new_n1030_), .Y(new_new_n1035_));
  NO2        g1013(.A(new_new_n482_), .B(new_new_n275_), .Y(new_new_n1036_));
  NO4        g1014(.A(new_new_n237_), .B(new_new_n146_), .C(new_new_n704_), .D(new_new_n37_), .Y(new_new_n1037_));
  NO2        g1015(.A(new_new_n1037_), .B(new_new_n1036_), .Y(new_new_n1038_));
  OAI210     g1016(.A0(new_new_n1017_), .A1(new_new_n149_), .B0(new_new_n1038_), .Y(new_new_n1039_));
  AOI210     g1017(.A0(new_new_n1035_), .A1(new_new_n49_), .B0(new_new_n1039_), .Y(new_new_n1040_));
  AOI210     g1018(.A0(new_new_n1040_), .A1(new_new_n1028_), .B0(new_new_n73_), .Y(new_new_n1041_));
  NO2        g1019(.A(new_new_n598_), .B(new_new_n390_), .Y(new_new_n1042_));
  NO2        g1020(.A(new_new_n1042_), .B(new_new_n776_), .Y(new_new_n1043_));
  OAI210     g1021(.A0(new_new_n80_), .A1(new_new_n55_), .B0(new_new_n110_), .Y(new_new_n1044_));
  NA2        g1022(.A(new_new_n1044_), .B(new_new_n76_), .Y(new_new_n1045_));
  AOI210     g1023(.A0(new_new_n994_), .A1(new_new_n912_), .B0(new_new_n927_), .Y(new_new_n1046_));
  AOI210     g1024(.A0(new_new_n1046_), .A1(new_new_n1045_), .B0(new_new_n704_), .Y(new_new_n1047_));
  INV        g1025(.A(new_new_n269_), .Y(new_new_n1048_));
  AOI220     g1026(.A0(new_new_n1048_), .A1(new_new_n76_), .B0(new_new_n357_), .B1(new_new_n261_), .Y(new_new_n1049_));
  NO2        g1027(.A(new_new_n1049_), .B(new_new_n241_), .Y(new_new_n1050_));
  NA3        g1028(.A(new_new_n98_), .B(new_new_n315_), .C(new_new_n31_), .Y(new_new_n1051_));
  INV        g1029(.A(new_new_n1051_), .Y(new_new_n1052_));
  NO3        g1030(.A(new_new_n1052_), .B(new_new_n1050_), .C(new_new_n1047_), .Y(new_new_n1053_));
  NA2        g1031(.A(new_new_n159_), .B(new_new_n89_), .Y(new_new_n1054_));
  NA3        g1032(.A(new_new_n780_), .B(new_new_n297_), .C(new_new_n80_), .Y(new_new_n1055_));
  AOI210     g1033(.A0(new_new_n1055_), .A1(new_new_n1054_), .B0(i_11_), .Y(new_new_n1056_));
  NA2        g1034(.A(new_new_n635_), .B(new_new_n218_), .Y(new_new_n1057_));
  OAI210     g1035(.A0(new_new_n1057_), .A1(new_new_n923_), .B0(new_new_n209_), .Y(new_new_n1058_));
  NA2        g1036(.A(new_new_n165_), .B(i_5_), .Y(new_new_n1059_));
  NO2        g1037(.A(new_new_n1058_), .B(new_new_n1059_), .Y(new_new_n1060_));
  NO4        g1038(.A(new_new_n951_), .B(new_new_n499_), .C(new_new_n258_), .D(new_new_n257_), .Y(new_new_n1061_));
  NO2        g1039(.A(new_new_n1061_), .B(new_new_n595_), .Y(new_new_n1062_));
  INV        g1040(.A(new_new_n375_), .Y(new_new_n1063_));
  AOI210     g1041(.A0(new_new_n1063_), .A1(new_new_n1062_), .B0(new_new_n41_), .Y(new_new_n1064_));
  NO3        g1042(.A(new_new_n1064_), .B(new_new_n1060_), .C(new_new_n1056_), .Y(new_new_n1065_));
  OAI210     g1043(.A0(new_new_n1053_), .A1(i_4_), .B0(new_new_n1065_), .Y(new_new_n1066_));
  NO3        g1044(.A(new_new_n1066_), .B(new_new_n1043_), .C(new_new_n1041_), .Y(new_new_n1067_));
  NA4        g1045(.A(new_new_n1067_), .B(new_new_n1024_), .C(new_new_n958_), .D(new_new_n888_), .Y(mai4));
  INV        g1046(.A(new_new_n724_), .Y(new_new_n1071_));
  INV        g1047(.A(i_2_), .Y(new_new_n1072_));
endmodule


