//Benchmark atmr_misex3_1774_0.0156

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1374_, ori_ori_n1378_, ori_ori_n1379_, ori_ori_n1380_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1521_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1533_, mai_mai_n1534_, mai_mai_n1535_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1540_, mai_mai_n1541_, mai_mai_n1542_, mai_mai_n1543_, mai_mai_n1544_, mai_mai_n1545_, mai_mai_n1546_, mai_mai_n1547_, mai_mai_n1548_, mai_mai_n1549_, mai_mai_n1550_, mai_mai_n1551_, mai_mai_n1552_, mai_mai_n1553_, mai_mai_n1555_, mai_mai_n1556_, mai_mai_n1557_, mai_mai_n1558_, mai_mai_n1559_, mai_mai_n1560_, mai_mai_n1561_, mai_mai_n1562_, mai_mai_n1566_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1597_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, men_men_n1605_, men_men_n1606_, men_men_n1608_, men_men_n1609_, men_men_n1610_, men_men_n1611_, men_men_n1612_, men_men_n1613_, men_men_n1614_, men_men_n1615_, men_men_n1619_, men_men_n1620_, men_men_n1621_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  NO2        o0001(.A(d), .B(c), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(o), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(o), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  NO2        o0010(.A(ori_ori_n38_), .B(n), .Y(ori_ori_n39_));
  INV        o0011(.A(h), .Y(ori_ori_n40_));
  NAi21      o0012(.An(j), .B(l), .Y(ori_ori_n41_));
  NAi32      o0013(.An(n), .Bn(o), .C(m), .Y(ori_ori_n42_));
  NO3        o0014(.A(ori_ori_n42_), .B(ori_ori_n41_), .C(ori_ori_n40_), .Y(ori_ori_n43_));
  NAi31      o0015(.An(n), .B(m), .C(l), .Y(ori_ori_n44_));
  INV        o0016(.A(i), .Y(ori_ori_n45_));
  AN2        o0017(.A(h), .B(o), .Y(ori_ori_n46_));
  NA2        o0018(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o0019(.A(ori_ori_n47_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NAi21      o0020(.An(n), .B(m), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(l), .Y(ori_ori_n50_));
  NOi32      o0022(.An(k), .Bn(h), .C(o), .Y(ori_ori_n51_));
  INV        o0023(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NO2        o0024(.A(ori_ori_n52_), .B(ori_ori_n49_), .Y(ori_ori_n53_));
  NO4        o0025(.A(ori_ori_n53_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n54_));
  AOI210     o0026(.A0(ori_ori_n54_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n55_));
  INV        o0027(.A(c), .Y(ori_ori_n56_));
  NA2        o0028(.A(e), .B(b), .Y(ori_ori_n57_));
  NO2        o0029(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0030(.A(d), .Y(ori_ori_n59_));
  NAi21      o0031(.An(i), .B(h), .Y(ori_ori_n60_));
  NAi41      o0032(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n61_));
  NA2        o0033(.A(o), .B(f), .Y(ori_ori_n62_));
  NO2        o0034(.A(ori_ori_n62_), .B(ori_ori_n61_), .Y(ori_ori_n63_));
  NAi21      o0035(.An(i), .B(j), .Y(ori_ori_n64_));
  NAi32      o0036(.An(n), .Bn(k), .C(m), .Y(ori_ori_n65_));
  NAi31      o0037(.An(l), .B(m), .C(k), .Y(ori_ori_n66_));
  NAi21      o0038(.An(e), .B(h), .Y(ori_ori_n67_));
  NAi41      o0039(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n68_));
  INV        o0040(.A(m), .Y(ori_ori_n69_));
  NOi21      o0041(.An(k), .B(l), .Y(ori_ori_n70_));
  NA2        o0042(.A(ori_ori_n70_), .B(ori_ori_n69_), .Y(ori_ori_n71_));
  AN4        o0043(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n72_));
  NOi31      o0044(.An(h), .B(o), .C(f), .Y(ori_ori_n73_));
  NA2        o0045(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  NAi32      o0046(.An(m), .Bn(k), .C(j), .Y(ori_ori_n75_));
  NOi32      o0047(.An(h), .Bn(o), .C(f), .Y(ori_ori_n76_));
  NA2        o0048(.A(ori_ori_n76_), .B(ori_ori_n72_), .Y(ori_ori_n77_));
  OA220      o0049(.A0(ori_ori_n77_), .A1(ori_ori_n75_), .B0(ori_ori_n74_), .B1(ori_ori_n71_), .Y(ori_ori_n78_));
  INV        o0050(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  INV        o0051(.A(n), .Y(ori_ori_n80_));
  NOi32      o0052(.An(e), .Bn(b), .C(d), .Y(ori_ori_n81_));
  NA2        o0053(.A(ori_ori_n81_), .B(ori_ori_n80_), .Y(ori_ori_n82_));
  INV        o0054(.A(j), .Y(ori_ori_n83_));
  AN3        o0055(.A(m), .B(k), .C(i), .Y(ori_ori_n84_));
  NA3        o0056(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(o), .Y(ori_ori_n85_));
  NO2        o0057(.A(ori_ori_n85_), .B(f), .Y(ori_ori_n86_));
  NAi32      o0058(.An(o), .Bn(f), .C(h), .Y(ori_ori_n87_));
  NAi31      o0059(.An(j), .B(m), .C(l), .Y(ori_ori_n88_));
  NO2        o0060(.A(ori_ori_n88_), .B(ori_ori_n87_), .Y(ori_ori_n89_));
  NA2        o0061(.A(m), .B(l), .Y(ori_ori_n90_));
  NAi31      o0062(.An(k), .B(j), .C(o), .Y(ori_ori_n91_));
  NO3        o0063(.A(ori_ori_n91_), .B(ori_ori_n90_), .C(f), .Y(ori_ori_n92_));
  AN2        o0064(.A(j), .B(o), .Y(ori_ori_n93_));
  NOi32      o0065(.An(m), .Bn(l), .C(i), .Y(ori_ori_n94_));
  NOi21      o0066(.An(o), .B(i), .Y(ori_ori_n95_));
  NOi32      o0067(.An(m), .Bn(j), .C(k), .Y(ori_ori_n96_));
  AOI220     o0068(.A0(ori_ori_n96_), .A1(ori_ori_n95_), .B0(ori_ori_n94_), .B1(ori_ori_n93_), .Y(ori_ori_n97_));
  NO2        o0069(.A(ori_ori_n97_), .B(f), .Y(ori_ori_n98_));
  NO4        o0070(.A(ori_ori_n98_), .B(ori_ori_n92_), .C(ori_ori_n89_), .D(ori_ori_n86_), .Y(ori_ori_n99_));
  NAi41      o0071(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n100_));
  AN2        o0072(.A(e), .B(b), .Y(ori_ori_n101_));
  NOi31      o0073(.An(c), .B(h), .C(f), .Y(ori_ori_n102_));
  NA2        o0074(.A(ori_ori_n102_), .B(ori_ori_n101_), .Y(ori_ori_n103_));
  NO3        o0075(.A(ori_ori_n103_), .B(ori_ori_n100_), .C(o), .Y(ori_ori_n104_));
  NOi21      o0076(.An(o), .B(f), .Y(ori_ori_n105_));
  NOi21      o0077(.An(i), .B(h), .Y(ori_ori_n106_));
  INV        o0078(.A(a), .Y(ori_ori_n107_));
  NA2        o0079(.A(ori_ori_n101_), .B(ori_ori_n107_), .Y(ori_ori_n108_));
  INV        o0080(.A(l), .Y(ori_ori_n109_));
  NOi21      o0081(.An(m), .B(n), .Y(ori_ori_n110_));
  AN2        o0082(.A(k), .B(h), .Y(ori_ori_n111_));
  INV        o0083(.A(b), .Y(ori_ori_n112_));
  NA2        o0084(.A(l), .B(j), .Y(ori_ori_n113_));
  AN2        o0085(.A(k), .B(i), .Y(ori_ori_n114_));
  NA2        o0086(.A(ori_ori_n114_), .B(ori_ori_n113_), .Y(ori_ori_n115_));
  NA2        o0087(.A(o), .B(e), .Y(ori_ori_n116_));
  NOi32      o0088(.An(c), .Bn(a), .C(d), .Y(ori_ori_n117_));
  NA2        o0089(.A(ori_ori_n117_), .B(ori_ori_n110_), .Y(ori_ori_n118_));
  INV        o0090(.A(ori_ori_n104_), .Y(ori_ori_n119_));
  OAI210     o0091(.A0(ori_ori_n99_), .A1(ori_ori_n82_), .B0(ori_ori_n119_), .Y(ori_ori_n120_));
  NOi31      o0092(.An(k), .B(m), .C(j), .Y(ori_ori_n121_));
  NA3        o0093(.A(ori_ori_n121_), .B(ori_ori_n73_), .C(ori_ori_n72_), .Y(ori_ori_n122_));
  NOi31      o0094(.An(k), .B(m), .C(i), .Y(ori_ori_n123_));
  NA3        o0095(.A(ori_ori_n123_), .B(ori_ori_n76_), .C(ori_ori_n72_), .Y(ori_ori_n124_));
  NA2        o0096(.A(ori_ori_n124_), .B(ori_ori_n122_), .Y(ori_ori_n125_));
  NOi32      o0097(.An(f), .Bn(b), .C(e), .Y(ori_ori_n126_));
  NAi21      o0098(.An(o), .B(h), .Y(ori_ori_n127_));
  NAi21      o0099(.An(m), .B(n), .Y(ori_ori_n128_));
  NAi21      o0100(.An(j), .B(k), .Y(ori_ori_n129_));
  NO3        o0101(.A(ori_ori_n129_), .B(ori_ori_n128_), .C(ori_ori_n127_), .Y(ori_ori_n130_));
  NAi41      o0102(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n131_));
  NAi31      o0103(.An(j), .B(k), .C(h), .Y(ori_ori_n132_));
  NA2        o0104(.A(ori_ori_n130_), .B(ori_ori_n126_), .Y(ori_ori_n133_));
  NO2        o0105(.A(k), .B(j), .Y(ori_ori_n134_));
  NO2        o0106(.A(ori_ori_n134_), .B(ori_ori_n128_), .Y(ori_ori_n135_));
  AN2        o0107(.A(k), .B(j), .Y(ori_ori_n136_));
  NAi21      o0108(.An(c), .B(b), .Y(ori_ori_n137_));
  NA2        o0109(.A(f), .B(d), .Y(ori_ori_n138_));
  NO4        o0110(.A(ori_ori_n138_), .B(ori_ori_n137_), .C(ori_ori_n136_), .D(ori_ori_n127_), .Y(ori_ori_n139_));
  NA2        o0111(.A(h), .B(c), .Y(ori_ori_n140_));
  NAi31      o0112(.An(f), .B(e), .C(b), .Y(ori_ori_n141_));
  NA2        o0113(.A(ori_ori_n139_), .B(ori_ori_n135_), .Y(ori_ori_n142_));
  NA2        o0114(.A(d), .B(b), .Y(ori_ori_n143_));
  NAi21      o0115(.An(e), .B(f), .Y(ori_ori_n144_));
  NO2        o0116(.A(ori_ori_n144_), .B(ori_ori_n143_), .Y(ori_ori_n145_));
  NA2        o0117(.A(b), .B(a), .Y(ori_ori_n146_));
  NAi21      o0118(.An(e), .B(o), .Y(ori_ori_n147_));
  NAi21      o0119(.An(c), .B(d), .Y(ori_ori_n148_));
  NAi31      o0120(.An(l), .B(k), .C(h), .Y(ori_ori_n149_));
  NO2        o0121(.A(ori_ori_n128_), .B(ori_ori_n149_), .Y(ori_ori_n150_));
  NA2        o0122(.A(ori_ori_n150_), .B(ori_ori_n145_), .Y(ori_ori_n151_));
  NAi41      o0123(.An(ori_ori_n125_), .B(ori_ori_n151_), .C(ori_ori_n142_), .D(ori_ori_n133_), .Y(ori_ori_n152_));
  NAi31      o0124(.An(e), .B(f), .C(b), .Y(ori_ori_n153_));
  NOi21      o0125(.An(o), .B(d), .Y(ori_ori_n154_));
  NO2        o0126(.A(ori_ori_n154_), .B(ori_ori_n153_), .Y(ori_ori_n155_));
  NOi21      o0127(.An(h), .B(i), .Y(ori_ori_n156_));
  NOi21      o0128(.An(k), .B(m), .Y(ori_ori_n157_));
  NA3        o0129(.A(ori_ori_n157_), .B(ori_ori_n156_), .C(n), .Y(ori_ori_n158_));
  NOi21      o0130(.An(ori_ori_n155_), .B(ori_ori_n158_), .Y(ori_ori_n159_));
  NOi21      o0131(.An(h), .B(o), .Y(ori_ori_n160_));
  NO2        o0132(.A(ori_ori_n138_), .B(ori_ori_n137_), .Y(ori_ori_n161_));
  NAi31      o0133(.An(l), .B(j), .C(h), .Y(ori_ori_n162_));
  NO2        o0134(.A(ori_ori_n162_), .B(ori_ori_n49_), .Y(ori_ori_n163_));
  NA2        o0135(.A(ori_ori_n163_), .B(ori_ori_n63_), .Y(ori_ori_n164_));
  NOi32      o0136(.An(n), .Bn(k), .C(m), .Y(ori_ori_n165_));
  NA2        o0137(.A(l), .B(i), .Y(ori_ori_n166_));
  INV        o0138(.A(ori_ori_n164_), .Y(ori_ori_n167_));
  NAi31      o0139(.An(d), .B(f), .C(c), .Y(ori_ori_n168_));
  NAi31      o0140(.An(e), .B(f), .C(c), .Y(ori_ori_n169_));
  NA2        o0141(.A(ori_ori_n169_), .B(ori_ori_n168_), .Y(ori_ori_n170_));
  NA2        o0142(.A(j), .B(h), .Y(ori_ori_n171_));
  OR3        o0143(.A(n), .B(m), .C(k), .Y(ori_ori_n172_));
  NO2        o0144(.A(ori_ori_n172_), .B(ori_ori_n171_), .Y(ori_ori_n173_));
  NAi32      o0145(.An(m), .Bn(k), .C(n), .Y(ori_ori_n174_));
  NO2        o0146(.A(ori_ori_n174_), .B(ori_ori_n171_), .Y(ori_ori_n175_));
  AOI220     o0147(.A0(ori_ori_n175_), .A1(ori_ori_n155_), .B0(ori_ori_n173_), .B1(ori_ori_n170_), .Y(ori_ori_n176_));
  NO2        o0148(.A(n), .B(m), .Y(ori_ori_n177_));
  NA2        o0149(.A(ori_ori_n177_), .B(ori_ori_n50_), .Y(ori_ori_n178_));
  NAi21      o0150(.An(f), .B(e), .Y(ori_ori_n179_));
  NA2        o0151(.A(d), .B(c), .Y(ori_ori_n180_));
  NO2        o0152(.A(ori_ori_n180_), .B(ori_ori_n179_), .Y(ori_ori_n181_));
  NOi21      o0153(.An(ori_ori_n181_), .B(ori_ori_n178_), .Y(ori_ori_n182_));
  NAi31      o0154(.An(m), .B(n), .C(b), .Y(ori_ori_n183_));
  NA2        o0155(.A(k), .B(i), .Y(ori_ori_n184_));
  NAi21      o0156(.An(h), .B(f), .Y(ori_ori_n185_));
  NO2        o0157(.A(ori_ori_n185_), .B(ori_ori_n184_), .Y(ori_ori_n186_));
  NO2        o0158(.A(ori_ori_n183_), .B(ori_ori_n148_), .Y(ori_ori_n187_));
  NA2        o0159(.A(ori_ori_n187_), .B(ori_ori_n186_), .Y(ori_ori_n188_));
  NOi32      o0160(.An(f), .Bn(c), .C(d), .Y(ori_ori_n189_));
  NOi32      o0161(.An(f), .Bn(c), .C(e), .Y(ori_ori_n190_));
  NO2        o0162(.A(ori_ori_n190_), .B(ori_ori_n189_), .Y(ori_ori_n191_));
  NO3        o0163(.A(n), .B(m), .C(j), .Y(ori_ori_n192_));
  NA2        o0164(.A(ori_ori_n192_), .B(ori_ori_n111_), .Y(ori_ori_n193_));
  AO210      o0165(.A0(ori_ori_n193_), .A1(ori_ori_n178_), .B0(ori_ori_n191_), .Y(ori_ori_n194_));
  NAi41      o0166(.An(ori_ori_n182_), .B(ori_ori_n194_), .C(ori_ori_n188_), .D(ori_ori_n176_), .Y(ori_ori_n195_));
  OR4        o0167(.A(ori_ori_n195_), .B(ori_ori_n167_), .C(ori_ori_n159_), .D(ori_ori_n152_), .Y(ori_ori_n196_));
  NO4        o0168(.A(ori_ori_n196_), .B(ori_ori_n120_), .C(ori_ori_n79_), .D(ori_ori_n55_), .Y(ori_ori_n197_));
  NA3        o0169(.A(m), .B(ori_ori_n109_), .C(j), .Y(ori_ori_n198_));
  NAi31      o0170(.An(n), .B(h), .C(o), .Y(ori_ori_n199_));
  NO2        o0171(.A(ori_ori_n199_), .B(ori_ori_n198_), .Y(ori_ori_n200_));
  NOi32      o0172(.An(m), .Bn(k), .C(l), .Y(ori_ori_n201_));
  NA3        o0173(.A(ori_ori_n201_), .B(ori_ori_n83_), .C(o), .Y(ori_ori_n202_));
  NO2        o0174(.A(ori_ori_n202_), .B(n), .Y(ori_ori_n203_));
  NOi21      o0175(.An(k), .B(j), .Y(ori_ori_n204_));
  NA4        o0176(.A(ori_ori_n204_), .B(ori_ori_n110_), .C(i), .D(o), .Y(ori_ori_n205_));
  AN2        o0177(.A(i), .B(o), .Y(ori_ori_n206_));
  NA3        o0178(.A(ori_ori_n70_), .B(ori_ori_n206_), .C(ori_ori_n110_), .Y(ori_ori_n207_));
  NA2        o0179(.A(ori_ori_n207_), .B(ori_ori_n205_), .Y(ori_ori_n208_));
  NO3        o0180(.A(ori_ori_n208_), .B(ori_ori_n203_), .C(ori_ori_n200_), .Y(ori_ori_n209_));
  NAi41      o0181(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n210_));
  INV        o0182(.A(ori_ori_n210_), .Y(ori_ori_n211_));
  INV        o0183(.A(f), .Y(ori_ori_n212_));
  INV        o0184(.A(o), .Y(ori_ori_n213_));
  NOi31      o0185(.An(i), .B(j), .C(h), .Y(ori_ori_n214_));
  NOi21      o0186(.An(l), .B(m), .Y(ori_ori_n215_));
  NA2        o0187(.A(ori_ori_n215_), .B(ori_ori_n214_), .Y(ori_ori_n216_));
  NO3        o0188(.A(ori_ori_n216_), .B(ori_ori_n213_), .C(ori_ori_n212_), .Y(ori_ori_n217_));
  NA2        o0189(.A(ori_ori_n217_), .B(ori_ori_n211_), .Y(ori_ori_n218_));
  OAI210     o0190(.A0(ori_ori_n209_), .A1(ori_ori_n32_), .B0(ori_ori_n218_), .Y(ori_ori_n219_));
  NOi21      o0191(.An(n), .B(m), .Y(ori_ori_n220_));
  NOi32      o0192(.An(l), .Bn(i), .C(j), .Y(ori_ori_n221_));
  NA2        o0193(.A(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  OA220      o0194(.A0(ori_ori_n222_), .A1(ori_ori_n103_), .B0(ori_ori_n75_), .B1(ori_ori_n74_), .Y(ori_ori_n223_));
  NAi21      o0195(.An(j), .B(h), .Y(ori_ori_n224_));
  XN2        o0196(.A(i), .B(h), .Y(ori_ori_n225_));
  NA2        o0197(.A(ori_ori_n225_), .B(ori_ori_n224_), .Y(ori_ori_n226_));
  NOi31      o0198(.An(k), .B(n), .C(m), .Y(ori_ori_n227_));
  NOi31      o0199(.An(ori_ori_n227_), .B(ori_ori_n180_), .C(ori_ori_n179_), .Y(ori_ori_n228_));
  NA2        o0200(.A(ori_ori_n228_), .B(ori_ori_n226_), .Y(ori_ori_n229_));
  NAi31      o0201(.An(f), .B(e), .C(c), .Y(ori_ori_n230_));
  NO4        o0202(.A(ori_ori_n230_), .B(ori_ori_n172_), .C(ori_ori_n171_), .D(ori_ori_n59_), .Y(ori_ori_n231_));
  NA4        o0203(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n232_));
  NAi32      o0204(.An(m), .Bn(i), .C(k), .Y(ori_ori_n233_));
  NA2        o0205(.A(k), .B(h), .Y(ori_ori_n234_));
  INV        o0206(.A(ori_ori_n231_), .Y(ori_ori_n235_));
  NAi21      o0207(.An(n), .B(a), .Y(ori_ori_n236_));
  NO2        o0208(.A(ori_ori_n236_), .B(ori_ori_n143_), .Y(ori_ori_n237_));
  NAi41      o0209(.An(o), .B(m), .C(k), .D(h), .Y(ori_ori_n238_));
  NO2        o0210(.A(ori_ori_n238_), .B(e), .Y(ori_ori_n239_));
  NA2        o0211(.A(ori_ori_n239_), .B(ori_ori_n237_), .Y(ori_ori_n240_));
  AN4        o0212(.A(ori_ori_n240_), .B(ori_ori_n235_), .C(ori_ori_n229_), .D(ori_ori_n223_), .Y(ori_ori_n241_));
  OR2        o0213(.A(h), .B(o), .Y(ori_ori_n242_));
  NO2        o0214(.A(ori_ori_n242_), .B(ori_ori_n100_), .Y(ori_ori_n243_));
  NA2        o0215(.A(ori_ori_n243_), .B(ori_ori_n126_), .Y(ori_ori_n244_));
  NAi41      o0216(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n245_));
  NO2        o0217(.A(ori_ori_n245_), .B(ori_ori_n212_), .Y(ori_ori_n246_));
  NA2        o0218(.A(ori_ori_n157_), .B(ori_ori_n106_), .Y(ori_ori_n247_));
  NAi21      o0219(.An(ori_ori_n247_), .B(ori_ori_n246_), .Y(ori_ori_n248_));
  NO2        o0220(.A(n), .B(a), .Y(ori_ori_n249_));
  NAi31      o0221(.An(ori_ori_n238_), .B(ori_ori_n249_), .C(ori_ori_n101_), .Y(ori_ori_n250_));
  AN2        o0222(.A(ori_ori_n250_), .B(ori_ori_n248_), .Y(ori_ori_n251_));
  NAi21      o0223(.An(h), .B(i), .Y(ori_ori_n252_));
  NA2        o0224(.A(ori_ori_n177_), .B(k), .Y(ori_ori_n253_));
  NO2        o0225(.A(ori_ori_n253_), .B(ori_ori_n252_), .Y(ori_ori_n254_));
  NA2        o0226(.A(ori_ori_n254_), .B(ori_ori_n189_), .Y(ori_ori_n255_));
  NA3        o0227(.A(ori_ori_n255_), .B(ori_ori_n251_), .C(ori_ori_n244_), .Y(ori_ori_n256_));
  NOi21      o0228(.An(o), .B(e), .Y(ori_ori_n257_));
  NO2        o0229(.A(ori_ori_n68_), .B(ori_ori_n69_), .Y(ori_ori_n258_));
  NA2        o0230(.A(ori_ori_n258_), .B(ori_ori_n257_), .Y(ori_ori_n259_));
  NOi32      o0231(.An(l), .Bn(j), .C(i), .Y(ori_ori_n260_));
  AOI210     o0232(.A0(ori_ori_n70_), .A1(ori_ori_n83_), .B0(ori_ori_n260_), .Y(ori_ori_n261_));
  NAi21      o0233(.An(f), .B(o), .Y(ori_ori_n262_));
  NO2        o0234(.A(ori_ori_n262_), .B(ori_ori_n61_), .Y(ori_ori_n263_));
  NO2        o0235(.A(ori_ori_n261_), .B(ori_ori_n259_), .Y(ori_ori_n264_));
  NOi41      o0236(.An(ori_ori_n241_), .B(ori_ori_n264_), .C(ori_ori_n256_), .D(ori_ori_n219_), .Y(ori_ori_n265_));
  NO4        o0237(.A(ori_ori_n200_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n266_));
  NO2        o0238(.A(ori_ori_n266_), .B(ori_ori_n108_), .Y(ori_ori_n267_));
  NA3        o0239(.A(ori_ori_n59_), .B(c), .C(b), .Y(ori_ori_n268_));
  NAi21      o0240(.An(h), .B(o), .Y(ori_ori_n269_));
  NO2        o0241(.A(ori_ori_n247_), .B(ori_ori_n262_), .Y(ori_ori_n270_));
  NA2        o0242(.A(ori_ori_n270_), .B(ori_ori_n72_), .Y(ori_ori_n271_));
  NAi31      o0243(.An(o), .B(k), .C(h), .Y(ori_ori_n272_));
  NO3        o0244(.A(ori_ori_n128_), .B(ori_ori_n272_), .C(l), .Y(ori_ori_n273_));
  NAi31      o0245(.An(e), .B(d), .C(a), .Y(ori_ori_n274_));
  NA2        o0246(.A(ori_ori_n273_), .B(ori_ori_n126_), .Y(ori_ori_n275_));
  NA2        o0247(.A(ori_ori_n275_), .B(ori_ori_n271_), .Y(ori_ori_n276_));
  NA4        o0248(.A(ori_ori_n157_), .B(ori_ori_n76_), .C(ori_ori_n72_), .D(ori_ori_n113_), .Y(ori_ori_n277_));
  NA3        o0249(.A(ori_ori_n157_), .B(ori_ori_n156_), .C(ori_ori_n80_), .Y(ori_ori_n278_));
  NO2        o0250(.A(ori_ori_n278_), .B(ori_ori_n191_), .Y(ori_ori_n279_));
  NOi21      o0251(.An(ori_ori_n277_), .B(ori_ori_n279_), .Y(ori_ori_n280_));
  NA3        o0252(.A(e), .B(c), .C(b), .Y(ori_ori_n281_));
  NAi32      o0253(.An(k), .Bn(i), .C(j), .Y(ori_ori_n282_));
  NAi31      o0254(.An(h), .B(l), .C(i), .Y(ori_ori_n283_));
  NA3        o0255(.A(ori_ori_n283_), .B(ori_ori_n282_), .C(ori_ori_n162_), .Y(ori_ori_n284_));
  NOi21      o0256(.An(ori_ori_n284_), .B(ori_ori_n49_), .Y(ori_ori_n285_));
  NA2        o0257(.A(ori_ori_n263_), .B(ori_ori_n285_), .Y(ori_ori_n286_));
  NAi21      o0258(.An(l), .B(k), .Y(ori_ori_n287_));
  NO2        o0259(.A(ori_ori_n287_), .B(ori_ori_n49_), .Y(ori_ori_n288_));
  NOi21      o0260(.An(l), .B(j), .Y(ori_ori_n289_));
  NA2        o0261(.A(ori_ori_n160_), .B(ori_ori_n289_), .Y(ori_ori_n290_));
  NA3        o0262(.A(ori_ori_n114_), .B(ori_ori_n113_), .C(o), .Y(ori_ori_n291_));
  OR3        o0263(.A(ori_ori_n68_), .B(ori_ori_n69_), .C(e), .Y(ori_ori_n292_));
  AOI210     o0264(.A0(ori_ori_n291_), .A1(ori_ori_n290_), .B0(ori_ori_n292_), .Y(ori_ori_n293_));
  INV        o0265(.A(ori_ori_n293_), .Y(ori_ori_n294_));
  NAi32      o0266(.An(j), .Bn(h), .C(i), .Y(ori_ori_n295_));
  NAi21      o0267(.An(m), .B(l), .Y(ori_ori_n296_));
  NO3        o0268(.A(ori_ori_n296_), .B(ori_ori_n295_), .C(ori_ori_n80_), .Y(ori_ori_n297_));
  NA2        o0269(.A(h), .B(o), .Y(ori_ori_n298_));
  NA2        o0270(.A(ori_ori_n165_), .B(ori_ori_n45_), .Y(ori_ori_n299_));
  NO2        o0271(.A(ori_ori_n299_), .B(ori_ori_n298_), .Y(ori_ori_n300_));
  OAI210     o0272(.A0(ori_ori_n300_), .A1(ori_ori_n297_), .B0(ori_ori_n161_), .Y(ori_ori_n301_));
  NA4        o0273(.A(ori_ori_n301_), .B(ori_ori_n294_), .C(ori_ori_n286_), .D(ori_ori_n280_), .Y(ori_ori_n302_));
  NO2        o0274(.A(ori_ori_n141_), .B(d), .Y(ori_ori_n303_));
  NA2        o0275(.A(ori_ori_n303_), .B(ori_ori_n53_), .Y(ori_ori_n304_));
  NO2        o0276(.A(ori_ori_n103_), .B(ori_ori_n100_), .Y(ori_ori_n305_));
  NAi32      o0277(.An(n), .Bn(m), .C(l), .Y(ori_ori_n306_));
  NO2        o0278(.A(ori_ori_n306_), .B(ori_ori_n295_), .Y(ori_ori_n307_));
  NA2        o0279(.A(ori_ori_n307_), .B(ori_ori_n181_), .Y(ori_ori_n308_));
  NAi31      o0280(.An(k), .B(l), .C(j), .Y(ori_ori_n309_));
  OAI210     o0281(.A0(ori_ori_n287_), .A1(j), .B0(ori_ori_n309_), .Y(ori_ori_n310_));
  NOi21      o0282(.An(ori_ori_n310_), .B(ori_ori_n116_), .Y(ori_ori_n311_));
  NA2        o0283(.A(ori_ori_n308_), .B(ori_ori_n304_), .Y(ori_ori_n312_));
  NO4        o0284(.A(ori_ori_n312_), .B(ori_ori_n302_), .C(ori_ori_n276_), .D(ori_ori_n267_), .Y(ori_ori_n313_));
  NA2        o0285(.A(ori_ori_n254_), .B(ori_ori_n190_), .Y(ori_ori_n314_));
  NAi21      o0286(.An(m), .B(k), .Y(ori_ori_n315_));
  NO2        o0287(.A(ori_ori_n225_), .B(ori_ori_n315_), .Y(ori_ori_n316_));
  NAi41      o0288(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n317_));
  NO2        o0289(.A(ori_ori_n317_), .B(ori_ori_n147_), .Y(ori_ori_n318_));
  NA2        o0290(.A(ori_ori_n318_), .B(ori_ori_n316_), .Y(ori_ori_n319_));
  NAi31      o0291(.An(i), .B(l), .C(h), .Y(ori_ori_n320_));
  NO4        o0292(.A(ori_ori_n320_), .B(ori_ori_n147_), .C(ori_ori_n68_), .D(ori_ori_n69_), .Y(ori_ori_n321_));
  NA2        o0293(.A(e), .B(c), .Y(ori_ori_n322_));
  NO3        o0294(.A(ori_ori_n322_), .B(n), .C(d), .Y(ori_ori_n323_));
  NOi21      o0295(.An(f), .B(h), .Y(ori_ori_n324_));
  NA2        o0296(.A(ori_ori_n324_), .B(ori_ori_n114_), .Y(ori_ori_n325_));
  NO2        o0297(.A(ori_ori_n325_), .B(ori_ori_n213_), .Y(ori_ori_n326_));
  NAi31      o0298(.An(d), .B(e), .C(b), .Y(ori_ori_n327_));
  NO2        o0299(.A(ori_ori_n128_), .B(ori_ori_n327_), .Y(ori_ori_n328_));
  NA2        o0300(.A(ori_ori_n328_), .B(ori_ori_n326_), .Y(ori_ori_n329_));
  NAi41      o0301(.An(ori_ori_n321_), .B(ori_ori_n329_), .C(ori_ori_n319_), .D(ori_ori_n314_), .Y(ori_ori_n330_));
  NO4        o0302(.A(ori_ori_n317_), .B(ori_ori_n75_), .C(ori_ori_n67_), .D(ori_ori_n213_), .Y(ori_ori_n331_));
  NA2        o0303(.A(ori_ori_n249_), .B(ori_ori_n101_), .Y(ori_ori_n332_));
  OR2        o0304(.A(ori_ori_n332_), .B(ori_ori_n202_), .Y(ori_ori_n333_));
  NOi31      o0305(.An(l), .B(n), .C(m), .Y(ori_ori_n334_));
  NA2        o0306(.A(ori_ori_n334_), .B(ori_ori_n214_), .Y(ori_ori_n335_));
  NO2        o0307(.A(ori_ori_n335_), .B(ori_ori_n191_), .Y(ori_ori_n336_));
  NAi32      o0308(.An(ori_ori_n336_), .Bn(ori_ori_n331_), .C(ori_ori_n333_), .Y(ori_ori_n337_));
  NAi32      o0309(.An(m), .Bn(j), .C(k), .Y(ori_ori_n338_));
  NAi41      o0310(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n339_));
  OAI210     o0311(.A0(ori_ori_n210_), .A1(ori_ori_n338_), .B0(ori_ori_n339_), .Y(ori_ori_n340_));
  NOi31      o0312(.An(j), .B(m), .C(k), .Y(ori_ori_n341_));
  NO2        o0313(.A(ori_ori_n121_), .B(ori_ori_n341_), .Y(ori_ori_n342_));
  AN3        o0314(.A(h), .B(o), .C(f), .Y(ori_ori_n343_));
  NAi31      o0315(.An(ori_ori_n342_), .B(ori_ori_n343_), .C(ori_ori_n340_), .Y(ori_ori_n344_));
  NOi32      o0316(.An(m), .Bn(j), .C(l), .Y(ori_ori_n345_));
  NO2        o0317(.A(ori_ori_n345_), .B(ori_ori_n94_), .Y(ori_ori_n346_));
  NAi32      o0318(.An(ori_ori_n346_), .Bn(ori_ori_n199_), .C(ori_ori_n303_), .Y(ori_ori_n347_));
  NO2        o0319(.A(ori_ori_n296_), .B(ori_ori_n295_), .Y(ori_ori_n348_));
  NO2        o0320(.A(ori_ori_n216_), .B(o), .Y(ori_ori_n349_));
  NO2        o0321(.A(ori_ori_n153_), .B(ori_ori_n80_), .Y(ori_ori_n350_));
  AOI220     o0322(.A0(ori_ori_n350_), .A1(ori_ori_n349_), .B0(ori_ori_n246_), .B1(ori_ori_n348_), .Y(ori_ori_n351_));
  NA2        o0323(.A(ori_ori_n233_), .B(ori_ori_n75_), .Y(ori_ori_n352_));
  NA3        o0324(.A(ori_ori_n352_), .B(ori_ori_n343_), .C(ori_ori_n211_), .Y(ori_ori_n353_));
  NA4        o0325(.A(ori_ori_n353_), .B(ori_ori_n351_), .C(ori_ori_n347_), .D(ori_ori_n344_), .Y(ori_ori_n354_));
  NA3        o0326(.A(h), .B(o), .C(f), .Y(ori_ori_n355_));
  NO2        o0327(.A(ori_ori_n355_), .B(ori_ori_n71_), .Y(ori_ori_n356_));
  NA2        o0328(.A(ori_ori_n339_), .B(ori_ori_n210_), .Y(ori_ori_n357_));
  NA2        o0329(.A(ori_ori_n160_), .B(e), .Y(ori_ori_n358_));
  NO2        o0330(.A(ori_ori_n358_), .B(ori_ori_n41_), .Y(ori_ori_n359_));
  NA2        o0331(.A(ori_ori_n357_), .B(ori_ori_n356_), .Y(ori_ori_n360_));
  NOi32      o0332(.An(j), .Bn(o), .C(i), .Y(ori_ori_n361_));
  NA3        o0333(.A(ori_ori_n361_), .B(ori_ori_n287_), .C(ori_ori_n110_), .Y(ori_ori_n362_));
  AO210      o0334(.A0(ori_ori_n108_), .A1(ori_ori_n32_), .B0(ori_ori_n362_), .Y(ori_ori_n363_));
  NOi32      o0335(.An(e), .Bn(b), .C(a), .Y(ori_ori_n364_));
  AN2        o0336(.A(l), .B(j), .Y(ori_ori_n365_));
  NO2        o0337(.A(ori_ori_n315_), .B(ori_ori_n365_), .Y(ori_ori_n366_));
  NO3        o0338(.A(ori_ori_n317_), .B(ori_ori_n67_), .C(ori_ori_n213_), .Y(ori_ori_n367_));
  NA3        o0339(.A(ori_ori_n207_), .B(ori_ori_n205_), .C(ori_ori_n35_), .Y(ori_ori_n368_));
  AOI220     o0340(.A0(ori_ori_n368_), .A1(ori_ori_n364_), .B0(ori_ori_n367_), .B1(ori_ori_n366_), .Y(ori_ori_n369_));
  NO2        o0341(.A(ori_ori_n327_), .B(n), .Y(ori_ori_n370_));
  NA2        o0342(.A(ori_ori_n206_), .B(k), .Y(ori_ori_n371_));
  NA3        o0343(.A(m), .B(ori_ori_n109_), .C(ori_ori_n212_), .Y(ori_ori_n372_));
  NA4        o0344(.A(ori_ori_n201_), .B(ori_ori_n83_), .C(o), .D(ori_ori_n212_), .Y(ori_ori_n373_));
  INV        o0345(.A(ori_ori_n373_), .Y(ori_ori_n374_));
  NA2        o0346(.A(ori_ori_n51_), .B(ori_ori_n110_), .Y(ori_ori_n375_));
  NA2        o0347(.A(ori_ori_n374_), .B(ori_ori_n370_), .Y(ori_ori_n376_));
  NA4        o0348(.A(ori_ori_n376_), .B(ori_ori_n369_), .C(ori_ori_n363_), .D(ori_ori_n360_), .Y(ori_ori_n377_));
  NO4        o0349(.A(ori_ori_n377_), .B(ori_ori_n354_), .C(ori_ori_n337_), .D(ori_ori_n330_), .Y(ori_ori_n378_));
  NA4        o0350(.A(ori_ori_n378_), .B(ori_ori_n313_), .C(ori_ori_n265_), .D(ori_ori_n197_), .Y(ori10));
  NA3        o0351(.A(m), .B(k), .C(i), .Y(ori_ori_n380_));
  NO3        o0352(.A(ori_ori_n380_), .B(j), .C(ori_ori_n213_), .Y(ori_ori_n381_));
  NOi21      o0353(.An(e), .B(f), .Y(ori_ori_n382_));
  NO4        o0354(.A(ori_ori_n148_), .B(ori_ori_n382_), .C(n), .D(ori_ori_n107_), .Y(ori_ori_n383_));
  NAi31      o0355(.An(b), .B(f), .C(c), .Y(ori_ori_n384_));
  INV        o0356(.A(ori_ori_n384_), .Y(ori_ori_n385_));
  NOi32      o0357(.An(k), .Bn(h), .C(j), .Y(ori_ori_n386_));
  NA2        o0358(.A(ori_ori_n386_), .B(ori_ori_n220_), .Y(ori_ori_n387_));
  NA2        o0359(.A(ori_ori_n158_), .B(ori_ori_n387_), .Y(ori_ori_n388_));
  AOI220     o0360(.A0(ori_ori_n388_), .A1(ori_ori_n385_), .B0(ori_ori_n383_), .B1(ori_ori_n381_), .Y(ori_ori_n389_));
  AN2        o0361(.A(j), .B(h), .Y(ori_ori_n390_));
  NO3        o0362(.A(n), .B(m), .C(k), .Y(ori_ori_n391_));
  NA2        o0363(.A(ori_ori_n391_), .B(ori_ori_n390_), .Y(ori_ori_n392_));
  NO3        o0364(.A(ori_ori_n392_), .B(ori_ori_n148_), .C(ori_ori_n212_), .Y(ori_ori_n393_));
  OR2        o0365(.A(m), .B(k), .Y(ori_ori_n394_));
  NO2        o0366(.A(ori_ori_n171_), .B(ori_ori_n394_), .Y(ori_ori_n395_));
  NA4        o0367(.A(n), .B(f), .C(c), .D(ori_ori_n112_), .Y(ori_ori_n396_));
  NOi21      o0368(.An(ori_ori_n395_), .B(ori_ori_n396_), .Y(ori_ori_n397_));
  NOi32      o0369(.An(d), .Bn(a), .C(c), .Y(ori_ori_n398_));
  NA2        o0370(.A(ori_ori_n398_), .B(ori_ori_n179_), .Y(ori_ori_n399_));
  NAi21      o0371(.An(i), .B(o), .Y(ori_ori_n400_));
  NAi31      o0372(.An(k), .B(m), .C(j), .Y(ori_ori_n401_));
  NO3        o0373(.A(ori_ori_n401_), .B(ori_ori_n400_), .C(n), .Y(ori_ori_n402_));
  NOi21      o0374(.An(ori_ori_n402_), .B(ori_ori_n399_), .Y(ori_ori_n403_));
  NO3        o0375(.A(ori_ori_n403_), .B(ori_ori_n397_), .C(ori_ori_n393_), .Y(ori_ori_n404_));
  NO2        o0376(.A(ori_ori_n396_), .B(ori_ori_n296_), .Y(ori_ori_n405_));
  NOi32      o0377(.An(f), .Bn(d), .C(c), .Y(ori_ori_n406_));
  AOI220     o0378(.A0(ori_ori_n406_), .A1(ori_ori_n307_), .B0(ori_ori_n405_), .B1(ori_ori_n214_), .Y(ori_ori_n407_));
  NA3        o0379(.A(ori_ori_n407_), .B(ori_ori_n404_), .C(ori_ori_n389_), .Y(ori_ori_n408_));
  NO2        o0380(.A(ori_ori_n59_), .B(ori_ori_n112_), .Y(ori_ori_n409_));
  NA2        o0381(.A(ori_ori_n249_), .B(ori_ori_n409_), .Y(ori_ori_n410_));
  INV        o0382(.A(e), .Y(ori_ori_n411_));
  NA2        o0383(.A(ori_ori_n46_), .B(e), .Y(ori_ori_n412_));
  OAI220     o0384(.A0(ori_ori_n412_), .A1(ori_ori_n198_), .B0(ori_ori_n202_), .B1(ori_ori_n411_), .Y(ori_ori_n413_));
  AN2        o0385(.A(o), .B(e), .Y(ori_ori_n414_));
  NA3        o0386(.A(ori_ori_n414_), .B(ori_ori_n201_), .C(i), .Y(ori_ori_n415_));
  OAI210     o0387(.A0(ori_ori_n85_), .A1(ori_ori_n411_), .B0(ori_ori_n415_), .Y(ori_ori_n416_));
  NO2        o0388(.A(ori_ori_n97_), .B(ori_ori_n411_), .Y(ori_ori_n417_));
  NO3        o0389(.A(ori_ori_n417_), .B(ori_ori_n416_), .C(ori_ori_n413_), .Y(ori_ori_n418_));
  NOi32      o0390(.An(h), .Bn(e), .C(o), .Y(ori_ori_n419_));
  NA3        o0391(.A(ori_ori_n419_), .B(ori_ori_n289_), .C(m), .Y(ori_ori_n420_));
  NOi21      o0392(.An(o), .B(h), .Y(ori_ori_n421_));
  AN3        o0393(.A(m), .B(l), .C(i), .Y(ori_ori_n422_));
  NA3        o0394(.A(ori_ori_n422_), .B(ori_ori_n421_), .C(e), .Y(ori_ori_n423_));
  AN3        o0395(.A(h), .B(o), .C(e), .Y(ori_ori_n424_));
  NA2        o0396(.A(ori_ori_n424_), .B(ori_ori_n94_), .Y(ori_ori_n425_));
  AN3        o0397(.A(ori_ori_n425_), .B(ori_ori_n423_), .C(ori_ori_n420_), .Y(ori_ori_n426_));
  AOI210     o0398(.A0(ori_ori_n426_), .A1(ori_ori_n418_), .B0(ori_ori_n410_), .Y(ori_ori_n427_));
  NA3        o0399(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(e), .Y(ori_ori_n428_));
  NO2        o0400(.A(ori_ori_n428_), .B(ori_ori_n410_), .Y(ori_ori_n429_));
  NA3        o0401(.A(ori_ori_n398_), .B(ori_ori_n179_), .C(ori_ori_n80_), .Y(ori_ori_n430_));
  NAi31      o0402(.An(b), .B(c), .C(a), .Y(ori_ori_n431_));
  NO2        o0403(.A(ori_ori_n431_), .B(n), .Y(ori_ori_n432_));
  NA2        o0404(.A(ori_ori_n51_), .B(m), .Y(ori_ori_n433_));
  NO2        o0405(.A(ori_ori_n433_), .B(ori_ori_n144_), .Y(ori_ori_n434_));
  NA2        o0406(.A(ori_ori_n434_), .B(ori_ori_n432_), .Y(ori_ori_n435_));
  INV        o0407(.A(ori_ori_n435_), .Y(ori_ori_n436_));
  NO4        o0408(.A(ori_ori_n436_), .B(ori_ori_n429_), .C(ori_ori_n427_), .D(ori_ori_n408_), .Y(ori_ori_n437_));
  NA2        o0409(.A(i), .B(o), .Y(ori_ori_n438_));
  NOi21      o0410(.An(a), .B(n), .Y(ori_ori_n439_));
  NOi21      o0411(.An(d), .B(c), .Y(ori_ori_n440_));
  NA2        o0412(.A(ori_ori_n440_), .B(ori_ori_n439_), .Y(ori_ori_n441_));
  NA3        o0413(.A(i), .B(o), .C(f), .Y(ori_ori_n442_));
  OR2        o0414(.A(ori_ori_n442_), .B(ori_ori_n66_), .Y(ori_ori_n443_));
  NA3        o0415(.A(ori_ori_n422_), .B(ori_ori_n421_), .C(ori_ori_n179_), .Y(ori_ori_n444_));
  AOI210     o0416(.A0(ori_ori_n444_), .A1(ori_ori_n443_), .B0(ori_ori_n441_), .Y(ori_ori_n445_));
  INV        o0417(.A(ori_ori_n445_), .Y(ori_ori_n446_));
  OR2        o0418(.A(n), .B(m), .Y(ori_ori_n447_));
  NO2        o0419(.A(ori_ori_n447_), .B(ori_ori_n149_), .Y(ori_ori_n448_));
  NO2        o0420(.A(ori_ori_n180_), .B(ori_ori_n144_), .Y(ori_ori_n449_));
  OAI210     o0421(.A0(ori_ori_n448_), .A1(ori_ori_n173_), .B0(ori_ori_n449_), .Y(ori_ori_n450_));
  INV        o0422(.A(ori_ori_n375_), .Y(ori_ori_n451_));
  NA3        o0423(.A(ori_ori_n451_), .B(ori_ori_n364_), .C(d), .Y(ori_ori_n452_));
  NO2        o0424(.A(ori_ori_n431_), .B(ori_ori_n49_), .Y(ori_ori_n453_));
  NO3        o0425(.A(ori_ori_n62_), .B(ori_ori_n109_), .C(e), .Y(ori_ori_n454_));
  NAi21      o0426(.An(k), .B(j), .Y(ori_ori_n455_));
  NA2        o0427(.A(ori_ori_n252_), .B(ori_ori_n455_), .Y(ori_ori_n456_));
  NA3        o0428(.A(ori_ori_n456_), .B(ori_ori_n454_), .C(ori_ori_n453_), .Y(ori_ori_n457_));
  NAi21      o0429(.An(e), .B(d), .Y(ori_ori_n458_));
  NO2        o0430(.A(ori_ori_n458_), .B(ori_ori_n56_), .Y(ori_ori_n459_));
  NO2        o0431(.A(ori_ori_n253_), .B(ori_ori_n212_), .Y(ori_ori_n460_));
  NA3        o0432(.A(ori_ori_n460_), .B(ori_ori_n459_), .C(ori_ori_n226_), .Y(ori_ori_n461_));
  NA4        o0433(.A(ori_ori_n461_), .B(ori_ori_n457_), .C(ori_ori_n452_), .D(ori_ori_n450_), .Y(ori_ori_n462_));
  NO2        o0434(.A(ori_ori_n335_), .B(ori_ori_n212_), .Y(ori_ori_n463_));
  NA2        o0435(.A(ori_ori_n463_), .B(ori_ori_n459_), .Y(ori_ori_n464_));
  NOi31      o0436(.An(n), .B(m), .C(k), .Y(ori_ori_n465_));
  AOI220     o0437(.A0(ori_ori_n465_), .A1(ori_ori_n390_), .B0(ori_ori_n220_), .B1(ori_ori_n50_), .Y(ori_ori_n466_));
  NAi31      o0438(.An(o), .B(f), .C(c), .Y(ori_ori_n467_));
  OR3        o0439(.A(ori_ori_n467_), .B(ori_ori_n466_), .C(e), .Y(ori_ori_n468_));
  NA3        o0440(.A(ori_ori_n468_), .B(ori_ori_n464_), .C(ori_ori_n308_), .Y(ori_ori_n469_));
  NOi41      o0441(.An(ori_ori_n446_), .B(ori_ori_n469_), .C(ori_ori_n462_), .D(ori_ori_n264_), .Y(ori_ori_n470_));
  NOi32      o0442(.An(c), .Bn(a), .C(b), .Y(ori_ori_n471_));
  NA2        o0443(.A(ori_ori_n471_), .B(ori_ori_n110_), .Y(ori_ori_n472_));
  NA2        o0444(.A(ori_ori_n272_), .B(ori_ori_n149_), .Y(ori_ori_n473_));
  AN2        o0445(.A(e), .B(d), .Y(ori_ori_n474_));
  NA2        o0446(.A(ori_ori_n474_), .B(ori_ori_n473_), .Y(ori_ori_n475_));
  INV        o0447(.A(ori_ori_n144_), .Y(ori_ori_n476_));
  NO2        o0448(.A(ori_ori_n127_), .B(ori_ori_n41_), .Y(ori_ori_n477_));
  NO2        o0449(.A(ori_ori_n62_), .B(e), .Y(ori_ori_n478_));
  NOi31      o0450(.An(j), .B(k), .C(i), .Y(ori_ori_n479_));
  NOi21      o0451(.An(ori_ori_n162_), .B(ori_ori_n479_), .Y(ori_ori_n480_));
  NA4        o0452(.A(ori_ori_n320_), .B(ori_ori_n480_), .C(ori_ori_n261_), .D(ori_ori_n115_), .Y(ori_ori_n481_));
  AOI220     o0453(.A0(ori_ori_n481_), .A1(ori_ori_n478_), .B0(ori_ori_n477_), .B1(ori_ori_n476_), .Y(ori_ori_n482_));
  AOI210     o0454(.A0(ori_ori_n482_), .A1(ori_ori_n475_), .B0(ori_ori_n472_), .Y(ori_ori_n483_));
  NO2        o0455(.A(ori_ori_n208_), .B(ori_ori_n203_), .Y(ori_ori_n484_));
  NOi21      o0456(.An(a), .B(b), .Y(ori_ori_n485_));
  NA3        o0457(.A(e), .B(d), .C(c), .Y(ori_ori_n486_));
  NAi21      o0458(.An(ori_ori_n486_), .B(ori_ori_n485_), .Y(ori_ori_n487_));
  NO2        o0459(.A(ori_ori_n430_), .B(ori_ori_n202_), .Y(ori_ori_n488_));
  NOi21      o0460(.An(ori_ori_n487_), .B(ori_ori_n488_), .Y(ori_ori_n489_));
  AOI210     o0461(.A0(ori_ori_n266_), .A1(ori_ori_n484_), .B0(ori_ori_n489_), .Y(ori_ori_n490_));
  NO4        o0462(.A(ori_ori_n185_), .B(ori_ori_n100_), .C(ori_ori_n56_), .D(b), .Y(ori_ori_n491_));
  NA2        o0463(.A(ori_ori_n385_), .B(ori_ori_n150_), .Y(ori_ori_n492_));
  OR2        o0464(.A(k), .B(j), .Y(ori_ori_n493_));
  NA2        o0465(.A(l), .B(k), .Y(ori_ori_n494_));
  NA3        o0466(.A(ori_ori_n494_), .B(ori_ori_n493_), .C(ori_ori_n220_), .Y(ori_ori_n495_));
  AOI210     o0467(.A0(ori_ori_n233_), .A1(ori_ori_n338_), .B0(ori_ori_n80_), .Y(ori_ori_n496_));
  NOi21      o0468(.An(ori_ori_n495_), .B(ori_ori_n496_), .Y(ori_ori_n497_));
  OR3        o0469(.A(ori_ori_n497_), .B(ori_ori_n140_), .C(ori_ori_n131_), .Y(ori_ori_n498_));
  NA3        o0470(.A(ori_ori_n277_), .B(ori_ori_n124_), .C(ori_ori_n122_), .Y(ori_ori_n499_));
  NO3        o0471(.A(ori_ori_n430_), .B(ori_ori_n88_), .C(ori_ori_n127_), .Y(ori_ori_n500_));
  NO3        o0472(.A(ori_ori_n500_), .B(ori_ori_n499_), .C(ori_ori_n321_), .Y(ori_ori_n501_));
  NA3        o0473(.A(ori_ori_n501_), .B(ori_ori_n498_), .C(ori_ori_n492_), .Y(ori_ori_n502_));
  NO4        o0474(.A(ori_ori_n502_), .B(ori_ori_n491_), .C(ori_ori_n490_), .D(ori_ori_n483_), .Y(ori_ori_n503_));
  NOi21      o0475(.An(d), .B(e), .Y(ori_ori_n504_));
  NO2        o0476(.A(ori_ori_n185_), .B(ori_ori_n56_), .Y(ori_ori_n505_));
  NAi31      o0477(.An(j), .B(l), .C(i), .Y(ori_ori_n506_));
  OAI210     o0478(.A0(ori_ori_n506_), .A1(ori_ori_n128_), .B0(ori_ori_n100_), .Y(ori_ori_n507_));
  NA4        o0479(.A(ori_ori_n507_), .B(ori_ori_n505_), .C(ori_ori_n504_), .D(b), .Y(ori_ori_n508_));
  NO3        o0480(.A(ori_ori_n399_), .B(ori_ori_n346_), .C(ori_ori_n199_), .Y(ori_ori_n509_));
  NO2        o0481(.A(ori_ori_n399_), .B(ori_ori_n375_), .Y(ori_ori_n510_));
  NO4        o0482(.A(ori_ori_n510_), .B(ori_ori_n509_), .C(ori_ori_n182_), .D(ori_ori_n305_), .Y(ori_ori_n511_));
  NA3        o0483(.A(ori_ori_n511_), .B(ori_ori_n508_), .C(ori_ori_n241_), .Y(ori_ori_n512_));
  OAI210     o0484(.A0(ori_ori_n123_), .A1(ori_ori_n121_), .B0(n), .Y(ori_ori_n513_));
  NO2        o0485(.A(ori_ori_n513_), .B(ori_ori_n127_), .Y(ori_ori_n514_));
  OA210      o0486(.A0(ori_ori_n243_), .A1(ori_ori_n514_), .B0(ori_ori_n190_), .Y(ori_ori_n515_));
  XO2        o0487(.A(i), .B(h), .Y(ori_ori_n516_));
  NA3        o0488(.A(ori_ori_n516_), .B(ori_ori_n157_), .C(n), .Y(ori_ori_n517_));
  NAi41      o0489(.An(ori_ori_n297_), .B(ori_ori_n517_), .C(ori_ori_n466_), .D(ori_ori_n387_), .Y(ori_ori_n518_));
  NOi32      o0490(.An(ori_ori_n518_), .Bn(ori_ori_n478_), .C(ori_ori_n268_), .Y(ori_ori_n519_));
  NAi31      o0491(.An(c), .B(f), .C(d), .Y(ori_ori_n520_));
  AOI210     o0492(.A0(ori_ori_n278_), .A1(ori_ori_n193_), .B0(ori_ori_n520_), .Y(ori_ori_n521_));
  NOi21      o0493(.An(ori_ori_n78_), .B(ori_ori_n521_), .Y(ori_ori_n522_));
  NA2        o0494(.A(ori_ori_n227_), .B(ori_ori_n106_), .Y(ori_ori_n523_));
  AOI210     o0495(.A0(ori_ori_n523_), .A1(ori_ori_n178_), .B0(ori_ori_n520_), .Y(ori_ori_n524_));
  AOI210     o0496(.A0(ori_ori_n362_), .A1(ori_ori_n35_), .B0(ori_ori_n487_), .Y(ori_ori_n525_));
  NO2        o0497(.A(ori_ori_n525_), .B(ori_ori_n524_), .Y(ori_ori_n526_));
  AO220      o0498(.A0(ori_ori_n285_), .A1(ori_ori_n263_), .B0(ori_ori_n163_), .B1(ori_ori_n63_), .Y(ori_ori_n527_));
  NA3        o0499(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(f), .Y(ori_ori_n528_));
  INV        o0500(.A(ori_ori_n293_), .Y(ori_ori_n529_));
  NAi41      o0501(.An(ori_ori_n527_), .B(ori_ori_n529_), .C(ori_ori_n526_), .D(ori_ori_n522_), .Y(ori_ori_n530_));
  NO4        o0502(.A(ori_ori_n530_), .B(ori_ori_n519_), .C(ori_ori_n515_), .D(ori_ori_n512_), .Y(ori_ori_n531_));
  NA4        o0503(.A(ori_ori_n531_), .B(ori_ori_n503_), .C(ori_ori_n470_), .D(ori_ori_n437_), .Y(ori11));
  NO2        o0504(.A(ori_ori_n68_), .B(f), .Y(ori_ori_n533_));
  NA2        o0505(.A(j), .B(o), .Y(ori_ori_n534_));
  NAi31      o0506(.An(i), .B(m), .C(l), .Y(ori_ori_n535_));
  NA3        o0507(.A(m), .B(k), .C(j), .Y(ori_ori_n536_));
  OAI220     o0508(.A0(ori_ori_n536_), .A1(ori_ori_n127_), .B0(ori_ori_n535_), .B1(ori_ori_n534_), .Y(ori_ori_n537_));
  NA2        o0509(.A(ori_ori_n537_), .B(ori_ori_n533_), .Y(ori_ori_n538_));
  NOi32      o0510(.An(e), .Bn(b), .C(f), .Y(ori_ori_n539_));
  NA2        o0511(.A(ori_ori_n46_), .B(j), .Y(ori_ori_n540_));
  NO2        o0512(.A(ori_ori_n540_), .B(ori_ori_n299_), .Y(ori_ori_n541_));
  NAi31      o0513(.An(d), .B(e), .C(a), .Y(ori_ori_n542_));
  NO2        o0514(.A(ori_ori_n542_), .B(n), .Y(ori_ori_n543_));
  AOI220     o0515(.A0(ori_ori_n543_), .A1(ori_ori_n98_), .B0(ori_ori_n541_), .B1(ori_ori_n539_), .Y(ori_ori_n544_));
  NA2        o0516(.A(j), .B(i), .Y(ori_ori_n545_));
  NAi31      o0517(.An(n), .B(m), .C(k), .Y(ori_ori_n546_));
  NO3        o0518(.A(ori_ori_n546_), .B(ori_ori_n545_), .C(ori_ori_n109_), .Y(ori_ori_n547_));
  NO4        o0519(.A(n), .B(d), .C(ori_ori_n112_), .D(a), .Y(ori_ori_n548_));
  OR2        o0520(.A(n), .B(c), .Y(ori_ori_n549_));
  NO2        o0521(.A(ori_ori_n549_), .B(ori_ori_n146_), .Y(ori_ori_n550_));
  NO2        o0522(.A(ori_ori_n550_), .B(ori_ori_n548_), .Y(ori_ori_n551_));
  NOi32      o0523(.An(o), .Bn(f), .C(i), .Y(ori_ori_n552_));
  AOI220     o0524(.A0(ori_ori_n552_), .A1(ori_ori_n96_), .B0(ori_ori_n537_), .B1(f), .Y(ori_ori_n553_));
  NO2        o0525(.A(ori_ori_n272_), .B(ori_ori_n49_), .Y(ori_ori_n554_));
  NO2        o0526(.A(ori_ori_n553_), .B(ori_ori_n551_), .Y(ori_ori_n555_));
  INV        o0527(.A(ori_ori_n555_), .Y(ori_ori_n556_));
  NA2        o0528(.A(ori_ori_n136_), .B(ori_ori_n34_), .Y(ori_ori_n557_));
  OAI220     o0529(.A0(ori_ori_n557_), .A1(m), .B0(ori_ori_n540_), .B1(ori_ori_n233_), .Y(ori_ori_n558_));
  NOi41      o0530(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n559_));
  NAi32      o0531(.An(e), .Bn(b), .C(c), .Y(ori_ori_n560_));
  OR2        o0532(.A(ori_ori_n560_), .B(ori_ori_n80_), .Y(ori_ori_n561_));
  AN2        o0533(.A(ori_ori_n339_), .B(ori_ori_n317_), .Y(ori_ori_n562_));
  NA2        o0534(.A(ori_ori_n562_), .B(ori_ori_n561_), .Y(ori_ori_n563_));
  OA210      o0535(.A0(ori_ori_n563_), .A1(ori_ori_n559_), .B0(ori_ori_n558_), .Y(ori_ori_n564_));
  OAI220     o0536(.A0(ori_ori_n401_), .A1(ori_ori_n400_), .B0(ori_ori_n535_), .B1(ori_ori_n534_), .Y(ori_ori_n565_));
  NAi31      o0537(.An(d), .B(c), .C(a), .Y(ori_ori_n566_));
  NO2        o0538(.A(ori_ori_n566_), .B(n), .Y(ori_ori_n567_));
  NO2        o0539(.A(ori_ori_n230_), .B(ori_ori_n107_), .Y(ori_ori_n568_));
  NA2        o0540(.A(ori_ori_n402_), .B(ori_ori_n568_), .Y(ori_ori_n569_));
  INV        o0541(.A(ori_ori_n569_), .Y(ori_ori_n570_));
  NO2        o0542(.A(ori_ori_n274_), .B(n), .Y(ori_ori_n571_));
  NO2        o0543(.A(ori_ori_n432_), .B(ori_ori_n571_), .Y(ori_ori_n572_));
  NA2        o0544(.A(ori_ori_n565_), .B(f), .Y(ori_ori_n573_));
  NAi32      o0545(.An(d), .Bn(a), .C(b), .Y(ori_ori_n574_));
  NO2        o0546(.A(ori_ori_n574_), .B(ori_ori_n49_), .Y(ori_ori_n575_));
  NA2        o0547(.A(h), .B(f), .Y(ori_ori_n576_));
  NO2        o0548(.A(ori_ori_n576_), .B(ori_ori_n91_), .Y(ori_ori_n577_));
  NO3        o0549(.A(ori_ori_n174_), .B(ori_ori_n171_), .C(o), .Y(ori_ori_n578_));
  AOI220     o0550(.A0(ori_ori_n578_), .A1(ori_ori_n58_), .B0(ori_ori_n577_), .B1(ori_ori_n575_), .Y(ori_ori_n579_));
  OAI210     o0551(.A0(ori_ori_n573_), .A1(ori_ori_n572_), .B0(ori_ori_n579_), .Y(ori_ori_n580_));
  AN3        o0552(.A(j), .B(h), .C(o), .Y(ori_ori_n581_));
  NO2        o0553(.A(ori_ori_n143_), .B(c), .Y(ori_ori_n582_));
  NA3        o0554(.A(ori_ori_n582_), .B(ori_ori_n581_), .C(ori_ori_n465_), .Y(ori_ori_n583_));
  NA3        o0555(.A(f), .B(d), .C(b), .Y(ori_ori_n584_));
  NO4        o0556(.A(ori_ori_n584_), .B(ori_ori_n174_), .C(ori_ori_n171_), .D(o), .Y(ori_ori_n585_));
  NAi21      o0557(.An(ori_ori_n585_), .B(ori_ori_n583_), .Y(ori_ori_n586_));
  NO4        o0558(.A(ori_ori_n586_), .B(ori_ori_n580_), .C(ori_ori_n570_), .D(ori_ori_n564_), .Y(ori_ori_n587_));
  AN4        o0559(.A(ori_ori_n587_), .B(ori_ori_n556_), .C(ori_ori_n544_), .D(ori_ori_n538_), .Y(ori_ori_n588_));
  INV        o0560(.A(k), .Y(ori_ori_n589_));
  NA3        o0561(.A(l), .B(ori_ori_n589_), .C(i), .Y(ori_ori_n590_));
  INV        o0562(.A(ori_ori_n590_), .Y(ori_ori_n591_));
  NA4        o0563(.A(ori_ori_n398_), .B(ori_ori_n421_), .C(ori_ori_n179_), .D(ori_ori_n110_), .Y(ori_ori_n592_));
  NAi32      o0564(.An(h), .Bn(f), .C(o), .Y(ori_ori_n593_));
  NAi41      o0565(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n594_));
  OAI210     o0566(.A0(ori_ori_n542_), .A1(n), .B0(ori_ori_n594_), .Y(ori_ori_n595_));
  NA2        o0567(.A(ori_ori_n595_), .B(m), .Y(ori_ori_n596_));
  NAi31      o0568(.An(h), .B(o), .C(f), .Y(ori_ori_n597_));
  OR2        o0569(.A(ori_ori_n596_), .B(ori_ori_n593_), .Y(ori_ori_n598_));
  NO3        o0570(.A(ori_ori_n593_), .B(ori_ori_n68_), .C(ori_ori_n69_), .Y(ori_ori_n599_));
  NO4        o0571(.A(ori_ori_n597_), .B(ori_ori_n549_), .C(ori_ori_n146_), .D(ori_ori_n69_), .Y(ori_ori_n600_));
  OR2        o0572(.A(ori_ori_n600_), .B(ori_ori_n599_), .Y(ori_ori_n601_));
  NAi31      o0573(.An(ori_ori_n601_), .B(ori_ori_n598_), .C(ori_ori_n592_), .Y(ori_ori_n602_));
  NAi31      o0574(.An(f), .B(h), .C(o), .Y(ori_ori_n603_));
  NOi32      o0575(.An(b), .Bn(a), .C(c), .Y(ori_ori_n604_));
  NOi32      o0576(.An(d), .Bn(a), .C(e), .Y(ori_ori_n605_));
  NA2        o0577(.A(ori_ori_n605_), .B(ori_ori_n110_), .Y(ori_ori_n606_));
  NO2        o0578(.A(n), .B(c), .Y(ori_ori_n607_));
  NA3        o0579(.A(ori_ori_n607_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n608_));
  NA2        o0580(.A(ori_ori_n608_), .B(ori_ori_n606_), .Y(ori_ori_n609_));
  NOi32      o0581(.An(e), .Bn(a), .C(d), .Y(ori_ori_n610_));
  AOI210     o0582(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n610_), .Y(ori_ori_n611_));
  AOI210     o0583(.A0(ori_ori_n611_), .A1(ori_ori_n212_), .B0(ori_ori_n557_), .Y(ori_ori_n612_));
  NA2        o0584(.A(ori_ori_n612_), .B(ori_ori_n609_), .Y(ori_ori_n613_));
  OAI210     o0585(.A0(ori_ori_n248_), .A1(ori_ori_n83_), .B0(ori_ori_n613_), .Y(ori_ori_n614_));
  AOI210     o0586(.A0(ori_ori_n602_), .A1(ori_ori_n591_), .B0(ori_ori_n614_), .Y(ori_ori_n615_));
  NO3        o0587(.A(ori_ori_n315_), .B(ori_ori_n60_), .C(n), .Y(ori_ori_n616_));
  NA3        o0588(.A(ori_ori_n520_), .B(ori_ori_n169_), .C(ori_ori_n168_), .Y(ori_ori_n617_));
  NA2        o0589(.A(ori_ori_n467_), .B(ori_ori_n230_), .Y(ori_ori_n618_));
  OR2        o0590(.A(ori_ori_n618_), .B(ori_ori_n617_), .Y(ori_ori_n619_));
  NA2        o0591(.A(ori_ori_n70_), .B(ori_ori_n110_), .Y(ori_ori_n620_));
  NA2        o0592(.A(ori_ori_n619_), .B(ori_ori_n616_), .Y(ori_ori_n621_));
  NO2        o0593(.A(ori_ori_n621_), .B(ori_ori_n83_), .Y(ori_ori_n622_));
  NA3        o0594(.A(ori_ori_n559_), .B(ori_ori_n341_), .C(ori_ori_n46_), .Y(ori_ori_n623_));
  NOi32      o0595(.An(e), .Bn(c), .C(f), .Y(ori_ori_n624_));
  NOi21      o0596(.An(f), .B(o), .Y(ori_ori_n625_));
  NO2        o0597(.A(ori_ori_n625_), .B(ori_ori_n210_), .Y(ori_ori_n626_));
  AOI220     o0598(.A0(ori_ori_n626_), .A1(ori_ori_n395_), .B0(ori_ori_n624_), .B1(ori_ori_n173_), .Y(ori_ori_n627_));
  NA3        o0599(.A(ori_ori_n627_), .B(ori_ori_n623_), .C(ori_ori_n176_), .Y(ori_ori_n628_));
  NOi21      o0600(.An(j), .B(l), .Y(ori_ori_n629_));
  NAi21      o0601(.An(k), .B(h), .Y(ori_ori_n630_));
  NO2        o0602(.A(ori_ori_n630_), .B(ori_ori_n262_), .Y(ori_ori_n631_));
  NA2        o0603(.A(ori_ori_n631_), .B(ori_ori_n629_), .Y(ori_ori_n632_));
  OR2        o0604(.A(ori_ori_n632_), .B(ori_ori_n596_), .Y(ori_ori_n633_));
  NOi31      o0605(.An(m), .B(n), .C(k), .Y(ori_ori_n634_));
  NA2        o0606(.A(ori_ori_n629_), .B(ori_ori_n634_), .Y(ori_ori_n635_));
  NO2        o0607(.A(ori_ori_n274_), .B(ori_ori_n49_), .Y(ori_ori_n636_));
  NO2        o0608(.A(ori_ori_n309_), .B(ori_ori_n603_), .Y(ori_ori_n637_));
  NO2        o0609(.A(ori_ori_n542_), .B(ori_ori_n49_), .Y(ori_ori_n638_));
  AOI220     o0610(.A0(ori_ori_n638_), .A1(ori_ori_n637_), .B0(ori_ori_n636_), .B1(ori_ori_n577_), .Y(ori_ori_n639_));
  NA2        o0611(.A(ori_ori_n639_), .B(ori_ori_n633_), .Y(ori_ori_n640_));
  NA2        o0612(.A(ori_ori_n106_), .B(ori_ori_n36_), .Y(ori_ori_n641_));
  NO2        o0613(.A(k), .B(ori_ori_n213_), .Y(ori_ori_n642_));
  INV        o0614(.A(ori_ori_n364_), .Y(ori_ori_n643_));
  NO2        o0615(.A(ori_ori_n643_), .B(n), .Y(ori_ori_n644_));
  NAi31      o0616(.An(ori_ori_n641_), .B(ori_ori_n644_), .C(ori_ori_n642_), .Y(ori_ori_n645_));
  NO2        o0617(.A(ori_ori_n540_), .B(ori_ori_n174_), .Y(ori_ori_n646_));
  NA3        o0618(.A(ori_ori_n560_), .B(ori_ori_n268_), .C(ori_ori_n141_), .Y(ori_ori_n647_));
  NA2        o0619(.A(ori_ori_n516_), .B(ori_ori_n157_), .Y(ori_ori_n648_));
  NO3        o0620(.A(ori_ori_n396_), .B(ori_ori_n648_), .C(ori_ori_n83_), .Y(ori_ori_n649_));
  AOI210     o0621(.A0(ori_ori_n647_), .A1(ori_ori_n646_), .B0(ori_ori_n649_), .Y(ori_ori_n650_));
  AN3        o0622(.A(f), .B(d), .C(b), .Y(ori_ori_n651_));
  OAI210     o0623(.A0(ori_ori_n651_), .A1(ori_ori_n126_), .B0(n), .Y(ori_ori_n652_));
  NA3        o0624(.A(ori_ori_n516_), .B(ori_ori_n157_), .C(ori_ori_n213_), .Y(ori_ori_n653_));
  AOI210     o0625(.A0(ori_ori_n652_), .A1(ori_ori_n232_), .B0(ori_ori_n653_), .Y(ori_ori_n654_));
  NAi31      o0626(.An(m), .B(n), .C(k), .Y(ori_ori_n655_));
  OR2        o0627(.A(ori_ori_n131_), .B(ori_ori_n60_), .Y(ori_ori_n656_));
  OAI210     o0628(.A0(ori_ori_n656_), .A1(ori_ori_n655_), .B0(ori_ori_n250_), .Y(ori_ori_n657_));
  OAI210     o0629(.A0(ori_ori_n657_), .A1(ori_ori_n654_), .B0(j), .Y(ori_ori_n658_));
  NA3        o0630(.A(ori_ori_n658_), .B(ori_ori_n650_), .C(ori_ori_n645_), .Y(ori_ori_n659_));
  NO4        o0631(.A(ori_ori_n659_), .B(ori_ori_n640_), .C(ori_ori_n628_), .D(ori_ori_n622_), .Y(ori_ori_n660_));
  NA2        o0632(.A(ori_ori_n383_), .B(ori_ori_n160_), .Y(ori_ori_n661_));
  NAi31      o0633(.An(o), .B(h), .C(f), .Y(ori_ori_n662_));
  OA210      o0634(.A0(ori_ori_n542_), .A1(n), .B0(ori_ori_n594_), .Y(ori_ori_n663_));
  NO2        o0635(.A(ori_ori_n663_), .B(ori_ori_n87_), .Y(ori_ori_n664_));
  INV        o0636(.A(ori_ori_n664_), .Y(ori_ori_n665_));
  AOI210     o0637(.A0(ori_ori_n665_), .A1(ori_ori_n661_), .B0(ori_ori_n536_), .Y(ori_ori_n666_));
  NO3        o0638(.A(o), .B(ori_ori_n212_), .C(ori_ori_n56_), .Y(ori_ori_n667_));
  NAi21      o0639(.An(h), .B(j), .Y(ori_ori_n668_));
  NO2        o0640(.A(ori_ori_n523_), .B(ori_ori_n83_), .Y(ori_ori_n669_));
  OAI210     o0641(.A0(ori_ori_n669_), .A1(ori_ori_n395_), .B0(ori_ori_n667_), .Y(ori_ori_n670_));
  OR2        o0642(.A(ori_ori_n68_), .B(ori_ori_n69_), .Y(ori_ori_n671_));
  NA2        o0643(.A(ori_ori_n604_), .B(ori_ori_n343_), .Y(ori_ori_n672_));
  OA220      o0644(.A0(ori_ori_n635_), .A1(ori_ori_n672_), .B0(ori_ori_n632_), .B1(ori_ori_n671_), .Y(ori_ori_n673_));
  AN2        o0645(.A(h), .B(f), .Y(ori_ori_n674_));
  NA2        o0646(.A(ori_ori_n674_), .B(ori_ori_n37_), .Y(ori_ori_n675_));
  NA2        o0647(.A(ori_ori_n96_), .B(ori_ori_n46_), .Y(ori_ori_n676_));
  OAI220     o0648(.A0(ori_ori_n676_), .A1(ori_ori_n332_), .B0(ori_ori_n675_), .B1(ori_ori_n472_), .Y(ori_ori_n677_));
  AOI210     o0649(.A0(ori_ori_n574_), .A1(ori_ori_n431_), .B0(ori_ori_n49_), .Y(ori_ori_n678_));
  OAI220     o0650(.A0(ori_ori_n597_), .A1(ori_ori_n590_), .B0(ori_ori_n325_), .B1(ori_ori_n534_), .Y(ori_ori_n679_));
  AOI210     o0651(.A0(ori_ori_n679_), .A1(ori_ori_n678_), .B0(ori_ori_n677_), .Y(ori_ori_n680_));
  NA3        o0652(.A(ori_ori_n680_), .B(ori_ori_n673_), .C(ori_ori_n670_), .Y(ori_ori_n681_));
  NO2        o0653(.A(ori_ori_n252_), .B(f), .Y(ori_ori_n682_));
  NO2        o0654(.A(ori_ori_n625_), .B(ori_ori_n60_), .Y(ori_ori_n683_));
  NO3        o0655(.A(ori_ori_n683_), .B(ori_ori_n682_), .C(ori_ori_n34_), .Y(ori_ori_n684_));
  NA2        o0656(.A(ori_ori_n328_), .B(ori_ori_n136_), .Y(ori_ori_n685_));
  NA2        o0657(.A(ori_ori_n128_), .B(ori_ori_n49_), .Y(ori_ori_n686_));
  AOI220     o0658(.A0(ori_ori_n686_), .A1(ori_ori_n539_), .B0(ori_ori_n364_), .B1(ori_ori_n110_), .Y(ori_ori_n687_));
  OA220      o0659(.A0(ori_ori_n687_), .A1(ori_ori_n557_), .B0(ori_ori_n362_), .B1(ori_ori_n108_), .Y(ori_ori_n688_));
  OAI210     o0660(.A0(ori_ori_n685_), .A1(ori_ori_n684_), .B0(ori_ori_n688_), .Y(ori_ori_n689_));
  NO3        o0661(.A(ori_ori_n406_), .B(ori_ori_n190_), .C(ori_ori_n189_), .Y(ori_ori_n690_));
  NA2        o0662(.A(ori_ori_n690_), .B(ori_ori_n230_), .Y(ori_ori_n691_));
  NA3        o0663(.A(ori_ori_n691_), .B(ori_ori_n254_), .C(j), .Y(ori_ori_n692_));
  NO3        o0664(.A(ori_ori_n467_), .B(ori_ori_n171_), .C(i), .Y(ori_ori_n693_));
  NA2        o0665(.A(ori_ori_n471_), .B(ori_ori_n80_), .Y(ori_ori_n694_));
  NO4        o0666(.A(ori_ori_n536_), .B(ori_ori_n694_), .C(ori_ori_n127_), .D(ori_ori_n212_), .Y(ori_ori_n695_));
  INV        o0667(.A(ori_ori_n695_), .Y(ori_ori_n696_));
  NA3        o0668(.A(ori_ori_n696_), .B(ori_ori_n692_), .C(ori_ori_n404_), .Y(ori_ori_n697_));
  NO4        o0669(.A(ori_ori_n697_), .B(ori_ori_n689_), .C(ori_ori_n681_), .D(ori_ori_n666_), .Y(ori_ori_n698_));
  NA4        o0670(.A(ori_ori_n698_), .B(ori_ori_n660_), .C(ori_ori_n615_), .D(ori_ori_n588_), .Y(ori08));
  NO2        o0671(.A(k), .B(h), .Y(ori_ori_n700_));
  AO210      o0672(.A0(ori_ori_n252_), .A1(ori_ori_n455_), .B0(ori_ori_n700_), .Y(ori_ori_n701_));
  NO2        o0673(.A(ori_ori_n701_), .B(ori_ori_n296_), .Y(ori_ori_n702_));
  NA2        o0674(.A(ori_ori_n624_), .B(ori_ori_n80_), .Y(ori_ori_n703_));
  NA2        o0675(.A(ori_ori_n703_), .B(ori_ori_n467_), .Y(ori_ori_n704_));
  AOI210     o0676(.A0(ori_ori_n704_), .A1(ori_ori_n702_), .B0(ori_ori_n500_), .Y(ori_ori_n705_));
  NA2        o0677(.A(ori_ori_n80_), .B(ori_ori_n107_), .Y(ori_ori_n706_));
  NO2        o0678(.A(ori_ori_n706_), .B(ori_ori_n57_), .Y(ori_ori_n707_));
  NO4        o0679(.A(ori_ori_n380_), .B(ori_ori_n109_), .C(j), .D(ori_ori_n213_), .Y(ori_ori_n708_));
  NA2        o0680(.A(ori_ori_n584_), .B(ori_ori_n232_), .Y(ori_ori_n709_));
  AOI220     o0681(.A0(ori_ori_n709_), .A1(ori_ori_n349_), .B0(ori_ori_n708_), .B1(ori_ori_n707_), .Y(ori_ori_n710_));
  AOI210     o0682(.A0(ori_ori_n584_), .A1(ori_ori_n153_), .B0(ori_ori_n80_), .Y(ori_ori_n711_));
  NA4        o0683(.A(ori_ori_n215_), .B(ori_ori_n136_), .C(ori_ori_n45_), .D(h), .Y(ori_ori_n712_));
  AN2        o0684(.A(l), .B(k), .Y(ori_ori_n713_));
  NA4        o0685(.A(ori_ori_n713_), .B(ori_ori_n106_), .C(ori_ori_n69_), .D(ori_ori_n213_), .Y(ori_ori_n714_));
  OAI210     o0686(.A0(ori_ori_n712_), .A1(o), .B0(ori_ori_n714_), .Y(ori_ori_n715_));
  NA2        o0687(.A(ori_ori_n715_), .B(ori_ori_n711_), .Y(ori_ori_n716_));
  NA4        o0688(.A(ori_ori_n716_), .B(ori_ori_n710_), .C(ori_ori_n705_), .D(ori_ori_n351_), .Y(ori_ori_n717_));
  AN2        o0689(.A(ori_ori_n543_), .B(ori_ori_n92_), .Y(ori_ori_n718_));
  NO4        o0690(.A(ori_ori_n171_), .B(ori_ori_n394_), .C(ori_ori_n109_), .D(o), .Y(ori_ori_n719_));
  NA2        o0691(.A(ori_ori_n719_), .B(ori_ori_n709_), .Y(ori_ori_n720_));
  NO2        o0692(.A(ori_ori_n38_), .B(ori_ori_n212_), .Y(ori_ori_n721_));
  AOI220     o0693(.A0(ori_ori_n626_), .A1(ori_ori_n348_), .B0(ori_ori_n721_), .B1(ori_ori_n571_), .Y(ori_ori_n722_));
  NAi31      o0694(.An(ori_ori_n718_), .B(ori_ori_n722_), .C(ori_ori_n720_), .Y(ori_ori_n723_));
  OAI210     o0695(.A0(ori_ori_n560_), .A1(ori_ori_n47_), .B0(ori_ori_n656_), .Y(ori_ori_n724_));
  NO2        o0696(.A(ori_ori_n494_), .B(ori_ori_n128_), .Y(ori_ori_n725_));
  NA2        o0697(.A(ori_ori_n725_), .B(ori_ori_n724_), .Y(ori_ori_n726_));
  NO3        o0698(.A(ori_ori_n315_), .B(ori_ori_n127_), .C(ori_ori_n41_), .Y(ori_ori_n727_));
  NAi21      o0699(.An(ori_ori_n727_), .B(ori_ori_n714_), .Y(ori_ori_n728_));
  NA2        o0700(.A(ori_ori_n701_), .B(ori_ori_n132_), .Y(ori_ori_n729_));
  AOI220     o0701(.A0(ori_ori_n729_), .A1(ori_ori_n405_), .B0(ori_ori_n728_), .B1(ori_ori_n72_), .Y(ori_ori_n730_));
  NA2        o0702(.A(ori_ori_n726_), .B(ori_ori_n730_), .Y(ori_ori_n731_));
  NA2        o0703(.A(ori_ori_n364_), .B(ori_ori_n43_), .Y(ori_ori_n732_));
  NA3        o0704(.A(ori_ori_n691_), .B(ori_ori_n334_), .C(ori_ori_n386_), .Y(ori_ori_n733_));
  NA3        o0705(.A(m), .B(l), .C(k), .Y(ori_ori_n734_));
  NA4        o0706(.A(ori_ori_n110_), .B(l), .C(k), .D(ori_ori_n83_), .Y(ori_ori_n735_));
  NA2        o0707(.A(ori_ori_n733_), .B(ori_ori_n732_), .Y(ori_ori_n736_));
  NO4        o0708(.A(ori_ori_n736_), .B(ori_ori_n731_), .C(ori_ori_n723_), .D(ori_ori_n717_), .Y(ori_ori_n737_));
  NA2        o0709(.A(ori_ori_n626_), .B(ori_ori_n395_), .Y(ori_ori_n738_));
  NO3        o0710(.A(ori_ori_n399_), .B(ori_ori_n534_), .C(h), .Y(ori_ori_n739_));
  AOI210     o0711(.A0(ori_ori_n739_), .A1(ori_ori_n110_), .B0(ori_ori_n510_), .Y(ori_ori_n740_));
  NA3        o0712(.A(ori_ori_n740_), .B(ori_ori_n738_), .C(ori_ori_n251_), .Y(ori_ori_n741_));
  NA2        o0713(.A(ori_ori_n713_), .B(ori_ori_n69_), .Y(ori_ori_n742_));
  NO4        o0714(.A(ori_ori_n690_), .B(ori_ori_n171_), .C(n), .D(i), .Y(ori_ori_n743_));
  NOi21      o0715(.An(h), .B(j), .Y(ori_ori_n744_));
  NA2        o0716(.A(ori_ori_n744_), .B(f), .Y(ori_ori_n745_));
  NO2        o0717(.A(ori_ori_n743_), .B(ori_ori_n693_), .Y(ori_ori_n746_));
  NO2        o0718(.A(ori_ori_n746_), .B(ori_ori_n742_), .Y(ori_ori_n747_));
  AOI210     o0719(.A0(ori_ori_n741_), .A1(l), .B0(ori_ori_n747_), .Y(ori_ori_n748_));
  NO2        o0720(.A(j), .B(i), .Y(ori_ori_n749_));
  NA3        o0721(.A(ori_ori_n749_), .B(ori_ori_n76_), .C(l), .Y(ori_ori_n750_));
  NA2        o0722(.A(ori_ori_n749_), .B(ori_ori_n33_), .Y(ori_ori_n751_));
  OR2        o0723(.A(ori_ori_n750_), .B(ori_ori_n596_), .Y(ori_ori_n752_));
  NO3        o0724(.A(ori_ori_n148_), .B(ori_ori_n49_), .C(ori_ori_n107_), .Y(ori_ori_n753_));
  NO3        o0725(.A(ori_ori_n549_), .B(ori_ori_n146_), .C(ori_ori_n69_), .Y(ori_ori_n754_));
  NO3        o0726(.A(ori_ori_n494_), .B(ori_ori_n442_), .C(j), .Y(ori_ori_n755_));
  OAI210     o0727(.A0(ori_ori_n754_), .A1(ori_ori_n753_), .B0(ori_ori_n755_), .Y(ori_ori_n756_));
  INV        o0728(.A(ori_ori_n756_), .Y(ori_ori_n757_));
  NA2        o0729(.A(k), .B(j), .Y(ori_ori_n758_));
  NO3        o0730(.A(ori_ori_n296_), .B(ori_ori_n758_), .C(ori_ori_n40_), .Y(ori_ori_n759_));
  AOI210     o0731(.A0(ori_ori_n539_), .A1(n), .B0(ori_ori_n559_), .Y(ori_ori_n760_));
  NA2        o0732(.A(ori_ori_n760_), .B(ori_ori_n562_), .Y(ori_ori_n761_));
  AN3        o0733(.A(ori_ori_n761_), .B(ori_ori_n759_), .C(ori_ori_n95_), .Y(ori_ori_n762_));
  NO3        o0734(.A(ori_ori_n171_), .B(ori_ori_n394_), .C(ori_ori_n109_), .Y(ori_ori_n763_));
  AOI220     o0735(.A0(ori_ori_n763_), .A1(ori_ori_n246_), .B0(ori_ori_n618_), .B1(ori_ori_n307_), .Y(ori_ori_n764_));
  NAi31      o0736(.An(ori_ori_n611_), .B(ori_ori_n89_), .C(ori_ori_n80_), .Y(ori_ori_n765_));
  NA2        o0737(.A(ori_ori_n765_), .B(ori_ori_n764_), .Y(ori_ori_n766_));
  NO2        o0738(.A(ori_ori_n296_), .B(ori_ori_n132_), .Y(ori_ori_n767_));
  AOI220     o0739(.A0(ori_ori_n767_), .A1(ori_ori_n626_), .B0(ori_ori_n727_), .B1(ori_ori_n711_), .Y(ori_ori_n768_));
  NO2        o0740(.A(ori_ori_n734_), .B(ori_ori_n87_), .Y(ori_ori_n769_));
  NA2        o0741(.A(ori_ori_n769_), .B(ori_ori_n595_), .Y(ori_ori_n770_));
  NO2        o0742(.A(ori_ori_n597_), .B(ori_ori_n113_), .Y(ori_ori_n771_));
  OAI210     o0743(.A0(ori_ori_n771_), .A1(ori_ori_n755_), .B0(ori_ori_n678_), .Y(ori_ori_n772_));
  NA3        o0744(.A(ori_ori_n772_), .B(ori_ori_n770_), .C(ori_ori_n768_), .Y(ori_ori_n773_));
  OR4        o0745(.A(ori_ori_n773_), .B(ori_ori_n766_), .C(ori_ori_n762_), .D(ori_ori_n757_), .Y(ori_ori_n774_));
  NA3        o0746(.A(ori_ori_n760_), .B(ori_ori_n562_), .C(ori_ori_n561_), .Y(ori_ori_n775_));
  NA4        o0747(.A(ori_ori_n775_), .B(ori_ori_n215_), .C(ori_ori_n455_), .D(ori_ori_n34_), .Y(ori_ori_n776_));
  NO4        o0748(.A(ori_ori_n494_), .B(ori_ori_n438_), .C(j), .D(f), .Y(ori_ori_n777_));
  OAI220     o0749(.A0(ori_ori_n712_), .A1(ori_ori_n703_), .B0(ori_ori_n332_), .B1(ori_ori_n38_), .Y(ori_ori_n778_));
  AOI210     o0750(.A0(ori_ori_n777_), .A1(ori_ori_n258_), .B0(ori_ori_n778_), .Y(ori_ori_n779_));
  NA3        o0751(.A(ori_ori_n552_), .B(ori_ori_n289_), .C(h), .Y(ori_ori_n780_));
  NOi21      o0752(.An(ori_ori_n678_), .B(ori_ori_n780_), .Y(ori_ori_n781_));
  NO2        o0753(.A(ori_ori_n88_), .B(ori_ori_n47_), .Y(ori_ori_n782_));
  OAI220     o0754(.A0(ori_ori_n780_), .A1(ori_ori_n608_), .B0(ori_ori_n750_), .B1(ori_ori_n671_), .Y(ori_ori_n783_));
  AOI210     o0755(.A0(ori_ori_n782_), .A1(ori_ori_n644_), .B0(ori_ori_n783_), .Y(ori_ori_n784_));
  NAi41      o0756(.An(ori_ori_n781_), .B(ori_ori_n784_), .C(ori_ori_n779_), .D(ori_ori_n776_), .Y(ori_ori_n785_));
  AOI220     o0757(.A0(ori_ori_n769_), .A1(ori_ori_n237_), .B0(ori_ori_n755_), .B1(ori_ori_n636_), .Y(ori_ori_n786_));
  NO2        o0758(.A(ori_ori_n663_), .B(ori_ori_n69_), .Y(ori_ori_n787_));
  AOI210     o0759(.A0(ori_ori_n777_), .A1(ori_ori_n787_), .B0(ori_ori_n336_), .Y(ori_ori_n788_));
  OAI210     o0760(.A0(ori_ori_n734_), .A1(ori_ori_n662_), .B0(ori_ori_n528_), .Y(ori_ori_n789_));
  NA3        o0761(.A(ori_ori_n249_), .B(ori_ori_n59_), .C(b), .Y(ori_ori_n790_));
  AOI220     o0762(.A0(ori_ori_n607_), .A1(ori_ori_n29_), .B0(ori_ori_n471_), .B1(ori_ori_n80_), .Y(ori_ori_n791_));
  NA2        o0763(.A(ori_ori_n791_), .B(ori_ori_n790_), .Y(ori_ori_n792_));
  NA2        o0764(.A(ori_ori_n792_), .B(ori_ori_n789_), .Y(ori_ori_n793_));
  NA3        o0765(.A(ori_ori_n793_), .B(ori_ori_n788_), .C(ori_ori_n786_), .Y(ori_ori_n794_));
  NOi41      o0766(.An(ori_ori_n752_), .B(ori_ori_n794_), .C(ori_ori_n785_), .D(ori_ori_n774_), .Y(ori_ori_n795_));
  NO3        o0767(.A(ori_ori_n342_), .B(ori_ori_n298_), .C(ori_ori_n109_), .Y(ori_ori_n796_));
  NA2        o0768(.A(ori_ori_n796_), .B(ori_ori_n761_), .Y(ori_ori_n797_));
  NO3        o0769(.A(ori_ori_n534_), .B(ori_ori_n90_), .C(h), .Y(ori_ori_n798_));
  NA2        o0770(.A(ori_ori_n798_), .B(ori_ori_n707_), .Y(ori_ori_n799_));
  NA3        o0771(.A(ori_ori_n799_), .B(ori_ori_n797_), .C(ori_ori_n407_), .Y(ori_ori_n800_));
  OR2        o0772(.A(ori_ori_n662_), .B(ori_ori_n88_), .Y(ori_ori_n801_));
  NOi31      o0773(.An(b), .B(d), .C(a), .Y(ori_ori_n802_));
  NO2        o0774(.A(ori_ori_n802_), .B(ori_ori_n605_), .Y(ori_ori_n803_));
  NO2        o0775(.A(ori_ori_n803_), .B(n), .Y(ori_ori_n804_));
  NOi21      o0776(.An(ori_ori_n791_), .B(ori_ori_n804_), .Y(ori_ori_n805_));
  OAI220     o0777(.A0(ori_ori_n805_), .A1(ori_ori_n801_), .B0(ori_ori_n780_), .B1(ori_ori_n606_), .Y(ori_ori_n806_));
  NO2        o0778(.A(ori_ori_n560_), .B(ori_ori_n80_), .Y(ori_ori_n807_));
  NA2        o0779(.A(ori_ori_n796_), .B(ori_ori_n807_), .Y(ori_ori_n808_));
  OAI210     o0780(.A0(ori_ori_n712_), .A1(ori_ori_n396_), .B0(ori_ori_n808_), .Y(ori_ori_n809_));
  NO2        o0781(.A(ori_ori_n690_), .B(n), .Y(ori_ori_n810_));
  AOI220     o0782(.A0(ori_ori_n767_), .A1(ori_ori_n667_), .B0(ori_ori_n810_), .B1(ori_ori_n702_), .Y(ori_ori_n811_));
  NO2        o0783(.A(ori_ori_n322_), .B(ori_ori_n236_), .Y(ori_ori_n812_));
  OAI210     o0784(.A0(ori_ori_n92_), .A1(ori_ori_n89_), .B0(ori_ori_n812_), .Y(ori_ori_n813_));
  INV        o0785(.A(ori_ori_n813_), .Y(ori_ori_n814_));
  NA2        o0786(.A(ori_ori_n719_), .B(ori_ori_n350_), .Y(ori_ori_n815_));
  OAI210     o0787(.A0(ori_ori_n600_), .A1(ori_ori_n599_), .B0(ori_ori_n365_), .Y(ori_ori_n816_));
  AN2        o0788(.A(ori_ori_n816_), .B(ori_ori_n815_), .Y(ori_ori_n817_));
  NAi31      o0789(.An(ori_ori_n814_), .B(ori_ori_n817_), .C(ori_ori_n811_), .Y(ori_ori_n818_));
  NO4        o0790(.A(ori_ori_n818_), .B(ori_ori_n809_), .C(ori_ori_n806_), .D(ori_ori_n800_), .Y(ori_ori_n819_));
  NA4        o0791(.A(ori_ori_n819_), .B(ori_ori_n795_), .C(ori_ori_n748_), .D(ori_ori_n737_), .Y(ori09));
  INV        o0792(.A(ori_ori_n118_), .Y(ori_ori_n821_));
  NA2        o0793(.A(f), .B(e), .Y(ori_ori_n822_));
  NO2        o0794(.A(ori_ori_n225_), .B(ori_ori_n109_), .Y(ori_ori_n823_));
  NA2        o0795(.A(ori_ori_n823_), .B(o), .Y(ori_ori_n824_));
  NA4        o0796(.A(ori_ori_n309_), .B(ori_ori_n480_), .C(ori_ori_n261_), .D(ori_ori_n115_), .Y(ori_ori_n825_));
  AOI210     o0797(.A0(ori_ori_n825_), .A1(o), .B0(ori_ori_n477_), .Y(ori_ori_n826_));
  AOI210     o0798(.A0(ori_ori_n826_), .A1(ori_ori_n824_), .B0(ori_ori_n822_), .Y(ori_ori_n827_));
  NA2        o0799(.A(ori_ori_n448_), .B(e), .Y(ori_ori_n828_));
  NO2        o0800(.A(ori_ori_n828_), .B(ori_ori_n520_), .Y(ori_ori_n829_));
  AOI210     o0801(.A0(ori_ori_n827_), .A1(ori_ori_n821_), .B0(ori_ori_n829_), .Y(ori_ori_n830_));
  NO2        o0802(.A(ori_ori_n202_), .B(ori_ori_n212_), .Y(ori_ori_n831_));
  NA3        o0803(.A(m), .B(l), .C(i), .Y(ori_ori_n832_));
  OAI220     o0804(.A0(ori_ori_n597_), .A1(ori_ori_n832_), .B0(ori_ori_n355_), .B1(ori_ori_n535_), .Y(ori_ori_n833_));
  NA4        o0805(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(o), .D(f), .Y(ori_ori_n834_));
  NAi31      o0806(.An(ori_ori_n833_), .B(ori_ori_n834_), .C(ori_ori_n443_), .Y(ori_ori_n835_));
  OA210      o0807(.A0(ori_ori_n835_), .A1(ori_ori_n831_), .B0(ori_ori_n571_), .Y(ori_ori_n836_));
  NA3        o0808(.A(ori_ori_n801_), .B(ori_ori_n573_), .C(ori_ori_n528_), .Y(ori_ori_n837_));
  OA210      o0809(.A0(ori_ori_n837_), .A1(ori_ori_n836_), .B0(ori_ori_n804_), .Y(ori_ori_n838_));
  INV        o0810(.A(ori_ori_n339_), .Y(ori_ori_n839_));
  NO2        o0811(.A(ori_ori_n123_), .B(ori_ori_n121_), .Y(ori_ori_n840_));
  NOi31      o0812(.An(k), .B(m), .C(l), .Y(ori_ori_n841_));
  NO2        o0813(.A(ori_ori_n341_), .B(ori_ori_n841_), .Y(ori_ori_n842_));
  AOI210     o0814(.A0(ori_ori_n842_), .A1(ori_ori_n840_), .B0(ori_ori_n603_), .Y(ori_ori_n843_));
  NA2        o0815(.A(ori_ori_n790_), .B(ori_ori_n332_), .Y(ori_ori_n844_));
  NA2        o0816(.A(ori_ori_n343_), .B(ori_ori_n345_), .Y(ori_ori_n845_));
  OAI210     o0817(.A0(ori_ori_n202_), .A1(ori_ori_n212_), .B0(ori_ori_n845_), .Y(ori_ori_n846_));
  AOI220     o0818(.A0(ori_ori_n846_), .A1(ori_ori_n844_), .B0(ori_ori_n843_), .B1(ori_ori_n839_), .Y(ori_ori_n847_));
  NA2        o0819(.A(ori_ori_n166_), .B(ori_ori_n111_), .Y(ori_ori_n848_));
  NA3        o0820(.A(ori_ori_n848_), .B(ori_ori_n701_), .C(ori_ori_n132_), .Y(ori_ori_n849_));
  NA3        o0821(.A(ori_ori_n849_), .B(ori_ori_n187_), .C(ori_ori_n31_), .Y(ori_ori_n850_));
  NA4        o0822(.A(ori_ori_n850_), .B(ori_ori_n847_), .C(ori_ori_n627_), .D(ori_ori_n78_), .Y(ori_ori_n851_));
  NO2        o0823(.A(ori_ori_n593_), .B(ori_ori_n506_), .Y(ori_ori_n852_));
  NA2        o0824(.A(ori_ori_n852_), .B(ori_ori_n187_), .Y(ori_ori_n853_));
  NOi21      o0825(.An(f), .B(d), .Y(ori_ori_n854_));
  NA2        o0826(.A(ori_ori_n854_), .B(m), .Y(ori_ori_n855_));
  NO2        o0827(.A(ori_ori_n855_), .B(ori_ori_n52_), .Y(ori_ori_n856_));
  NOi32      o0828(.An(o), .Bn(f), .C(d), .Y(ori_ori_n857_));
  NA4        o0829(.A(ori_ori_n857_), .B(ori_ori_n607_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n858_));
  NOi21      o0830(.An(ori_ori_n310_), .B(ori_ori_n858_), .Y(ori_ori_n859_));
  AOI210     o0831(.A0(ori_ori_n856_), .A1(ori_ori_n550_), .B0(ori_ori_n859_), .Y(ori_ori_n860_));
  NA3        o0832(.A(ori_ori_n309_), .B(ori_ori_n261_), .C(ori_ori_n115_), .Y(ori_ori_n861_));
  AN2        o0833(.A(f), .B(d), .Y(ori_ori_n862_));
  NA3        o0834(.A(ori_ori_n485_), .B(ori_ori_n862_), .C(ori_ori_n80_), .Y(ori_ori_n863_));
  NO3        o0835(.A(ori_ori_n863_), .B(ori_ori_n69_), .C(ori_ori_n213_), .Y(ori_ori_n864_));
  NA2        o0836(.A(ori_ori_n861_), .B(ori_ori_n864_), .Y(ori_ori_n865_));
  NAi41      o0837(.An(ori_ori_n499_), .B(ori_ori_n865_), .C(ori_ori_n860_), .D(ori_ori_n853_), .Y(ori_ori_n866_));
  NO4        o0838(.A(ori_ori_n625_), .B(ori_ori_n128_), .C(ori_ori_n327_), .D(ori_ori_n149_), .Y(ori_ori_n867_));
  NO2        o0839(.A(ori_ori_n655_), .B(ori_ori_n327_), .Y(ori_ori_n868_));
  AN2        o0840(.A(ori_ori_n868_), .B(ori_ori_n682_), .Y(ori_ori_n869_));
  NO2        o0841(.A(ori_ori_n869_), .B(ori_ori_n867_), .Y(ori_ori_n870_));
  NA2        o0842(.A(ori_ori_n605_), .B(ori_ori_n80_), .Y(ori_ori_n871_));
  OAI220     o0843(.A0(ori_ori_n845_), .A1(ori_ori_n871_), .B0(ori_ori_n790_), .B1(ori_ori_n443_), .Y(ori_ori_n872_));
  NA3        o0844(.A(ori_ori_n157_), .B(ori_ori_n106_), .C(ori_ori_n105_), .Y(ori_ori_n873_));
  OAI220     o0845(.A0(ori_ori_n863_), .A1(ori_ori_n433_), .B0(ori_ori_n339_), .B1(ori_ori_n873_), .Y(ori_ori_n874_));
  NOi41      o0846(.An(ori_ori_n223_), .B(ori_ori_n874_), .C(ori_ori_n872_), .D(ori_ori_n305_), .Y(ori_ori_n875_));
  NA2        o0847(.A(c), .B(ori_ori_n112_), .Y(ori_ori_n876_));
  NO2        o0848(.A(ori_ori_n876_), .B(ori_ori_n411_), .Y(ori_ori_n877_));
  NA3        o0849(.A(ori_ori_n877_), .B(ori_ori_n518_), .C(f), .Y(ori_ori_n878_));
  OR2        o0850(.A(ori_ori_n662_), .B(ori_ori_n546_), .Y(ori_ori_n879_));
  INV        o0851(.A(ori_ori_n879_), .Y(ori_ori_n880_));
  NA2        o0852(.A(ori_ori_n803_), .B(ori_ori_n108_), .Y(ori_ori_n881_));
  NA2        o0853(.A(ori_ori_n881_), .B(ori_ori_n880_), .Y(ori_ori_n882_));
  NA4        o0854(.A(ori_ori_n882_), .B(ori_ori_n878_), .C(ori_ori_n875_), .D(ori_ori_n870_), .Y(ori_ori_n883_));
  NO4        o0855(.A(ori_ori_n883_), .B(ori_ori_n866_), .C(ori_ori_n851_), .D(ori_ori_n838_), .Y(ori_ori_n884_));
  OR2        o0856(.A(ori_ori_n863_), .B(ori_ori_n69_), .Y(ori_ori_n885_));
  NA2        o0857(.A(ori_ori_n823_), .B(o), .Y(ori_ori_n886_));
  AOI210     o0858(.A0(ori_ori_n886_), .A1(ori_ori_n290_), .B0(ori_ori_n885_), .Y(ori_ori_n887_));
  AOI210     o0859(.A0(ori_ori_n790_), .A1(ori_ori_n332_), .B0(ori_ori_n834_), .Y(ori_ori_n888_));
  NO2        o0860(.A(ori_ori_n132_), .B(ori_ori_n128_), .Y(ori_ori_n889_));
  NO2        o0861(.A(ori_ori_n230_), .B(ori_ori_n224_), .Y(ori_ori_n890_));
  AOI220     o0862(.A0(ori_ori_n890_), .A1(ori_ori_n227_), .B0(ori_ori_n303_), .B1(ori_ori_n889_), .Y(ori_ori_n891_));
  NO2        o0863(.A(ori_ori_n433_), .B(ori_ori_n822_), .Y(ori_ori_n892_));
  NA2        o0864(.A(ori_ori_n892_), .B(ori_ori_n567_), .Y(ori_ori_n893_));
  NA2        o0865(.A(ori_ori_n893_), .B(ori_ori_n891_), .Y(ori_ori_n894_));
  NA2        o0866(.A(e), .B(d), .Y(ori_ori_n895_));
  OAI220     o0867(.A0(ori_ori_n895_), .A1(c), .B0(ori_ori_n322_), .B1(d), .Y(ori_ori_n896_));
  NA3        o0868(.A(ori_ori_n896_), .B(ori_ori_n460_), .C(ori_ori_n516_), .Y(ori_ori_n897_));
  AOI210     o0869(.A0(ori_ori_n523_), .A1(ori_ori_n178_), .B0(ori_ori_n230_), .Y(ori_ori_n898_));
  AOI210     o0870(.A0(ori_ori_n626_), .A1(ori_ori_n348_), .B0(ori_ori_n898_), .Y(ori_ori_n899_));
  NA2        o0871(.A(ori_ori_n282_), .B(ori_ori_n162_), .Y(ori_ori_n900_));
  NA2        o0872(.A(ori_ori_n864_), .B(ori_ori_n900_), .Y(ori_ori_n901_));
  NA3        o0873(.A(ori_ori_n165_), .B(ori_ori_n81_), .C(ori_ori_n34_), .Y(ori_ori_n902_));
  NA4        o0874(.A(ori_ori_n902_), .B(ori_ori_n901_), .C(ori_ori_n899_), .D(ori_ori_n897_), .Y(ori_ori_n903_));
  NO4        o0875(.A(ori_ori_n903_), .B(ori_ori_n894_), .C(ori_ori_n888_), .D(ori_ori_n887_), .Y(ori_ori_n904_));
  OR2        o0876(.A(ori_ori_n703_), .B(ori_ori_n216_), .Y(ori_ori_n905_));
  OAI220     o0877(.A0(ori_ori_n625_), .A1(ori_ori_n60_), .B0(ori_ori_n298_), .B1(j), .Y(ori_ori_n906_));
  AOI220     o0878(.A0(ori_ori_n906_), .A1(ori_ori_n868_), .B0(ori_ori_n616_), .B1(ori_ori_n624_), .Y(ori_ori_n907_));
  OAI210     o0879(.A0(ori_ori_n828_), .A1(ori_ori_n168_), .B0(ori_ori_n907_), .Y(ori_ori_n908_));
  OAI210     o0880(.A0(ori_ori_n823_), .A1(ori_ori_n900_), .B0(ori_ori_n857_), .Y(ori_ori_n909_));
  NO2        o0881(.A(ori_ori_n909_), .B(ori_ori_n608_), .Y(ori_ori_n910_));
  AOI210     o0882(.A0(ori_ori_n114_), .A1(ori_ori_n113_), .B0(ori_ori_n260_), .Y(ori_ori_n911_));
  NO2        o0883(.A(ori_ori_n911_), .B(ori_ori_n858_), .Y(ori_ori_n912_));
  AO210      o0884(.A0(ori_ori_n844_), .A1(ori_ori_n833_), .B0(ori_ori_n912_), .Y(ori_ori_n913_));
  NOi31      o0885(.An(ori_ori_n550_), .B(ori_ori_n855_), .C(ori_ori_n290_), .Y(ori_ori_n914_));
  NO4        o0886(.A(ori_ori_n914_), .B(ori_ori_n913_), .C(ori_ori_n910_), .D(ori_ori_n908_), .Y(ori_ori_n915_));
  AO220      o0887(.A0(ori_ori_n460_), .A1(ori_ori_n744_), .B0(ori_ori_n173_), .B1(f), .Y(ori_ori_n916_));
  OAI210     o0888(.A0(ori_ori_n916_), .A1(ori_ori_n463_), .B0(ori_ori_n896_), .Y(ori_ori_n917_));
  NO2        o0889(.A(ori_ori_n442_), .B(ori_ori_n66_), .Y(ori_ori_n918_));
  OAI210     o0890(.A0(ori_ori_n837_), .A1(ori_ori_n918_), .B0(ori_ori_n707_), .Y(ori_ori_n919_));
  AN4        o0891(.A(ori_ori_n919_), .B(ori_ori_n917_), .C(ori_ori_n915_), .D(ori_ori_n905_), .Y(ori_ori_n920_));
  NA4        o0892(.A(ori_ori_n920_), .B(ori_ori_n904_), .C(ori_ori_n884_), .D(ori_ori_n830_), .Y(ori12));
  NO2        o0893(.A(ori_ori_n458_), .B(c), .Y(ori_ori_n922_));
  NO4        o0894(.A(ori_ori_n447_), .B(ori_ori_n252_), .C(ori_ori_n589_), .D(ori_ori_n213_), .Y(ori_ori_n923_));
  NA2        o0895(.A(ori_ori_n923_), .B(ori_ori_n922_), .Y(ori_ori_n924_));
  NA2        o0896(.A(ori_ori_n550_), .B(ori_ori_n918_), .Y(ori_ori_n925_));
  NO2        o0897(.A(ori_ori_n458_), .B(ori_ori_n112_), .Y(ori_ori_n926_));
  NO2        o0898(.A(ori_ori_n840_), .B(ori_ori_n355_), .Y(ori_ori_n927_));
  NO2        o0899(.A(ori_ori_n662_), .B(ori_ori_n380_), .Y(ori_ori_n928_));
  AOI220     o0900(.A0(ori_ori_n928_), .A1(ori_ori_n548_), .B0(ori_ori_n927_), .B1(ori_ori_n926_), .Y(ori_ori_n929_));
  NA4        o0901(.A(ori_ori_n929_), .B(ori_ori_n925_), .C(ori_ori_n924_), .D(ori_ori_n446_), .Y(ori_ori_n930_));
  AOI210     o0902(.A0(ori_ori_n233_), .A1(ori_ori_n338_), .B0(ori_ori_n199_), .Y(ori_ori_n931_));
  OR2        o0903(.A(ori_ori_n931_), .B(ori_ori_n923_), .Y(ori_ori_n932_));
  AOI210     o0904(.A0(ori_ori_n335_), .A1(ori_ori_n392_), .B0(ori_ori_n213_), .Y(ori_ori_n933_));
  OAI210     o0905(.A0(ori_ori_n933_), .A1(ori_ori_n932_), .B0(ori_ori_n406_), .Y(ori_ori_n934_));
  NO2        o0906(.A(ori_ori_n641_), .B(ori_ori_n262_), .Y(ori_ori_n935_));
  NO2        o0907(.A(ori_ori_n597_), .B(ori_ori_n832_), .Y(ori_ori_n936_));
  NO2        o0908(.A(ori_ori_n148_), .B(ori_ori_n236_), .Y(ori_ori_n937_));
  NA3        o0909(.A(ori_ori_n937_), .B(ori_ori_n239_), .C(i), .Y(ori_ori_n938_));
  NA2        o0910(.A(ori_ori_n938_), .B(ori_ori_n934_), .Y(ori_ori_n939_));
  OR2        o0911(.A(ori_ori_n323_), .B(ori_ori_n926_), .Y(ori_ori_n940_));
  NA2        o0912(.A(ori_ori_n940_), .B(ori_ori_n356_), .Y(ori_ori_n941_));
  NO3        o0913(.A(ori_ori_n128_), .B(ori_ori_n149_), .C(ori_ori_n213_), .Y(ori_ori_n942_));
  NA2        o0914(.A(ori_ori_n942_), .B(ori_ori_n539_), .Y(ori_ori_n943_));
  NA4        o0915(.A(ori_ori_n448_), .B(ori_ori_n440_), .C(ori_ori_n179_), .D(o), .Y(ori_ori_n944_));
  NA3        o0916(.A(ori_ori_n944_), .B(ori_ori_n943_), .C(ori_ori_n941_), .Y(ori_ori_n945_));
  NO3        o0917(.A(ori_ori_n665_), .B(ori_ori_n88_), .C(ori_ori_n45_), .Y(ori_ori_n946_));
  NO4        o0918(.A(ori_ori_n946_), .B(ori_ori_n945_), .C(ori_ori_n939_), .D(ori_ori_n930_), .Y(ori_ori_n947_));
  NO2        o0919(.A(ori_ori_n372_), .B(ori_ori_n371_), .Y(ori_ori_n948_));
  INV        o0920(.A(ori_ori_n68_), .Y(ori_ori_n949_));
  NA2        o0921(.A(ori_ori_n560_), .B(ori_ori_n141_), .Y(ori_ori_n950_));
  NOi21      o0922(.An(ori_ori_n34_), .B(ori_ori_n655_), .Y(ori_ori_n951_));
  AOI220     o0923(.A0(ori_ori_n951_), .A1(ori_ori_n950_), .B0(ori_ori_n949_), .B1(ori_ori_n948_), .Y(ori_ori_n952_));
  OAI210     o0924(.A0(ori_ori_n250_), .A1(ori_ori_n45_), .B0(ori_ori_n952_), .Y(ori_ori_n953_));
  INV        o0925(.A(ori_ori_n319_), .Y(ori_ori_n954_));
  NO2        o0926(.A(ori_ori_n49_), .B(ori_ori_n45_), .Y(ori_ori_n955_));
  NO2        o0927(.A(ori_ori_n513_), .B(ori_ori_n298_), .Y(ori_ori_n956_));
  INV        o0928(.A(ori_ori_n956_), .Y(ori_ori_n957_));
  NO2        o0929(.A(ori_ori_n957_), .B(ori_ori_n141_), .Y(ori_ori_n958_));
  INV        o0930(.A(ori_ori_n369_), .Y(ori_ori_n959_));
  NO4        o0931(.A(ori_ori_n959_), .B(ori_ori_n958_), .C(ori_ori_n954_), .D(ori_ori_n953_), .Y(ori_ori_n960_));
  NA2        o0932(.A(ori_ori_n348_), .B(o), .Y(ori_ori_n961_));
  NA2        o0933(.A(ori_ori_n160_), .B(i), .Y(ori_ori_n962_));
  NA2        o0934(.A(ori_ori_n46_), .B(i), .Y(ori_ori_n963_));
  OAI220     o0935(.A0(ori_ori_n963_), .A1(ori_ori_n198_), .B0(ori_ori_n962_), .B1(ori_ori_n88_), .Y(ori_ori_n964_));
  AOI210     o0936(.A0(ori_ori_n422_), .A1(ori_ori_n37_), .B0(ori_ori_n964_), .Y(ori_ori_n965_));
  NO2        o0937(.A(ori_ori_n141_), .B(ori_ori_n80_), .Y(ori_ori_n966_));
  OR2        o0938(.A(ori_ori_n966_), .B(ori_ori_n559_), .Y(ori_ori_n967_));
  NA2        o0939(.A(ori_ori_n560_), .B(ori_ori_n384_), .Y(ori_ori_n968_));
  AOI210     o0940(.A0(ori_ori_n968_), .A1(n), .B0(ori_ori_n967_), .Y(ori_ori_n969_));
  OAI220     o0941(.A0(ori_ori_n969_), .A1(ori_ori_n961_), .B0(ori_ori_n965_), .B1(ori_ori_n332_), .Y(ori_ori_n970_));
  NO2        o0942(.A(ori_ori_n662_), .B(ori_ori_n506_), .Y(ori_ori_n971_));
  NA3        o0943(.A(ori_ori_n343_), .B(ori_ori_n629_), .C(i), .Y(ori_ori_n972_));
  OAI210     o0944(.A0(ori_ori_n442_), .A1(ori_ori_n309_), .B0(ori_ori_n972_), .Y(ori_ori_n973_));
  OAI220     o0945(.A0(ori_ori_n973_), .A1(ori_ori_n971_), .B0(ori_ori_n678_), .B1(ori_ori_n754_), .Y(ori_ori_n974_));
  NA2        o0946(.A(ori_ori_n610_), .B(ori_ori_n110_), .Y(ori_ori_n975_));
  OR3        o0947(.A(ori_ori_n309_), .B(ori_ori_n438_), .C(f), .Y(ori_ori_n976_));
  NA3        o0948(.A(ori_ori_n629_), .B(ori_ori_n76_), .C(i), .Y(ori_ori_n977_));
  OA220      o0949(.A0(ori_ori_n977_), .A1(ori_ori_n975_), .B0(ori_ori_n976_), .B1(ori_ori_n596_), .Y(ori_ori_n978_));
  NA3        o0950(.A(ori_ori_n324_), .B(ori_ori_n114_), .C(o), .Y(ori_ori_n979_));
  AOI210     o0951(.A0(ori_ori_n675_), .A1(ori_ori_n979_), .B0(m), .Y(ori_ori_n980_));
  OAI210     o0952(.A0(ori_ori_n980_), .A1(ori_ori_n927_), .B0(ori_ori_n323_), .Y(ori_ori_n981_));
  NA2        o0953(.A(ori_ori_n694_), .B(ori_ori_n871_), .Y(ori_ori_n982_));
  NA2        o0954(.A(ori_ori_n834_), .B(ori_ori_n443_), .Y(ori_ori_n983_));
  NA2        o0955(.A(ori_ori_n221_), .B(ori_ori_n73_), .Y(ori_ori_n984_));
  NA2        o0956(.A(ori_ori_n984_), .B(ori_ori_n977_), .Y(ori_ori_n985_));
  AOI220     o0957(.A0(ori_ori_n985_), .A1(ori_ori_n258_), .B0(ori_ori_n983_), .B1(ori_ori_n982_), .Y(ori_ori_n986_));
  NA4        o0958(.A(ori_ori_n986_), .B(ori_ori_n981_), .C(ori_ori_n978_), .D(ori_ori_n974_), .Y(ori_ori_n987_));
  NO2        o0959(.A(ori_ori_n380_), .B(ori_ori_n87_), .Y(ori_ori_n988_));
  OAI210     o0960(.A0(ori_ori_n988_), .A1(ori_ori_n935_), .B0(ori_ori_n237_), .Y(ori_ori_n989_));
  NA2        o0961(.A(ori_ori_n664_), .B(ori_ori_n84_), .Y(ori_ori_n990_));
  NO2        o0962(.A(ori_ori_n466_), .B(ori_ori_n213_), .Y(ori_ori_n991_));
  AOI220     o0963(.A0(ori_ori_n991_), .A1(ori_ori_n385_), .B0(ori_ori_n940_), .B1(ori_ori_n217_), .Y(ori_ori_n992_));
  AOI220     o0964(.A0(ori_ori_n928_), .A1(ori_ori_n937_), .B0(ori_ori_n595_), .B1(ori_ori_n86_), .Y(ori_ori_n993_));
  NA4        o0965(.A(ori_ori_n993_), .B(ori_ori_n992_), .C(ori_ori_n990_), .D(ori_ori_n989_), .Y(ori_ori_n994_));
  OAI210     o0966(.A0(ori_ori_n983_), .A1(ori_ori_n936_), .B0(ori_ori_n548_), .Y(ori_ori_n995_));
  NA2        o0967(.A(ori_ori_n980_), .B(ori_ori_n926_), .Y(ori_ori_n996_));
  NA2        o0968(.A(ori_ori_n646_), .B(ori_ori_n539_), .Y(ori_ori_n997_));
  NA3        o0969(.A(ori_ori_n997_), .B(ori_ori_n996_), .C(ori_ori_n995_), .Y(ori_ori_n998_));
  NO4        o0970(.A(ori_ori_n998_), .B(ori_ori_n994_), .C(ori_ori_n987_), .D(ori_ori_n970_), .Y(ori_ori_n999_));
  NAi31      o0971(.An(ori_ori_n137_), .B(ori_ori_n424_), .C(n), .Y(ori_ori_n1000_));
  NO3        o0972(.A(ori_ori_n121_), .B(ori_ori_n341_), .C(ori_ori_n841_), .Y(ori_ori_n1001_));
  NO2        o0973(.A(ori_ori_n1001_), .B(ori_ori_n1000_), .Y(ori_ori_n1002_));
  NO3        o0974(.A(ori_ori_n269_), .B(ori_ori_n137_), .C(ori_ori_n411_), .Y(ori_ori_n1003_));
  AOI210     o0975(.A0(ori_ori_n1003_), .A1(ori_ori_n507_), .B0(ori_ori_n1002_), .Y(ori_ori_n1004_));
  NA2        o0976(.A(ori_ori_n500_), .B(i), .Y(ori_ori_n1005_));
  NA2        o0977(.A(ori_ori_n1005_), .B(ori_ori_n1004_), .Y(ori_ori_n1006_));
  NA2        o0978(.A(ori_ori_n230_), .B(ori_ori_n169_), .Y(ori_ori_n1007_));
  NO3        o0979(.A(ori_ori_n307_), .B(ori_ori_n448_), .C(ori_ori_n173_), .Y(ori_ori_n1008_));
  NOi31      o0980(.An(ori_ori_n1007_), .B(ori_ori_n1008_), .C(ori_ori_n213_), .Y(ori_ori_n1009_));
  NAi21      o0981(.An(ori_ori_n560_), .B(ori_ori_n991_), .Y(ori_ori_n1010_));
  NA2        o0982(.A(ori_ori_n491_), .B(o), .Y(ori_ori_n1011_));
  NA2        o0983(.A(ori_ori_n1011_), .B(ori_ori_n1010_), .Y(ori_ori_n1012_));
  NO2        o0984(.A(ori_ori_n1000_), .B(ori_ori_n233_), .Y(ori_ori_n1013_));
  NA2        o0985(.A(ori_ori_n931_), .B(ori_ori_n922_), .Y(ori_ori_n1014_));
  OAI220     o0986(.A0(ori_ori_n928_), .A1(ori_ori_n936_), .B0(ori_ori_n550_), .B1(ori_ori_n432_), .Y(ori_ori_n1015_));
  NA3        o0987(.A(ori_ori_n1015_), .B(ori_ori_n1014_), .C(ori_ori_n623_), .Y(ori_ori_n1016_));
  OAI210     o0988(.A0(ori_ori_n931_), .A1(ori_ori_n923_), .B0(ori_ori_n1007_), .Y(ori_ori_n1017_));
  NA3        o0989(.A(ori_ori_n968_), .B(ori_ori_n496_), .C(ori_ori_n46_), .Y(ori_ori_n1018_));
  AOI210     o0990(.A0(ori_ori_n383_), .A1(ori_ori_n381_), .B0(ori_ori_n331_), .Y(ori_ori_n1019_));
  NA3        o0991(.A(ori_ori_n1019_), .B(ori_ori_n1018_), .C(ori_ori_n1017_), .Y(ori_ori_n1020_));
  OR3        o0992(.A(ori_ori_n1020_), .B(ori_ori_n1016_), .C(ori_ori_n1013_), .Y(ori_ori_n1021_));
  NO4        o0993(.A(ori_ori_n1021_), .B(ori_ori_n1012_), .C(ori_ori_n1009_), .D(ori_ori_n1006_), .Y(ori_ori_n1022_));
  NA4        o0994(.A(ori_ori_n1022_), .B(ori_ori_n999_), .C(ori_ori_n960_), .D(ori_ori_n947_), .Y(ori13));
  AN2        o0995(.A(c), .B(b), .Y(ori_ori_n1024_));
  NAi32      o0996(.An(d), .Bn(c), .C(e), .Y(ori_ori_n1025_));
  AN2        o0997(.A(d), .B(c), .Y(ori_ori_n1026_));
  NA2        o0998(.A(ori_ori_n1026_), .B(ori_ori_n112_), .Y(ori_ori_n1027_));
  NOi41      o0999(.An(n), .B(m), .C(i), .D(h), .Y(ori_ori_n1028_));
  NA3        o1000(.A(k), .B(j), .C(i), .Y(ori_ori_n1029_));
  OR3        o1001(.A(n), .B(m), .C(i), .Y(ori_ori_n1030_));
  AN3        o1002(.A(o), .B(f), .C(c), .Y(ori_ori_n1031_));
  NA3        o1003(.A(ori_ori_n1031_), .B(ori_ori_n474_), .C(h), .Y(ori_ori_n1032_));
  NA3        o1004(.A(l), .B(k), .C(j), .Y(ori_ori_n1033_));
  NA2        o1005(.A(i), .B(h), .Y(ori_ori_n1034_));
  NO3        o1006(.A(ori_ori_n1034_), .B(ori_ori_n1033_), .C(ori_ori_n128_), .Y(ori_ori_n1035_));
  NO3        o1007(.A(ori_ori_n138_), .B(ori_ori_n281_), .C(ori_ori_n213_), .Y(ori_ori_n1036_));
  NA3        o1008(.A(c), .B(b), .C(a), .Y(ori_ori_n1037_));
  NO2        o1009(.A(ori_ori_n535_), .B(ori_ori_n603_), .Y(ori_ori_n1038_));
  NA4        o1010(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(o), .D(ori_ori_n212_), .Y(ori_ori_n1039_));
  NA4        o1011(.A(ori_ori_n581_), .B(m), .C(ori_ori_n109_), .D(ori_ori_n212_), .Y(ori_ori_n1040_));
  NA3        o1012(.A(ori_ori_n1040_), .B(ori_ori_n373_), .C(ori_ori_n1039_), .Y(ori_ori_n1041_));
  NO2        o1013(.A(ori_ori_n1041_), .B(ori_ori_n1038_), .Y(ori_ori_n1042_));
  NOi41      o1014(.An(ori_ori_n801_), .B(ori_ori_n846_), .C(ori_ori_n835_), .D(ori_ori_n721_), .Y(ori_ori_n1043_));
  OAI220     o1015(.A0(ori_ori_n1043_), .A1(ori_ori_n694_), .B0(ori_ori_n1042_), .B1(ori_ori_n594_), .Y(ori_ori_n1044_));
  NOi31      o1016(.An(m), .B(n), .C(f), .Y(ori_ori_n1045_));
  NA2        o1017(.A(ori_ori_n1045_), .B(ori_ori_n51_), .Y(ori_ori_n1046_));
  AN2        o1018(.A(e), .B(c), .Y(ori_ori_n1047_));
  NA2        o1019(.A(ori_ori_n1047_), .B(a), .Y(ori_ori_n1048_));
  OAI220     o1020(.A0(ori_ori_n1048_), .A1(ori_ori_n1046_), .B0(ori_ori_n879_), .B1(ori_ori_n431_), .Y(ori_ori_n1049_));
  NA2        o1021(.A(ori_ori_n516_), .B(l), .Y(ori_ori_n1050_));
  NO2        o1022(.A(ori_ori_n281_), .B(a), .Y(ori_ori_n1051_));
  NO2        o1023(.A(ori_ori_n83_), .B(o), .Y(ori_ori_n1052_));
  NO4        o1024(.A(ori_ori_n1049_), .B(ori_ori_n1044_), .C(ori_ori_n814_), .D(ori_ori_n570_), .Y(ori_ori_n1053_));
  NA2        o1025(.A(c), .B(b), .Y(ori_ori_n1054_));
  NO2        o1026(.A(ori_ori_n706_), .B(ori_ori_n1054_), .Y(ori_ori_n1055_));
  OAI210     o1027(.A0(ori_ori_n855_), .A1(ori_ori_n826_), .B0(ori_ori_n418_), .Y(ori_ori_n1056_));
  OAI210     o1028(.A0(ori_ori_n1056_), .A1(ori_ori_n856_), .B0(ori_ori_n1055_), .Y(ori_ori_n1057_));
  NAi21      o1029(.An(ori_ori_n426_), .B(ori_ori_n1055_), .Y(ori_ori_n1058_));
  NA3        o1030(.A(ori_ori_n432_), .B(ori_ori_n565_), .C(f), .Y(ori_ori_n1059_));
  OAI210     o1031(.A0(ori_ori_n554_), .A1(ori_ori_n39_), .B0(ori_ori_n1051_), .Y(ori_ori_n1060_));
  NA3        o1032(.A(ori_ori_n1060_), .B(ori_ori_n1059_), .C(ori_ori_n1058_), .Y(ori_ori_n1061_));
  NA2        o1033(.A(ori_ori_n261_), .B(ori_ori_n115_), .Y(ori_ori_n1062_));
  OAI210     o1034(.A0(ori_ori_n1062_), .A1(ori_ori_n284_), .B0(o), .Y(ori_ori_n1063_));
  NAi21      o1035(.An(f), .B(d), .Y(ori_ori_n1064_));
  NO2        o1036(.A(ori_ori_n1064_), .B(ori_ori_n1037_), .Y(ori_ori_n1065_));
  INV        o1037(.A(ori_ori_n1065_), .Y(ori_ori_n1066_));
  AOI210     o1038(.A0(ori_ori_n1063_), .A1(ori_ori_n290_), .B0(ori_ori_n1066_), .Y(ori_ori_n1067_));
  AOI210     o1039(.A0(ori_ori_n1067_), .A1(ori_ori_n110_), .B0(ori_ori_n1061_), .Y(ori_ori_n1068_));
  NA2        o1040(.A(ori_ori_n477_), .B(ori_ori_n476_), .Y(ori_ori_n1069_));
  NO2        o1041(.A(ori_ori_n180_), .B(ori_ori_n236_), .Y(ori_ori_n1070_));
  NA2        o1042(.A(ori_ori_n1070_), .B(m), .Y(ori_ori_n1071_));
  NA3        o1043(.A(ori_ori_n911_), .B(ori_ori_n1050_), .C(ori_ori_n480_), .Y(ori_ori_n1072_));
  OAI210     o1044(.A0(ori_ori_n1072_), .A1(ori_ori_n310_), .B0(ori_ori_n478_), .Y(ori_ori_n1073_));
  AOI210     o1045(.A0(ori_ori_n1073_), .A1(ori_ori_n1069_), .B0(ori_ori_n1071_), .Y(ori_ori_n1074_));
  NA2        o1046(.A(ori_ori_n451_), .B(ori_ori_n1065_), .Y(ori_ori_n1075_));
  INV        o1047(.A(ori_ori_n1075_), .Y(ori_ori_n1076_));
  NO2        o1048(.A(ori_ori_n1076_), .B(ori_ori_n1074_), .Y(ori_ori_n1077_));
  NA4        o1049(.A(ori_ori_n1077_), .B(ori_ori_n1068_), .C(ori_ori_n1057_), .D(ori_ori_n1053_), .Y(ori00));
  NA2        o1050(.A(ori_ori_n892_), .B(ori_ori_n937_), .Y(ori_ori_n1079_));
  INV        o1051(.A(ori_ori_n718_), .Y(ori_ori_n1080_));
  NA2        o1052(.A(ori_ori_n1080_), .B(ori_ori_n1079_), .Y(ori_ori_n1081_));
  NA2        o1053(.A(ori_ori_n518_), .B(f), .Y(ori_ori_n1082_));
  OAI210     o1054(.A0(ori_ori_n1001_), .A1(ori_ori_n40_), .B0(ori_ori_n648_), .Y(ori_ori_n1083_));
  NA3        o1055(.A(ori_ori_n1083_), .B(ori_ori_n257_), .C(n), .Y(ori_ori_n1084_));
  AOI210     o1056(.A0(ori_ori_n1084_), .A1(ori_ori_n1082_), .B0(ori_ori_n1027_), .Y(ori_ori_n1085_));
  NO2        o1057(.A(ori_ori_n1085_), .B(ori_ori_n1081_), .Y(ori_ori_n1086_));
  NA3        o1058(.A(ori_ori_n165_), .B(ori_ori_n46_), .C(ori_ori_n45_), .Y(ori_ori_n1087_));
  NA3        o1059(.A(d), .B(ori_ori_n56_), .C(b), .Y(ori_ori_n1088_));
  NO2        o1060(.A(ori_ori_n1088_), .B(ori_ori_n1087_), .Y(ori_ori_n1089_));
  INV        o1061(.A(ori_ori_n583_), .Y(ori_ori_n1090_));
  NO3        o1062(.A(ori_ori_n1090_), .B(ori_ori_n1089_), .C(ori_ori_n914_), .Y(ori_ori_n1091_));
  NO4        o1063(.A(ori_ori_n497_), .B(ori_ori_n358_), .C(ori_ori_n1054_), .D(ori_ori_n59_), .Y(ori_ori_n1092_));
  NA3        o1064(.A(ori_ori_n386_), .B(ori_ori_n220_), .C(o), .Y(ori_ori_n1093_));
  OR2        o1065(.A(ori_ori_n1093_), .B(ori_ori_n1088_), .Y(ori_ori_n1094_));
  NO2        o1066(.A(h), .B(o), .Y(ori_ori_n1095_));
  NA4        o1067(.A(ori_ori_n507_), .B(ori_ori_n474_), .C(ori_ori_n1095_), .D(ori_ori_n1024_), .Y(ori_ori_n1096_));
  OAI220     o1068(.A0(ori_ori_n535_), .A1(ori_ori_n603_), .B0(ori_ori_n88_), .B1(ori_ori_n87_), .Y(ori_ori_n1097_));
  AOI220     o1069(.A0(ori_ori_n1097_), .A1(ori_ori_n543_), .B0(ori_ori_n942_), .B1(ori_ori_n582_), .Y(ori_ori_n1098_));
  AOI220     o1070(.A0(ori_ori_n316_), .A1(ori_ori_n246_), .B0(ori_ori_n175_), .B1(ori_ori_n145_), .Y(ori_ori_n1099_));
  NA4        o1071(.A(ori_ori_n1099_), .B(ori_ori_n1098_), .C(ori_ori_n1096_), .D(ori_ori_n1094_), .Y(ori_ori_n1100_));
  NO3        o1072(.A(ori_ori_n1100_), .B(ori_ori_n1092_), .C(ori_ori_n264_), .Y(ori_ori_n1101_));
  INV        o1073(.A(ori_ori_n321_), .Y(ori_ori_n1102_));
  AOI210     o1074(.A0(ori_ori_n246_), .A1(ori_ori_n348_), .B0(ori_ori_n585_), .Y(ori_ori_n1103_));
  NA3        o1075(.A(ori_ori_n1103_), .B(ori_ori_n1102_), .C(ori_ori_n151_), .Y(ori_ori_n1104_));
  NO2        o1076(.A(ori_ori_n238_), .B(ori_ori_n179_), .Y(ori_ori_n1105_));
  NA2        o1077(.A(ori_ori_n1105_), .B(ori_ori_n432_), .Y(ori_ori_n1106_));
  INV        o1078(.A(ori_ori_n1106_), .Y(ori_ori_n1107_));
  NO2        o1079(.A(ori_ori_n272_), .B(ori_ori_n69_), .Y(ori_ori_n1108_));
  NO3        o1080(.A(ori_ori_n431_), .B(ori_ori_n822_), .C(n), .Y(ori_ori_n1109_));
  NA2        o1081(.A(ori_ori_n1109_), .B(ori_ori_n1108_), .Y(ori_ori_n1110_));
  INV        o1082(.A(ori_ori_n1110_), .Y(ori_ori_n1111_));
  NO4        o1083(.A(ori_ori_n1111_), .B(ori_ori_n1107_), .C(ori_ori_n1104_), .D(ori_ori_n527_), .Y(ori_ori_n1112_));
  AN3        o1084(.A(ori_ori_n1112_), .B(ori_ori_n1101_), .C(ori_ori_n1091_), .Y(ori_ori_n1113_));
  NA2        o1085(.A(ori_ori_n543_), .B(ori_ori_n98_), .Y(ori_ori_n1114_));
  NA3        o1086(.A(ori_ori_n1045_), .B(ori_ori_n610_), .C(ori_ori_n473_), .Y(ori_ori_n1115_));
  NA3        o1087(.A(ori_ori_n1115_), .B(ori_ori_n1114_), .C(ori_ori_n240_), .Y(ori_ori_n1116_));
  NA2        o1088(.A(ori_ori_n1041_), .B(ori_ori_n543_), .Y(ori_ori_n1117_));
  NA4        o1089(.A(ori_ori_n651_), .B(ori_ori_n204_), .C(ori_ori_n220_), .D(ori_ori_n160_), .Y(ori_ori_n1118_));
  NA3        o1090(.A(ori_ori_n1118_), .B(ori_ori_n1117_), .C(ori_ori_n294_), .Y(ori_ori_n1119_));
  OAI210     o1091(.A0(ori_ori_n472_), .A1(ori_ori_n116_), .B0(ori_ori_n858_), .Y(ori_ori_n1120_));
  NA2        o1092(.A(ori_ori_n1120_), .B(ori_ori_n1072_), .Y(ori_ori_n1121_));
  NO2        o1093(.A(ori_ori_n216_), .B(ori_ori_n213_), .Y(ori_ori_n1122_));
  NA2        o1094(.A(n), .B(e), .Y(ori_ori_n1123_));
  NO2        o1095(.A(ori_ori_n1123_), .B(ori_ori_n143_), .Y(ori_ori_n1124_));
  AOI220     o1096(.A0(ori_ori_n1124_), .A1(ori_ori_n270_), .B0(ori_ori_n839_), .B1(ori_ori_n1122_), .Y(ori_ori_n1125_));
  OAI210     o1097(.A0(ori_ori_n359_), .A1(ori_ori_n311_), .B0(ori_ori_n453_), .Y(ori_ori_n1126_));
  NA3        o1098(.A(ori_ori_n1126_), .B(ori_ori_n1125_), .C(ori_ori_n1121_), .Y(ori_ori_n1127_));
  NA2        o1099(.A(ori_ori_n1124_), .B(ori_ori_n843_), .Y(ori_ori_n1128_));
  AOI220     o1100(.A0(ori_ori_n951_), .A1(ori_ori_n582_), .B0(ori_ori_n651_), .B1(ori_ori_n243_), .Y(ori_ori_n1129_));
  NO2        o1101(.A(ori_ori_n64_), .B(h), .Y(ori_ori_n1130_));
  NA3        o1102(.A(ori_ori_n1129_), .B(ori_ori_n1128_), .C(ori_ori_n860_), .Y(ori_ori_n1131_));
  NO4        o1103(.A(ori_ori_n1131_), .B(ori_ori_n1127_), .C(ori_ori_n1119_), .D(ori_ori_n1116_), .Y(ori_ori_n1132_));
  NA2        o1104(.A(ori_ori_n827_), .B(ori_ori_n753_), .Y(ori_ori_n1133_));
  NA4        o1105(.A(ori_ori_n1133_), .B(ori_ori_n1132_), .C(ori_ori_n1113_), .D(ori_ori_n1086_), .Y(ori01));
  NO2        o1106(.A(ori_ori_n488_), .B(ori_ori_n279_), .Y(ori_ori_n1135_));
  NA2        o1107(.A(ori_ori_n397_), .B(i), .Y(ori_ori_n1136_));
  NA3        o1108(.A(ori_ori_n1136_), .B(ori_ori_n1135_), .C(ori_ori_n1014_), .Y(ori_ori_n1137_));
  NA2        o1109(.A(ori_ori_n595_), .B(ori_ori_n86_), .Y(ori_ori_n1138_));
  NA2        o1110(.A(ori_ori_n560_), .B(ori_ori_n268_), .Y(ori_ori_n1139_));
  NA2        o1111(.A(ori_ori_n956_), .B(ori_ori_n1139_), .Y(ori_ori_n1140_));
  NA4        o1112(.A(ori_ori_n1140_), .B(ori_ori_n1138_), .C(ori_ori_n907_), .D(ori_ori_n333_), .Y(ori_ori_n1141_));
  NA2        o1113(.A(ori_ori_n45_), .B(f), .Y(ori_ori_n1142_));
  NA2        o1114(.A(ori_ori_n713_), .B(ori_ori_n93_), .Y(ori_ori_n1143_));
  NO2        o1115(.A(ori_ori_n1143_), .B(ori_ori_n1142_), .Y(ori_ori_n1144_));
  OAI210     o1116(.A0(ori_ori_n780_), .A1(ori_ori_n606_), .B0(ori_ori_n1118_), .Y(ori_ori_n1145_));
  AOI210     o1117(.A0(ori_ori_n1144_), .A1(ori_ori_n636_), .B0(ori_ori_n1145_), .Y(ori_ori_n1146_));
  OR2        o1118(.A(ori_ori_n663_), .B(ori_ori_n373_), .Y(ori_ori_n1147_));
  NAi41      o1119(.An(ori_ori_n159_), .B(ori_ori_n1147_), .C(ori_ori_n1146_), .D(ori_ori_n891_), .Y(ori_ori_n1148_));
  NO3        o1120(.A(ori_ori_n781_), .B(ori_ori_n677_), .C(ori_ori_n521_), .Y(ori_ori_n1149_));
  NA4        o1121(.A(ori_ori_n713_), .B(ori_ori_n93_), .C(ori_ori_n45_), .D(ori_ori_n212_), .Y(ori_ori_n1150_));
  OA220      o1122(.A0(ori_ori_n1150_), .A1(ori_ori_n671_), .B0(ori_ori_n193_), .B1(ori_ori_n191_), .Y(ori_ori_n1151_));
  NA3        o1123(.A(ori_ori_n1151_), .B(ori_ori_n1149_), .C(ori_ori_n133_), .Y(ori_ori_n1152_));
  NO4        o1124(.A(ori_ori_n1152_), .B(ori_ori_n1148_), .C(ori_ori_n1141_), .D(ori_ori_n1137_), .Y(ori_ori_n1153_));
  INV        o1125(.A(ori_ori_n1093_), .Y(ori_ori_n1154_));
  OAI210     o1126(.A0(ori_ori_n1154_), .A1(ori_ori_n300_), .B0(ori_ori_n539_), .Y(ori_ori_n1155_));
  AOI210     o1127(.A0(ori_ori_n202_), .A1(ori_ori_n85_), .B0(ori_ori_n212_), .Y(ori_ori_n1156_));
  OAI210     o1128(.A0(ori_ori_n804_), .A1(ori_ori_n432_), .B0(ori_ori_n1156_), .Y(ori_ori_n1157_));
  AN3        o1129(.A(m), .B(l), .C(k), .Y(ori_ori_n1158_));
  OAI210     o1130(.A0(ori_ori_n361_), .A1(ori_ori_n34_), .B0(ori_ori_n1158_), .Y(ori_ori_n1159_));
  NA2        o1131(.A(ori_ori_n201_), .B(ori_ori_n34_), .Y(ori_ori_n1160_));
  AO210      o1132(.A0(ori_ori_n1160_), .A1(ori_ori_n1159_), .B0(ori_ori_n332_), .Y(ori_ori_n1161_));
  NA3        o1133(.A(ori_ori_n1161_), .B(ori_ori_n1157_), .C(ori_ori_n1155_), .Y(ori_ori_n1162_));
  NA2        o1134(.A(ori_ori_n601_), .B(ori_ori_n114_), .Y(ori_ori_n1163_));
  INV        o1135(.A(ori_ori_n1163_), .Y(ori_ori_n1164_));
  NA2        o1136(.A(ori_ori_n278_), .B(ori_ori_n193_), .Y(ori_ori_n1165_));
  OAI210     o1137(.A0(ori_ori_n1165_), .A1(ori_ori_n388_), .B0(ori_ori_n667_), .Y(ori_ori_n1166_));
  OAI210     o1138(.A0(ori_ori_n1144_), .A1(ori_ori_n326_), .B0(ori_ori_n678_), .Y(ori_ori_n1167_));
  NA3        o1139(.A(ori_ori_n1167_), .B(ori_ori_n1166_), .C(ori_ori_n784_), .Y(ori_ori_n1168_));
  NO3        o1140(.A(ori_ori_n1168_), .B(ori_ori_n1164_), .C(ori_ori_n1162_), .Y(ori_ori_n1169_));
  NA3        o1141(.A(ori_ori_n607_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n1170_));
  NO2        o1142(.A(ori_ori_n1170_), .B(ori_ori_n202_), .Y(ori_ori_n1171_));
  AOI210     o1143(.A0(ori_ori_n514_), .A1(ori_ori_n58_), .B0(ori_ori_n1171_), .Y(ori_ori_n1172_));
  OR3        o1144(.A(ori_ori_n1143_), .B(ori_ori_n608_), .C(ori_ori_n1142_), .Y(ori_ori_n1173_));
  NO2        o1145(.A(ori_ori_n1150_), .B(ori_ori_n975_), .Y(ori_ori_n1174_));
  NO2        o1146(.A(ori_ori_n205_), .B(ori_ori_n108_), .Y(ori_ori_n1175_));
  NO3        o1147(.A(ori_ori_n1175_), .B(ori_ori_n1174_), .C(ori_ori_n1089_), .Y(ori_ori_n1176_));
  NA4        o1148(.A(ori_ori_n1176_), .B(ori_ori_n1173_), .C(ori_ori_n1172_), .D(ori_ori_n752_), .Y(ori_ori_n1177_));
  NO2        o1149(.A(ori_ori_n962_), .B(ori_ori_n232_), .Y(ori_ori_n1178_));
  NO2        o1150(.A(ori_ori_n963_), .B(ori_ori_n562_), .Y(ori_ori_n1179_));
  OAI210     o1151(.A0(ori_ori_n1179_), .A1(ori_ori_n1178_), .B0(ori_ori_n341_), .Y(ori_ori_n1180_));
  NA2        o1152(.A(ori_ori_n577_), .B(ori_ori_n575_), .Y(ori_ori_n1181_));
  NO3        o1153(.A(ori_ori_n75_), .B(ori_ori_n298_), .C(ori_ori_n45_), .Y(ori_ori_n1182_));
  NA2        o1154(.A(ori_ori_n1182_), .B(ori_ori_n559_), .Y(ori_ori_n1183_));
  NA3        o1155(.A(ori_ori_n1183_), .B(ori_ori_n1181_), .C(ori_ori_n673_), .Y(ori_ori_n1184_));
  OR2        o1156(.A(ori_ori_n1093_), .B(ori_ori_n1088_), .Y(ori_ori_n1185_));
  NO2        o1157(.A(ori_ori_n373_), .B(ori_ori_n68_), .Y(ori_ori_n1186_));
  INV        o1158(.A(ori_ori_n1186_), .Y(ori_ori_n1187_));
  NA2        o1159(.A(ori_ori_n1182_), .B(ori_ori_n807_), .Y(ori_ori_n1188_));
  NA4        o1160(.A(ori_ori_n1188_), .B(ori_ori_n1187_), .C(ori_ori_n1185_), .D(ori_ori_n389_), .Y(ori_ori_n1189_));
  NOi41      o1161(.An(ori_ori_n1180_), .B(ori_ori_n1189_), .C(ori_ori_n1184_), .D(ori_ori_n1177_), .Y(ori_ori_n1190_));
  NO2        o1162(.A(ori_ori_n127_), .B(ori_ori_n45_), .Y(ori_ori_n1191_));
  NO2        o1163(.A(ori_ori_n45_), .B(ori_ori_n40_), .Y(ori_ori_n1192_));
  AO220      o1164(.A0(ori_ori_n1192_), .A1(ori_ori_n626_), .B0(ori_ori_n1191_), .B1(ori_ori_n711_), .Y(ori_ori_n1193_));
  NA2        o1165(.A(ori_ori_n1193_), .B(ori_ori_n341_), .Y(ori_ori_n1194_));
  INV        o1166(.A(ori_ori_n131_), .Y(ori_ori_n1195_));
  NO3        o1167(.A(ori_ori_n1034_), .B(ori_ori_n174_), .C(ori_ori_n83_), .Y(ori_ori_n1196_));
  AOI220     o1168(.A0(ori_ori_n1196_), .A1(ori_ori_n1195_), .B0(ori_ori_n1182_), .B1(ori_ori_n966_), .Y(ori_ori_n1197_));
  NA2        o1169(.A(ori_ori_n1197_), .B(ori_ori_n1194_), .Y(ori_ori_n1198_));
  NO2        o1170(.A(ori_ori_n618_), .B(ori_ori_n617_), .Y(ori_ori_n1199_));
  NO4        o1171(.A(ori_ori_n1034_), .B(ori_ori_n1199_), .C(ori_ori_n172_), .D(ori_ori_n83_), .Y(ori_ori_n1200_));
  NO3        o1172(.A(ori_ori_n1200_), .B(ori_ori_n1198_), .C(ori_ori_n640_), .Y(ori_ori_n1201_));
  NA4        o1173(.A(ori_ori_n1201_), .B(ori_ori_n1190_), .C(ori_ori_n1169_), .D(ori_ori_n1153_), .Y(ori06));
  NO2        o1174(.A(ori_ori_n224_), .B(ori_ori_n100_), .Y(ori_ori_n1203_));
  OAI210     o1175(.A0(ori_ori_n1203_), .A1(ori_ori_n1196_), .B0(ori_ori_n385_), .Y(ori_ori_n1204_));
  NO3        o1176(.A(ori_ori_n604_), .B(ori_ori_n802_), .C(ori_ori_n605_), .Y(ori_ori_n1205_));
  OR2        o1177(.A(ori_ori_n1205_), .B(ori_ori_n879_), .Y(ori_ori_n1206_));
  NA3        o1178(.A(ori_ori_n1206_), .B(ori_ori_n1204_), .C(ori_ori_n1180_), .Y(ori_ori_n1207_));
  NO3        o1179(.A(ori_ori_n1207_), .B(ori_ori_n1184_), .C(ori_ori_n256_), .Y(ori_ori_n1208_));
  NO2        o1180(.A(ori_ori_n298_), .B(ori_ori_n45_), .Y(ori_ori_n1209_));
  AOI210     o1181(.A0(ori_ori_n1209_), .A1(ori_ori_n967_), .B0(ori_ori_n1178_), .Y(ori_ori_n1210_));
  AOI210     o1182(.A0(ori_ori_n1209_), .A1(ori_ori_n563_), .B0(ori_ori_n1193_), .Y(ori_ori_n1211_));
  AOI210     o1183(.A0(ori_ori_n1211_), .A1(ori_ori_n1210_), .B0(ori_ori_n338_), .Y(ori_ori_n1212_));
  OAI210     o1184(.A0(ori_ori_n85_), .A1(ori_ori_n40_), .B0(ori_ori_n676_), .Y(ori_ori_n1213_));
  NA2        o1185(.A(ori_ori_n1213_), .B(ori_ori_n644_), .Y(ori_ori_n1214_));
  NO2        o1186(.A(ori_ori_n523_), .B(ori_ori_n169_), .Y(ori_ori_n1215_));
  NO2        o1187(.A(ori_ori_n611_), .B(ori_ori_n1046_), .Y(ori_ori_n1216_));
  OAI210     o1188(.A0(ori_ori_n467_), .A1(ori_ori_n247_), .B0(ori_ori_n902_), .Y(ori_ori_n1217_));
  NO3        o1189(.A(ori_ori_n1217_), .B(ori_ori_n1216_), .C(ori_ori_n1215_), .Y(ori_ori_n1218_));
  NO2        o1190(.A(ori_ori_n372_), .B(ori_ori_n132_), .Y(ori_ori_n1219_));
  NA2        o1191(.A(ori_ori_n1219_), .B(ori_ori_n595_), .Y(ori_ori_n1220_));
  NA3        o1192(.A(ori_ori_n1220_), .B(ori_ori_n1218_), .C(ori_ori_n1214_), .Y(ori_ori_n1221_));
  NO2        o1193(.A(ori_ori_n745_), .B(ori_ori_n371_), .Y(ori_ori_n1222_));
  NO2        o1194(.A(ori_ori_n678_), .B(ori_ori_n636_), .Y(ori_ori_n1223_));
  NOi21      o1195(.An(ori_ori_n1222_), .B(ori_ori_n1223_), .Y(ori_ori_n1224_));
  AN2        o1196(.A(ori_ori_n951_), .B(ori_ori_n647_), .Y(ori_ori_n1225_));
  NO4        o1197(.A(ori_ori_n1225_), .B(ori_ori_n1224_), .C(ori_ori_n1221_), .D(ori_ori_n1212_), .Y(ori_ori_n1226_));
  OAI220     o1198(.A0(ori_ori_n735_), .A1(ori_ori_n47_), .B0(ori_ori_n224_), .B1(ori_ori_n620_), .Y(ori_ori_n1227_));
  OAI210     o1199(.A0(ori_ori_n274_), .A1(c), .B0(ori_ori_n643_), .Y(ori_ori_n1228_));
  NA2        o1200(.A(ori_ori_n1228_), .B(ori_ori_n1227_), .Y(ori_ori_n1229_));
  NO3        o1201(.A(ori_ori_n242_), .B(ori_ori_n100_), .C(ori_ori_n281_), .Y(ori_ori_n1230_));
  OAI220     o1202(.A0(ori_ori_n703_), .A1(ori_ori_n247_), .B0(ori_ori_n520_), .B1(ori_ori_n523_), .Y(ori_ori_n1231_));
  OAI210     o1203(.A0(l), .A1(i), .B0(k), .Y(ori_ori_n1232_));
  NO3        o1204(.A(ori_ori_n1232_), .B(ori_ori_n603_), .C(j), .Y(ori_ori_n1233_));
  NO3        o1205(.A(ori_ori_n1231_), .B(ori_ori_n1230_), .C(ori_ori_n1049_), .Y(ori_ori_n1234_));
  NA4        o1206(.A(ori_ori_n791_), .B(ori_ori_n790_), .C(ori_ori_n441_), .D(ori_ori_n871_), .Y(ori_ori_n1235_));
  NAi31      o1207(.An(ori_ori_n745_), .B(ori_ori_n1235_), .C(ori_ori_n201_), .Y(ori_ori_n1236_));
  NA4        o1208(.A(ori_ori_n1236_), .B(ori_ori_n1234_), .C(ori_ori_n1229_), .D(ori_ori_n1129_), .Y(ori_ori_n1237_));
  NOi21      o1209(.An(ori_ori_n1205_), .B(ori_ori_n471_), .Y(ori_ori_n1238_));
  OR3        o1210(.A(ori_ori_n1238_), .B(ori_ori_n780_), .C(ori_ori_n546_), .Y(ori_ori_n1239_));
  NA2        o1211(.A(ori_ori_n577_), .B(ori_ori_n453_), .Y(ori_ori_n1240_));
  NA2        o1212(.A(ori_ori_n1233_), .B(ori_ori_n787_), .Y(ori_ori_n1241_));
  NA3        o1213(.A(ori_ori_n1241_), .B(ori_ori_n1240_), .C(ori_ori_n1239_), .Y(ori_ori_n1242_));
  AOI220     o1214(.A0(ori_ori_n1222_), .A1(ori_ori_n753_), .B0(ori_ori_n1219_), .B1(ori_ori_n237_), .Y(ori_ori_n1243_));
  AN2        o1215(.A(ori_ori_n923_), .B(ori_ori_n922_), .Y(ori_ori_n1244_));
  NO4        o1216(.A(ori_ori_n1244_), .B(ori_ori_n869_), .C(ori_ori_n510_), .D(ori_ori_n491_), .Y(ori_ori_n1245_));
  NA3        o1217(.A(ori_ori_n1245_), .B(ori_ori_n1243_), .C(ori_ori_n1188_), .Y(ori_ori_n1246_));
  NAi21      o1218(.An(j), .B(i), .Y(ori_ori_n1247_));
  NO4        o1219(.A(ori_ori_n1199_), .B(ori_ori_n1247_), .C(ori_ori_n447_), .D(ori_ori_n234_), .Y(ori_ori_n1248_));
  NO4        o1220(.A(ori_ori_n1248_), .B(ori_ori_n1246_), .C(ori_ori_n1242_), .D(ori_ori_n1237_), .Y(ori_ori_n1249_));
  NA4        o1221(.A(ori_ori_n1249_), .B(ori_ori_n1226_), .C(ori_ori_n1208_), .D(ori_ori_n1201_), .Y(ori07));
  NAi32      o1222(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1251_));
  NO3        o1223(.A(ori_ori_n1251_), .B(o), .C(f), .Y(ori_ori_n1252_));
  NAi21      o1224(.An(f), .B(c), .Y(ori_ori_n1253_));
  NOi31      o1225(.An(n), .B(m), .C(b), .Y(ori_ori_n1254_));
  NOi41      o1226(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1255_));
  NO2        o1227(.A(k), .B(i), .Y(ori_ori_n1256_));
  NA3        o1228(.A(ori_ori_n1256_), .B(ori_ori_n890_), .C(ori_ori_n177_), .Y(ori_ori_n1257_));
  NO2        o1229(.A(ori_ori_n1029_), .B(ori_ori_n306_), .Y(ori_ori_n1258_));
  NA2        o1230(.A(ori_ori_n547_), .B(ori_ori_n76_), .Y(ori_ori_n1259_));
  NA2        o1231(.A(ori_ori_n1130_), .B(ori_ori_n288_), .Y(ori_ori_n1260_));
  NA3        o1232(.A(ori_ori_n1260_), .B(ori_ori_n1259_), .C(ori_ori_n1257_), .Y(ori_ori_n1261_));
  NO2        o1233(.A(ori_ori_n1261_), .B(ori_ori_n1252_), .Y(ori_ori_n1262_));
  NO3        o1234(.A(e), .B(d), .C(c), .Y(ori_ori_n1263_));
  NO2        o1235(.A(ori_ori_n128_), .B(ori_ori_n213_), .Y(ori_ori_n1264_));
  NA2        o1236(.A(ori_ori_n1264_), .B(ori_ori_n1263_), .Y(ori_ori_n1265_));
  NO2        o1237(.A(ori_ori_n1265_), .B(c), .Y(ori_ori_n1266_));
  NO3        o1238(.A(n), .B(m), .C(i), .Y(ori_ori_n1267_));
  NA3        o1239(.A(ori_ori_n700_), .B(ori_ori_n686_), .C(ori_ori_n109_), .Y(ori_ori_n1268_));
  NO2        o1240(.A(ori_ori_n1268_), .B(ori_ori_n45_), .Y(ori_ori_n1269_));
  INV        o1241(.A(ori_ori_n1267_), .Y(ori_ori_n1270_));
  NO2        o1242(.A(l), .B(k), .Y(ori_ori_n1271_));
  NO2        o1243(.A(ori_ori_n1269_), .B(ori_ori_n1266_), .Y(ori_ori_n1272_));
  NO2        o1244(.A(o), .B(c), .Y(ori_ori_n1273_));
  NO2        o1245(.A(ori_ori_n458_), .B(a), .Y(ori_ori_n1274_));
  NA2        o1246(.A(ori_ori_n1274_), .B(ori_ori_n110_), .Y(ori_ori_n1275_));
  NA2        o1247(.A(ori_ori_n134_), .B(ori_ori_n220_), .Y(ori_ori_n1276_));
  NO2        o1248(.A(ori_ori_n1276_), .B(ori_ori_n1380_), .Y(ori_ori_n1277_));
  NO2        o1249(.A(ori_ori_n751_), .B(ori_ori_n185_), .Y(ori_ori_n1278_));
  NOi31      o1250(.An(m), .B(n), .C(b), .Y(ori_ori_n1279_));
  NOi31      o1251(.An(f), .B(d), .C(c), .Y(ori_ori_n1280_));
  NA2        o1252(.A(ori_ori_n1280_), .B(ori_ori_n1279_), .Y(ori_ori_n1281_));
  INV        o1253(.A(ori_ori_n1281_), .Y(ori_ori_n1282_));
  NO3        o1254(.A(ori_ori_n1282_), .B(ori_ori_n1278_), .C(ori_ori_n1277_), .Y(ori_ori_n1283_));
  NA2        o1255(.A(ori_ori_n1031_), .B(ori_ori_n474_), .Y(ori_ori_n1284_));
  NO3        o1256(.A(ori_ori_n1284_), .B(ori_ori_n447_), .C(ori_ori_n45_), .Y(ori_ori_n1285_));
  NO3        o1257(.A(ori_ori_n41_), .B(i), .C(h), .Y(ori_ori_n1286_));
  NO2        o1258(.A(ori_ori_n1028_), .B(ori_ori_n1285_), .Y(ori_ori_n1287_));
  AN3        o1259(.A(ori_ori_n1287_), .B(ori_ori_n1283_), .C(ori_ori_n1275_), .Y(ori_ori_n1288_));
  NA2        o1260(.A(ori_ori_n1254_), .B(ori_ori_n382_), .Y(ori_ori_n1289_));
  INV        o1261(.A(ori_ori_n1289_), .Y(ori_ori_n1290_));
  INV        o1262(.A(ori_ori_n1035_), .Y(ori_ori_n1291_));
  NAi21      o1263(.An(ori_ori_n1290_), .B(ori_ori_n1291_), .Y(ori_ori_n1292_));
  NO4        o1264(.A(ori_ori_n128_), .B(o), .C(f), .D(e), .Y(ori_ori_n1293_));
  NA2        o1265(.A(ori_ori_n1255_), .B(ori_ori_n1271_), .Y(ori_ori_n1294_));
  INV        o1266(.A(ori_ori_n1294_), .Y(ori_ori_n1295_));
  OR3        o1267(.A(ori_ori_n546_), .B(ori_ori_n545_), .C(ori_ori_n109_), .Y(ori_ori_n1296_));
  NA2        o1268(.A(ori_ori_n1045_), .B(ori_ori_n411_), .Y(ori_ori_n1297_));
  NO2        o1269(.A(ori_ori_n1297_), .B(ori_ori_n440_), .Y(ori_ori_n1298_));
  AO210      o1270(.A0(ori_ori_n1298_), .A1(ori_ori_n112_), .B0(ori_ori_n1295_), .Y(ori_ori_n1299_));
  NO2        o1271(.A(ori_ori_n1299_), .B(ori_ori_n1292_), .Y(ori_ori_n1300_));
  NA4        o1272(.A(ori_ori_n1300_), .B(ori_ori_n1288_), .C(ori_ori_n1272_), .D(ori_ori_n1262_), .Y(ori_ori_n1301_));
  NO2        o1273(.A(ori_ori_n1054_), .B(ori_ori_n107_), .Y(ori_ori_n1302_));
  NA2        o1274(.A(ori_ori_n382_), .B(ori_ori_n56_), .Y(ori_ori_n1303_));
  NO2        o1275(.A(ori_ori_n1303_), .B(ori_ori_n1270_), .Y(ori_ori_n1304_));
  NA2        o1276(.A(ori_ori_n214_), .B(ori_ori_n177_), .Y(ori_ori_n1305_));
  NO2        o1277(.A(ori_ori_n1305_), .B(ori_ori_n1303_), .Y(ori_ori_n1306_));
  NO2        o1278(.A(ori_ori_n1032_), .B(ori_ori_n1030_), .Y(ori_ori_n1307_));
  NO3        o1279(.A(ori_ori_n1307_), .B(ori_ori_n1306_), .C(ori_ori_n1304_), .Y(ori_ori_n1308_));
  NO2        o1280(.A(ori_ori_n394_), .B(j), .Y(ori_ori_n1309_));
  NA2        o1281(.A(ori_ori_n1286_), .B(ori_ori_n1045_), .Y(ori_ori_n1310_));
  INV        o1282(.A(ori_ori_n1310_), .Y(ori_ori_n1311_));
  NA3        o1283(.A(o), .B(ori_ori_n1309_), .C(ori_ori_n156_), .Y(ori_ori_n1312_));
  INV        o1284(.A(ori_ori_n1312_), .Y(ori_ori_n1313_));
  NO2        o1285(.A(ori_ori_n745_), .B(ori_ori_n172_), .Y(ori_ori_n1314_));
  NO3        o1286(.A(ori_ori_n1314_), .B(ori_ori_n1313_), .C(ori_ori_n1311_), .Y(ori_ori_n1315_));
  INV        o1287(.A(ori_ori_n49_), .Y(ori_ori_n1316_));
  NA2        o1288(.A(ori_ori_n1316_), .B(ori_ori_n1095_), .Y(ori_ori_n1317_));
  INV        o1289(.A(ori_ori_n1317_), .Y(ori_ori_n1318_));
  NO2        o1290(.A(ori_ori_n668_), .B(ori_ori_n174_), .Y(ori_ori_n1319_));
  NO2        o1291(.A(ori_ori_n1319_), .B(ori_ori_n1318_), .Y(ori_ori_n1320_));
  NO3        o1292(.A(ori_ori_n1037_), .B(d), .C(ori_ori_n49_), .Y(ori_ori_n1321_));
  NO2        o1293(.A(ori_ori_n1030_), .B(h), .Y(ori_ori_n1322_));
  NA3        o1294(.A(ori_ori_n1302_), .B(ori_ori_n474_), .C(f), .Y(ori_ori_n1323_));
  INV        o1295(.A(ori_ori_n177_), .Y(ori_ori_n1324_));
  NO2        o1296(.A(ori_ori_n1378_), .B(ori_ori_n1323_), .Y(ori_ori_n1325_));
  NO2        o1297(.A(ori_ori_n1247_), .B(ori_ori_n172_), .Y(ori_ori_n1326_));
  NOi21      o1298(.An(d), .B(f), .Y(ori_ori_n1327_));
  NO2        o1299(.A(ori_ori_n1325_), .B(ori_ori_n1322_), .Y(ori_ori_n1328_));
  NA4        o1300(.A(ori_ori_n1328_), .B(ori_ori_n1320_), .C(ori_ori_n1315_), .D(ori_ori_n1308_), .Y(ori_ori_n1329_));
  NA2        o1301(.A(h), .B(ori_ori_n1258_), .Y(ori_ori_n1330_));
  OAI210     o1302(.A0(ori_ori_n1293_), .A1(ori_ori_n1254_), .B0(ori_ori_n876_), .Y(ori_ori_n1331_));
  NO2        o1303(.A(ori_ori_n1025_), .B(ori_ori_n128_), .Y(ori_ori_n1332_));
  NA2        o1304(.A(ori_ori_n1332_), .B(ori_ori_n625_), .Y(ori_ori_n1333_));
  NA3        o1305(.A(ori_ori_n1333_), .B(ori_ori_n1331_), .C(ori_ori_n1330_), .Y(ori_ori_n1334_));
  NA2        o1306(.A(ori_ori_n1273_), .B(ori_ori_n1327_), .Y(ori_ori_n1335_));
  NO2        o1307(.A(ori_ori_n1335_), .B(m), .Y(ori_ori_n1336_));
  NO2        o1308(.A(ori_ori_n148_), .B(ori_ori_n179_), .Y(ori_ori_n1337_));
  OAI210     o1309(.A0(ori_ori_n1337_), .A1(ori_ori_n107_), .B0(ori_ori_n1279_), .Y(ori_ori_n1338_));
  INV        o1310(.A(ori_ori_n1338_), .Y(ori_ori_n1339_));
  NO3        o1311(.A(ori_ori_n1339_), .B(ori_ori_n1336_), .C(ori_ori_n1334_), .Y(ori_ori_n1340_));
  NO2        o1312(.A(ori_ori_n1253_), .B(e), .Y(ori_ori_n1341_));
  NA2        o1313(.A(ori_ori_n1341_), .B(ori_ori_n409_), .Y(ori_ori_n1342_));
  BUFFER     o1314(.A(ori_ori_n128_), .Y(ori_ori_n1343_));
  NO2        o1315(.A(ori_ori_n1343_), .B(ori_ori_n1342_), .Y(ori_ori_n1344_));
  NO2        o1316(.A(ori_ori_n1296_), .B(ori_ori_n355_), .Y(ori_ori_n1345_));
  NO2        o1317(.A(ori_ori_n1345_), .B(ori_ori_n1344_), .Y(ori_ori_n1346_));
  NO2        o1318(.A(ori_ori_n179_), .B(c), .Y(ori_ori_n1347_));
  NA2        o1319(.A(ori_ori_n1347_), .B(ori_ori_n177_), .Y(ori_ori_n1348_));
  AOI210     o1320(.A0(ori_ori_n540_), .A1(ori_ori_n371_), .B0(ori_ori_n1348_), .Y(ori_ori_n1349_));
  INV        o1321(.A(ori_ori_n1321_), .Y(ori_ori_n1350_));
  INV        o1322(.A(ori_ori_n1052_), .Y(ori_ori_n1351_));
  OAI220     o1323(.A0(ori_ori_n1351_), .A1(ori_ori_n65_), .B0(ori_ori_n1350_), .B1(ori_ori_n212_), .Y(ori_ori_n1352_));
  OR2        o1324(.A(h), .B(ori_ori_n545_), .Y(ori_ori_n1353_));
  NO2        o1325(.A(ori_ori_n1353_), .B(ori_ori_n172_), .Y(ori_ori_n1354_));
  NA2        o1326(.A(ori_ori_n1036_), .B(ori_ori_n220_), .Y(ori_ori_n1355_));
  NO2        o1327(.A(ori_ori_n49_), .B(l), .Y(ori_ori_n1356_));
  INV        o1328(.A(ori_ori_n493_), .Y(ori_ori_n1357_));
  NA2        o1329(.A(ori_ori_n1357_), .B(ori_ori_n1356_), .Y(ori_ori_n1358_));
  NA2        o1330(.A(ori_ori_n1358_), .B(ori_ori_n1355_), .Y(ori_ori_n1359_));
  NO4        o1331(.A(ori_ori_n1359_), .B(ori_ori_n1354_), .C(ori_ori_n1352_), .D(ori_ori_n1349_), .Y(ori_ori_n1360_));
  NA3        o1332(.A(ori_ori_n1360_), .B(ori_ori_n1346_), .C(ori_ori_n1340_), .Y(ori_ori_n1361_));
  NA3        o1333(.A(ori_ori_n955_), .B(ori_ori_n134_), .C(ori_ori_n46_), .Y(ori_ori_n1362_));
  INV        o1334(.A(ori_ori_n1362_), .Y(ori_ori_n1363_));
  NA2        o1335(.A(c), .B(ori_ori_n1322_), .Y(ori_ori_n1364_));
  NA2        o1336(.A(ori_ori_n1326_), .B(h), .Y(ori_ori_n1365_));
  NA2        o1337(.A(ori_ori_n1365_), .B(ori_ori_n1364_), .Y(ori_ori_n1366_));
  NO2        o1338(.A(ori_ori_n1366_), .B(ori_ori_n1363_), .Y(ori_ori_n1367_));
  INV        o1339(.A(ori_ori_n1341_), .Y(ori_ori_n1368_));
  NO2        o1340(.A(ori_ori_n1368_), .B(ori_ori_n1324_), .Y(ori_ori_n1369_));
  INV        o1341(.A(ori_ori_n1369_), .Y(ori_ori_n1370_));
  NOi31      o1342(.An(ori_ori_n30_), .B(m), .C(n), .Y(ori_ori_n1371_));
  INV        o1343(.A(ori_ori_n1371_), .Y(ori_ori_n1372_));
  NO2        o1344(.A(ori_ori_n1297_), .B(d), .Y(ori_ori_n1373_));
  NA4        o1345(.A(ori_ori_n1379_), .B(ori_ori_n1372_), .C(ori_ori_n1370_), .D(ori_ori_n1367_), .Y(ori_ori_n1374_));
  OR4        o1346(.A(ori_ori_n1374_), .B(ori_ori_n1361_), .C(ori_ori_n1329_), .D(ori_ori_n1301_), .Y(ori04));
  INV        o1347(.A(ori_ori_n110_), .Y(ori_ori_n1378_));
  INV        o1348(.A(ori_ori_n1373_), .Y(ori_ori_n1379_));
  INV        o1349(.A(h), .Y(ori_ori_n1380_));
  ZERO       o1350(.Y(ori02));
  ZERO       o1351(.Y(ori03));
  ZERO       o1352(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(m), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(m), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(m), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(m), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(m), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO4        m0025(.A(mai_mai_n53_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n54_));
  AOI210     m0026(.A0(mai_mai_n54_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NA3        m0031(.A(m), .B(mai_mai_n59_), .C(a), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(h), .Y(mai_mai_n61_));
  NAi31      m0033(.An(i), .B(l), .C(j), .Y(mai_mai_n62_));
  OAI220     m0034(.A0(mai_mai_n62_), .A1(mai_mai_n49_), .B0(mai_mai_n61_), .B1(mai_mai_n44_), .Y(mai_mai_n63_));
  NAi31      m0035(.An(mai_mai_n60_), .B(mai_mai_n63_), .C(mai_mai_n58_), .Y(mai_mai_n64_));
  NAi41      m0036(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n65_));
  NA2        m0037(.A(m), .B(f), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi21      m0039(.An(i), .B(j), .Y(mai_mai_n68_));
  NAi32      m0040(.An(n), .Bn(k), .C(m), .Y(mai_mai_n69_));
  NO2        m0041(.A(mai_mai_n69_), .B(mai_mai_n68_), .Y(mai_mai_n70_));
  NAi31      m0042(.An(l), .B(m), .C(k), .Y(mai_mai_n71_));
  NAi21      m0043(.An(e), .B(h), .Y(mai_mai_n72_));
  NAi41      m0044(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n74_));
  INV        m0046(.A(m), .Y(mai_mai_n75_));
  NOi21      m0047(.An(k), .B(l), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n77_));
  AN4        m0049(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n78_));
  NOi31      m0050(.An(h), .B(m), .C(f), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  NAi32      m0052(.An(m), .Bn(k), .C(j), .Y(mai_mai_n81_));
  NOi32      m0053(.An(h), .Bn(m), .C(f), .Y(mai_mai_n82_));
  NA2        m0054(.A(mai_mai_n82_), .B(mai_mai_n78_), .Y(mai_mai_n83_));
  OA220      m0055(.A0(mai_mai_n83_), .A1(mai_mai_n81_), .B0(mai_mai_n80_), .B1(mai_mai_n77_), .Y(mai_mai_n84_));
  NA3        m0056(.A(mai_mai_n84_), .B(mai_mai_n74_), .C(mai_mai_n64_), .Y(mai_mai_n85_));
  INV        m0057(.A(n), .Y(mai_mai_n86_));
  NOi32      m0058(.An(e), .Bn(b), .C(d), .Y(mai_mai_n87_));
  NA2        m0059(.A(mai_mai_n87_), .B(mai_mai_n86_), .Y(mai_mai_n88_));
  INV        m0060(.A(j), .Y(mai_mai_n89_));
  AN3        m0061(.A(m), .B(k), .C(i), .Y(mai_mai_n90_));
  NA3        m0062(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(m), .Y(mai_mai_n91_));
  NAi32      m0063(.An(m), .Bn(f), .C(h), .Y(mai_mai_n92_));
  NAi31      m0064(.An(j), .B(m), .C(l), .Y(mai_mai_n93_));
  NA2        m0065(.A(m), .B(l), .Y(mai_mai_n94_));
  NAi31      m0066(.An(k), .B(j), .C(m), .Y(mai_mai_n95_));
  NO3        m0067(.A(mai_mai_n95_), .B(mai_mai_n94_), .C(f), .Y(mai_mai_n96_));
  AN2        m0068(.A(j), .B(m), .Y(mai_mai_n97_));
  NOi32      m0069(.An(m), .Bn(l), .C(i), .Y(mai_mai_n98_));
  NOi21      m0070(.An(m), .B(i), .Y(mai_mai_n99_));
  NOi32      m0071(.An(m), .Bn(j), .C(k), .Y(mai_mai_n100_));
  AOI220     m0072(.A0(mai_mai_n100_), .A1(mai_mai_n99_), .B0(mai_mai_n98_), .B1(mai_mai_n97_), .Y(mai_mai_n101_));
  NAi41      m0073(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n102_));
  AN2        m0074(.A(e), .B(b), .Y(mai_mai_n103_));
  NOi31      m0075(.An(c), .B(h), .C(f), .Y(mai_mai_n104_));
  NA2        m0076(.A(mai_mai_n104_), .B(mai_mai_n103_), .Y(mai_mai_n105_));
  NO3        m0077(.A(mai_mai_n105_), .B(mai_mai_n102_), .C(m), .Y(mai_mai_n106_));
  NOi21      m0078(.An(m), .B(f), .Y(mai_mai_n107_));
  NOi21      m0079(.An(i), .B(h), .Y(mai_mai_n108_));
  NA3        m0080(.A(mai_mai_n108_), .B(mai_mai_n107_), .C(mai_mai_n36_), .Y(mai_mai_n109_));
  INV        m0081(.A(a), .Y(mai_mai_n110_));
  NA2        m0082(.A(mai_mai_n103_), .B(mai_mai_n110_), .Y(mai_mai_n111_));
  INV        m0083(.A(l), .Y(mai_mai_n112_));
  NOi21      m0084(.An(m), .B(n), .Y(mai_mai_n113_));
  AN2        m0085(.A(k), .B(h), .Y(mai_mai_n114_));
  NO2        m0086(.A(mai_mai_n109_), .B(mai_mai_n88_), .Y(mai_mai_n115_));
  INV        m0087(.A(b), .Y(mai_mai_n116_));
  NA2        m0088(.A(l), .B(j), .Y(mai_mai_n117_));
  AN2        m0089(.A(k), .B(i), .Y(mai_mai_n118_));
  NA2        m0090(.A(mai_mai_n118_), .B(mai_mai_n117_), .Y(mai_mai_n119_));
  NA2        m0091(.A(m), .B(e), .Y(mai_mai_n120_));
  NOi32      m0092(.An(c), .Bn(a), .C(d), .Y(mai_mai_n121_));
  NA2        m0093(.A(mai_mai_n121_), .B(mai_mai_n113_), .Y(mai_mai_n122_));
  NO4        m0094(.A(mai_mai_n122_), .B(mai_mai_n120_), .C(mai_mai_n119_), .D(mai_mai_n116_), .Y(mai_mai_n123_));
  NO3        m0095(.A(mai_mai_n123_), .B(mai_mai_n115_), .C(mai_mai_n106_), .Y(mai_mai_n124_));
  OAI210     m0096(.A0(mai_mai_n101_), .A1(mai_mai_n88_), .B0(mai_mai_n124_), .Y(mai_mai_n125_));
  NOi31      m0097(.An(k), .B(m), .C(j), .Y(mai_mai_n126_));
  NOi31      m0098(.An(k), .B(m), .C(i), .Y(mai_mai_n127_));
  NOi32      m0099(.An(f), .Bn(b), .C(e), .Y(mai_mai_n128_));
  NAi21      m0100(.An(m), .B(h), .Y(mai_mai_n129_));
  NAi21      m0101(.An(m), .B(n), .Y(mai_mai_n130_));
  NAi21      m0102(.An(j), .B(k), .Y(mai_mai_n131_));
  NO3        m0103(.A(mai_mai_n131_), .B(mai_mai_n130_), .C(mai_mai_n129_), .Y(mai_mai_n132_));
  NAi41      m0104(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n133_));
  NAi31      m0105(.An(j), .B(k), .C(h), .Y(mai_mai_n134_));
  NO3        m0106(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n130_), .Y(mai_mai_n135_));
  AOI210     m0107(.A0(mai_mai_n132_), .A1(mai_mai_n128_), .B0(mai_mai_n135_), .Y(mai_mai_n136_));
  NO2        m0108(.A(k), .B(j), .Y(mai_mai_n137_));
  AN2        m0109(.A(k), .B(j), .Y(mai_mai_n138_));
  NAi21      m0110(.An(c), .B(b), .Y(mai_mai_n139_));
  NA2        m0111(.A(f), .B(d), .Y(mai_mai_n140_));
  NA2        m0112(.A(h), .B(c), .Y(mai_mai_n141_));
  NAi31      m0113(.An(f), .B(e), .C(b), .Y(mai_mai_n142_));
  NA2        m0114(.A(d), .B(b), .Y(mai_mai_n143_));
  NAi21      m0115(.An(e), .B(f), .Y(mai_mai_n144_));
  NO2        m0116(.A(mai_mai_n144_), .B(mai_mai_n143_), .Y(mai_mai_n145_));
  NA2        m0117(.A(b), .B(a), .Y(mai_mai_n146_));
  NAi21      m0118(.An(e), .B(m), .Y(mai_mai_n147_));
  NAi21      m0119(.An(c), .B(d), .Y(mai_mai_n148_));
  NAi31      m0120(.An(l), .B(k), .C(h), .Y(mai_mai_n149_));
  NO2        m0121(.A(mai_mai_n130_), .B(mai_mai_n149_), .Y(mai_mai_n150_));
  INV        m0122(.A(mai_mai_n136_), .Y(mai_mai_n151_));
  NAi31      m0123(.An(e), .B(f), .C(b), .Y(mai_mai_n152_));
  NOi21      m0124(.An(m), .B(d), .Y(mai_mai_n153_));
  NO2        m0125(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  NOi21      m0126(.An(h), .B(i), .Y(mai_mai_n155_));
  NOi21      m0127(.An(k), .B(m), .Y(mai_mai_n156_));
  NA3        m0128(.A(mai_mai_n156_), .B(mai_mai_n155_), .C(n), .Y(mai_mai_n157_));
  NOi21      m0129(.An(mai_mai_n154_), .B(mai_mai_n157_), .Y(mai_mai_n158_));
  NOi21      m0130(.An(h), .B(m), .Y(mai_mai_n159_));
  NO2        m0131(.A(mai_mai_n140_), .B(mai_mai_n139_), .Y(mai_mai_n160_));
  NA2        m0132(.A(mai_mai_n160_), .B(mai_mai_n159_), .Y(mai_mai_n161_));
  NAi31      m0133(.An(l), .B(j), .C(h), .Y(mai_mai_n162_));
  NOi32      m0134(.An(n), .Bn(k), .C(m), .Y(mai_mai_n163_));
  NA2        m0135(.A(l), .B(i), .Y(mai_mai_n164_));
  NA2        m0136(.A(mai_mai_n164_), .B(mai_mai_n163_), .Y(mai_mai_n165_));
  NO2        m0137(.A(mai_mai_n165_), .B(mai_mai_n161_), .Y(mai_mai_n166_));
  NAi31      m0138(.An(d), .B(f), .C(c), .Y(mai_mai_n167_));
  NAi31      m0139(.An(e), .B(f), .C(c), .Y(mai_mai_n168_));
  NA2        m0140(.A(mai_mai_n168_), .B(mai_mai_n167_), .Y(mai_mai_n169_));
  NA2        m0141(.A(j), .B(h), .Y(mai_mai_n170_));
  OR3        m0142(.A(n), .B(m), .C(k), .Y(mai_mai_n171_));
  NO2        m0143(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  NAi32      m0144(.An(m), .Bn(k), .C(n), .Y(mai_mai_n173_));
  NO2        m0145(.A(mai_mai_n173_), .B(mai_mai_n170_), .Y(mai_mai_n174_));
  AOI220     m0146(.A0(mai_mai_n174_), .A1(mai_mai_n154_), .B0(mai_mai_n172_), .B1(mai_mai_n169_), .Y(mai_mai_n175_));
  NO2        m0147(.A(n), .B(m), .Y(mai_mai_n176_));
  NA2        m0148(.A(mai_mai_n176_), .B(mai_mai_n50_), .Y(mai_mai_n177_));
  NAi21      m0149(.An(f), .B(e), .Y(mai_mai_n178_));
  NA2        m0150(.A(d), .B(c), .Y(mai_mai_n179_));
  NO2        m0151(.A(mai_mai_n179_), .B(mai_mai_n178_), .Y(mai_mai_n180_));
  NOi21      m0152(.An(mai_mai_n180_), .B(mai_mai_n177_), .Y(mai_mai_n181_));
  NAi21      m0153(.An(d), .B(c), .Y(mai_mai_n182_));
  NAi31      m0154(.An(m), .B(n), .C(b), .Y(mai_mai_n183_));
  NA2        m0155(.A(k), .B(i), .Y(mai_mai_n184_));
  NAi21      m0156(.An(h), .B(f), .Y(mai_mai_n185_));
  NO2        m0157(.A(mai_mai_n185_), .B(mai_mai_n184_), .Y(mai_mai_n186_));
  NO2        m0158(.A(mai_mai_n183_), .B(mai_mai_n148_), .Y(mai_mai_n187_));
  NA2        m0159(.A(mai_mai_n187_), .B(mai_mai_n186_), .Y(mai_mai_n188_));
  NOi32      m0160(.An(f), .Bn(c), .C(d), .Y(mai_mai_n189_));
  NOi32      m0161(.An(f), .Bn(c), .C(e), .Y(mai_mai_n190_));
  NO2        m0162(.A(mai_mai_n190_), .B(mai_mai_n189_), .Y(mai_mai_n191_));
  NO3        m0163(.A(n), .B(m), .C(j), .Y(mai_mai_n192_));
  NA2        m0164(.A(mai_mai_n192_), .B(mai_mai_n114_), .Y(mai_mai_n193_));
  AO210      m0165(.A0(mai_mai_n193_), .A1(mai_mai_n177_), .B0(mai_mai_n191_), .Y(mai_mai_n194_));
  NAi41      m0166(.An(mai_mai_n181_), .B(mai_mai_n194_), .C(mai_mai_n188_), .D(mai_mai_n175_), .Y(mai_mai_n195_));
  OR4        m0167(.A(mai_mai_n195_), .B(mai_mai_n166_), .C(mai_mai_n158_), .D(mai_mai_n151_), .Y(mai_mai_n196_));
  NO4        m0168(.A(mai_mai_n196_), .B(mai_mai_n125_), .C(mai_mai_n85_), .D(mai_mai_n55_), .Y(mai_mai_n197_));
  NA3        m0169(.A(m), .B(mai_mai_n112_), .C(j), .Y(mai_mai_n198_));
  NAi31      m0170(.An(n), .B(h), .C(m), .Y(mai_mai_n199_));
  NO2        m0171(.A(mai_mai_n199_), .B(mai_mai_n198_), .Y(mai_mai_n200_));
  NOi32      m0172(.An(m), .Bn(k), .C(l), .Y(mai_mai_n201_));
  NA3        m0173(.A(mai_mai_n201_), .B(mai_mai_n89_), .C(m), .Y(mai_mai_n202_));
  NO2        m0174(.A(mai_mai_n202_), .B(n), .Y(mai_mai_n203_));
  AN2        m0175(.A(i), .B(m), .Y(mai_mai_n204_));
  NA3        m0176(.A(mai_mai_n76_), .B(mai_mai_n204_), .C(mai_mai_n113_), .Y(mai_mai_n205_));
  INV        m0177(.A(mai_mai_n205_), .Y(mai_mai_n206_));
  NAi41      m0178(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n207_));
  INV        m0179(.A(mai_mai_n207_), .Y(mai_mai_n208_));
  INV        m0180(.A(f), .Y(mai_mai_n209_));
  INV        m0181(.A(m), .Y(mai_mai_n210_));
  NOi31      m0182(.An(i), .B(j), .C(h), .Y(mai_mai_n211_));
  NOi21      m0183(.An(l), .B(m), .Y(mai_mai_n212_));
  NA2        m0184(.A(mai_mai_n212_), .B(mai_mai_n211_), .Y(mai_mai_n213_));
  NO3        m0185(.A(mai_mai_n213_), .B(mai_mai_n210_), .C(mai_mai_n209_), .Y(mai_mai_n214_));
  NA2        m0186(.A(mai_mai_n214_), .B(mai_mai_n208_), .Y(mai_mai_n215_));
  INV        m0187(.A(mai_mai_n215_), .Y(mai_mai_n216_));
  NOi21      m0188(.An(n), .B(m), .Y(mai_mai_n217_));
  NOi32      m0189(.An(l), .Bn(i), .C(j), .Y(mai_mai_n218_));
  NA2        m0190(.A(mai_mai_n218_), .B(mai_mai_n217_), .Y(mai_mai_n219_));
  OA220      m0191(.A0(mai_mai_n219_), .A1(mai_mai_n105_), .B0(mai_mai_n81_), .B1(mai_mai_n80_), .Y(mai_mai_n220_));
  NAi21      m0192(.An(j), .B(h), .Y(mai_mai_n221_));
  XN2        m0193(.A(i), .B(h), .Y(mai_mai_n222_));
  NA2        m0194(.A(mai_mai_n222_), .B(mai_mai_n221_), .Y(mai_mai_n223_));
  NOi31      m0195(.An(k), .B(n), .C(m), .Y(mai_mai_n224_));
  NOi31      m0196(.An(mai_mai_n224_), .B(mai_mai_n179_), .C(mai_mai_n178_), .Y(mai_mai_n225_));
  NA2        m0197(.A(mai_mai_n225_), .B(mai_mai_n223_), .Y(mai_mai_n226_));
  NAi31      m0198(.An(f), .B(e), .C(c), .Y(mai_mai_n227_));
  NO4        m0199(.A(mai_mai_n227_), .B(mai_mai_n171_), .C(mai_mai_n170_), .D(mai_mai_n59_), .Y(mai_mai_n228_));
  NA4        m0200(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n229_));
  NAi32      m0201(.An(m), .Bn(i), .C(k), .Y(mai_mai_n230_));
  NO3        m0202(.A(mai_mai_n230_), .B(mai_mai_n92_), .C(mai_mai_n229_), .Y(mai_mai_n231_));
  NA2        m0203(.A(k), .B(h), .Y(mai_mai_n232_));
  NO2        m0204(.A(mai_mai_n231_), .B(mai_mai_n228_), .Y(mai_mai_n233_));
  NAi21      m0205(.An(n), .B(a), .Y(mai_mai_n234_));
  NO2        m0206(.A(mai_mai_n234_), .B(mai_mai_n143_), .Y(mai_mai_n235_));
  NAi41      m0207(.An(m), .B(m), .C(k), .D(h), .Y(mai_mai_n236_));
  NO2        m0208(.A(mai_mai_n236_), .B(e), .Y(mai_mai_n237_));
  NO3        m0209(.A(mai_mai_n144_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n238_));
  OAI210     m0210(.A0(mai_mai_n238_), .A1(mai_mai_n237_), .B0(mai_mai_n235_), .Y(mai_mai_n239_));
  AN4        m0211(.A(mai_mai_n239_), .B(mai_mai_n233_), .C(mai_mai_n226_), .D(mai_mai_n220_), .Y(mai_mai_n240_));
  OR2        m0212(.A(h), .B(m), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n241_), .B(mai_mai_n102_), .Y(mai_mai_n242_));
  NA2        m0214(.A(mai_mai_n242_), .B(mai_mai_n128_), .Y(mai_mai_n243_));
  NAi41      m0215(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n244_));
  NA2        m0216(.A(mai_mai_n156_), .B(mai_mai_n108_), .Y(mai_mai_n245_));
  NO2        m0217(.A(n), .B(a), .Y(mai_mai_n246_));
  NAi31      m0218(.An(mai_mai_n236_), .B(mai_mai_n246_), .C(mai_mai_n103_), .Y(mai_mai_n247_));
  NAi21      m0219(.An(h), .B(i), .Y(mai_mai_n248_));
  NA2        m0220(.A(mai_mai_n176_), .B(k), .Y(mai_mai_n249_));
  NO2        m0221(.A(mai_mai_n249_), .B(mai_mai_n248_), .Y(mai_mai_n250_));
  NA2        m0222(.A(mai_mai_n250_), .B(mai_mai_n189_), .Y(mai_mai_n251_));
  NA3        m0223(.A(mai_mai_n251_), .B(mai_mai_n247_), .C(mai_mai_n243_), .Y(mai_mai_n252_));
  NOi21      m0224(.An(m), .B(e), .Y(mai_mai_n253_));
  NO2        m0225(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n254_));
  NA2        m0226(.A(mai_mai_n254_), .B(mai_mai_n253_), .Y(mai_mai_n255_));
  NOi32      m0227(.An(l), .Bn(j), .C(i), .Y(mai_mai_n256_));
  AOI210     m0228(.A0(mai_mai_n76_), .A1(mai_mai_n89_), .B0(mai_mai_n256_), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n248_), .B(mai_mai_n44_), .Y(mai_mai_n258_));
  NAi21      m0230(.An(f), .B(m), .Y(mai_mai_n259_));
  NO2        m0231(.A(mai_mai_n259_), .B(mai_mai_n65_), .Y(mai_mai_n260_));
  NO2        m0232(.A(mai_mai_n69_), .B(mai_mai_n117_), .Y(mai_mai_n261_));
  AOI220     m0233(.A0(mai_mai_n261_), .A1(mai_mai_n260_), .B0(mai_mai_n258_), .B1(mai_mai_n67_), .Y(mai_mai_n262_));
  OAI210     m0234(.A0(mai_mai_n257_), .A1(mai_mai_n255_), .B0(mai_mai_n262_), .Y(mai_mai_n263_));
  NO3        m0235(.A(mai_mai_n131_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n264_));
  NOi41      m0236(.An(mai_mai_n240_), .B(mai_mai_n263_), .C(mai_mai_n252_), .D(mai_mai_n216_), .Y(mai_mai_n265_));
  NO4        m0237(.A(mai_mai_n200_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n266_));
  NO2        m0238(.A(mai_mai_n266_), .B(mai_mai_n111_), .Y(mai_mai_n267_));
  NA3        m0239(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n268_));
  NAi21      m0240(.An(h), .B(m), .Y(mai_mai_n269_));
  OR4        m0241(.A(mai_mai_n269_), .B(mai_mai_n268_), .C(mai_mai_n219_), .D(e), .Y(mai_mai_n270_));
  NO2        m0242(.A(mai_mai_n245_), .B(mai_mai_n259_), .Y(mai_mai_n271_));
  NA2        m0243(.A(mai_mai_n271_), .B(mai_mai_n78_), .Y(mai_mai_n272_));
  NAi31      m0244(.An(m), .B(k), .C(h), .Y(mai_mai_n273_));
  NO3        m0245(.A(mai_mai_n130_), .B(mai_mai_n273_), .C(l), .Y(mai_mai_n274_));
  NAi31      m0246(.An(e), .B(d), .C(a), .Y(mai_mai_n275_));
  NA2        m0247(.A(mai_mai_n274_), .B(mai_mai_n128_), .Y(mai_mai_n276_));
  NA3        m0248(.A(mai_mai_n276_), .B(mai_mai_n272_), .C(mai_mai_n270_), .Y(mai_mai_n277_));
  NA4        m0249(.A(mai_mai_n156_), .B(mai_mai_n82_), .C(mai_mai_n78_), .D(mai_mai_n117_), .Y(mai_mai_n278_));
  NA3        m0250(.A(mai_mai_n156_), .B(mai_mai_n155_), .C(mai_mai_n86_), .Y(mai_mai_n279_));
  NO2        m0251(.A(mai_mai_n279_), .B(mai_mai_n191_), .Y(mai_mai_n280_));
  NOi21      m0252(.An(mai_mai_n278_), .B(mai_mai_n280_), .Y(mai_mai_n281_));
  NA3        m0253(.A(e), .B(c), .C(b), .Y(mai_mai_n282_));
  NO2        m0254(.A(mai_mai_n60_), .B(mai_mai_n282_), .Y(mai_mai_n283_));
  NAi32      m0255(.An(k), .Bn(i), .C(j), .Y(mai_mai_n284_));
  NAi31      m0256(.An(h), .B(l), .C(i), .Y(mai_mai_n285_));
  NA3        m0257(.A(mai_mai_n285_), .B(mai_mai_n284_), .C(mai_mai_n162_), .Y(mai_mai_n286_));
  NOi21      m0258(.An(mai_mai_n286_), .B(mai_mai_n49_), .Y(mai_mai_n287_));
  OAI210     m0259(.A0(mai_mai_n260_), .A1(mai_mai_n283_), .B0(mai_mai_n287_), .Y(mai_mai_n288_));
  NAi21      m0260(.An(l), .B(k), .Y(mai_mai_n289_));
  NO2        m0261(.A(mai_mai_n289_), .B(mai_mai_n49_), .Y(mai_mai_n290_));
  NOi21      m0262(.An(l), .B(j), .Y(mai_mai_n291_));
  NA2        m0263(.A(mai_mai_n159_), .B(mai_mai_n291_), .Y(mai_mai_n292_));
  NA3        m0264(.A(mai_mai_n118_), .B(mai_mai_n117_), .C(m), .Y(mai_mai_n293_));
  OR3        m0265(.A(mai_mai_n73_), .B(mai_mai_n75_), .C(e), .Y(mai_mai_n294_));
  AOI210     m0266(.A0(mai_mai_n293_), .A1(mai_mai_n292_), .B0(mai_mai_n294_), .Y(mai_mai_n295_));
  INV        m0267(.A(mai_mai_n295_), .Y(mai_mai_n296_));
  NAi32      m0268(.An(j), .Bn(h), .C(i), .Y(mai_mai_n297_));
  NAi21      m0269(.An(m), .B(l), .Y(mai_mai_n298_));
  NO3        m0270(.A(mai_mai_n298_), .B(mai_mai_n297_), .C(mai_mai_n86_), .Y(mai_mai_n299_));
  NA2        m0271(.A(h), .B(m), .Y(mai_mai_n300_));
  NA2        m0272(.A(mai_mai_n299_), .B(mai_mai_n160_), .Y(mai_mai_n301_));
  NA4        m0273(.A(mai_mai_n301_), .B(mai_mai_n296_), .C(mai_mai_n288_), .D(mai_mai_n281_), .Y(mai_mai_n302_));
  NO2        m0274(.A(mai_mai_n142_), .B(d), .Y(mai_mai_n303_));
  NA2        m0275(.A(mai_mai_n303_), .B(mai_mai_n53_), .Y(mai_mai_n304_));
  NO2        m0276(.A(mai_mai_n105_), .B(mai_mai_n102_), .Y(mai_mai_n305_));
  NAi32      m0277(.An(n), .Bn(m), .C(l), .Y(mai_mai_n306_));
  NO2        m0278(.A(mai_mai_n306_), .B(mai_mai_n297_), .Y(mai_mai_n307_));
  NA2        m0279(.A(mai_mai_n307_), .B(mai_mai_n180_), .Y(mai_mai_n308_));
  NO2        m0280(.A(mai_mai_n122_), .B(mai_mai_n116_), .Y(mai_mai_n309_));
  NAi31      m0281(.An(k), .B(l), .C(j), .Y(mai_mai_n310_));
  OAI210     m0282(.A0(mai_mai_n289_), .A1(j), .B0(mai_mai_n310_), .Y(mai_mai_n311_));
  NOi21      m0283(.An(mai_mai_n311_), .B(mai_mai_n120_), .Y(mai_mai_n312_));
  NA2        m0284(.A(mai_mai_n312_), .B(mai_mai_n309_), .Y(mai_mai_n313_));
  NA3        m0285(.A(mai_mai_n313_), .B(mai_mai_n308_), .C(mai_mai_n304_), .Y(mai_mai_n314_));
  NO4        m0286(.A(mai_mai_n314_), .B(mai_mai_n302_), .C(mai_mai_n277_), .D(mai_mai_n267_), .Y(mai_mai_n315_));
  NA2        m0287(.A(mai_mai_n250_), .B(mai_mai_n190_), .Y(mai_mai_n316_));
  NAi21      m0288(.An(m), .B(k), .Y(mai_mai_n317_));
  NO2        m0289(.A(mai_mai_n222_), .B(mai_mai_n317_), .Y(mai_mai_n318_));
  NAi41      m0290(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n319_));
  NO2        m0291(.A(mai_mai_n319_), .B(mai_mai_n147_), .Y(mai_mai_n320_));
  NA2        m0292(.A(mai_mai_n320_), .B(mai_mai_n318_), .Y(mai_mai_n321_));
  NAi31      m0293(.An(i), .B(l), .C(h), .Y(mai_mai_n322_));
  NA2        m0294(.A(e), .B(c), .Y(mai_mai_n323_));
  NO3        m0295(.A(mai_mai_n323_), .B(n), .C(d), .Y(mai_mai_n324_));
  NOi21      m0296(.An(f), .B(h), .Y(mai_mai_n325_));
  NA2        m0297(.A(mai_mai_n325_), .B(mai_mai_n118_), .Y(mai_mai_n326_));
  NO2        m0298(.A(mai_mai_n326_), .B(mai_mai_n210_), .Y(mai_mai_n327_));
  NAi31      m0299(.An(d), .B(e), .C(b), .Y(mai_mai_n328_));
  NO2        m0300(.A(mai_mai_n130_), .B(mai_mai_n328_), .Y(mai_mai_n329_));
  NA2        m0301(.A(mai_mai_n329_), .B(mai_mai_n327_), .Y(mai_mai_n330_));
  NA3        m0302(.A(mai_mai_n330_), .B(mai_mai_n321_), .C(mai_mai_n316_), .Y(mai_mai_n331_));
  NO4        m0303(.A(mai_mai_n319_), .B(mai_mai_n81_), .C(mai_mai_n72_), .D(mai_mai_n210_), .Y(mai_mai_n332_));
  NA2        m0304(.A(mai_mai_n246_), .B(mai_mai_n103_), .Y(mai_mai_n333_));
  OR2        m0305(.A(mai_mai_n333_), .B(mai_mai_n202_), .Y(mai_mai_n334_));
  NOi31      m0306(.An(l), .B(n), .C(m), .Y(mai_mai_n335_));
  NA2        m0307(.A(mai_mai_n335_), .B(mai_mai_n211_), .Y(mai_mai_n336_));
  NO2        m0308(.A(mai_mai_n336_), .B(mai_mai_n191_), .Y(mai_mai_n337_));
  NAi32      m0309(.An(mai_mai_n337_), .Bn(mai_mai_n332_), .C(mai_mai_n334_), .Y(mai_mai_n338_));
  NAi32      m0310(.An(m), .Bn(j), .C(k), .Y(mai_mai_n339_));
  NAi41      m0311(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n340_));
  OAI210     m0312(.A0(mai_mai_n207_), .A1(mai_mai_n339_), .B0(mai_mai_n340_), .Y(mai_mai_n341_));
  NOi31      m0313(.An(j), .B(m), .C(k), .Y(mai_mai_n342_));
  NO2        m0314(.A(mai_mai_n126_), .B(mai_mai_n342_), .Y(mai_mai_n343_));
  AN3        m0315(.A(h), .B(m), .C(f), .Y(mai_mai_n344_));
  NAi31      m0316(.An(mai_mai_n343_), .B(mai_mai_n344_), .C(mai_mai_n341_), .Y(mai_mai_n345_));
  NOi32      m0317(.An(m), .Bn(j), .C(l), .Y(mai_mai_n346_));
  NO2        m0318(.A(mai_mai_n346_), .B(mai_mai_n98_), .Y(mai_mai_n347_));
  NO2        m0319(.A(mai_mai_n298_), .B(mai_mai_n297_), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n213_), .B(m), .Y(mai_mai_n349_));
  NO2        m0321(.A(mai_mai_n152_), .B(mai_mai_n86_), .Y(mai_mai_n350_));
  NA2        m0322(.A(mai_mai_n350_), .B(mai_mai_n349_), .Y(mai_mai_n351_));
  NA2        m0323(.A(mai_mai_n230_), .B(mai_mai_n81_), .Y(mai_mai_n352_));
  NA3        m0324(.A(mai_mai_n352_), .B(mai_mai_n344_), .C(mai_mai_n208_), .Y(mai_mai_n353_));
  NA3        m0325(.A(mai_mai_n353_), .B(mai_mai_n351_), .C(mai_mai_n345_), .Y(mai_mai_n354_));
  NA3        m0326(.A(h), .B(m), .C(f), .Y(mai_mai_n355_));
  NO2        m0327(.A(mai_mai_n355_), .B(mai_mai_n77_), .Y(mai_mai_n356_));
  NA2        m0328(.A(mai_mai_n340_), .B(mai_mai_n207_), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n159_), .B(e), .Y(mai_mai_n358_));
  NO2        m0330(.A(mai_mai_n358_), .B(mai_mai_n41_), .Y(mai_mai_n359_));
  AOI220     m0331(.A0(mai_mai_n359_), .A1(mai_mai_n309_), .B0(mai_mai_n357_), .B1(mai_mai_n356_), .Y(mai_mai_n360_));
  NOi32      m0332(.An(j), .Bn(m), .C(i), .Y(mai_mai_n361_));
  NA3        m0333(.A(mai_mai_n361_), .B(mai_mai_n289_), .C(mai_mai_n113_), .Y(mai_mai_n362_));
  AO210      m0334(.A0(mai_mai_n111_), .A1(mai_mai_n32_), .B0(mai_mai_n362_), .Y(mai_mai_n363_));
  NOi32      m0335(.An(e), .Bn(b), .C(a), .Y(mai_mai_n364_));
  AN2        m0336(.A(l), .B(j), .Y(mai_mai_n365_));
  NO2        m0337(.A(mai_mai_n317_), .B(mai_mai_n365_), .Y(mai_mai_n366_));
  NO3        m0338(.A(mai_mai_n319_), .B(mai_mai_n72_), .C(mai_mai_n210_), .Y(mai_mai_n367_));
  NA2        m0339(.A(mai_mai_n205_), .B(mai_mai_n35_), .Y(mai_mai_n368_));
  AOI220     m0340(.A0(mai_mai_n368_), .A1(mai_mai_n364_), .B0(mai_mai_n367_), .B1(mai_mai_n366_), .Y(mai_mai_n369_));
  NO2        m0341(.A(mai_mai_n328_), .B(n), .Y(mai_mai_n370_));
  NA2        m0342(.A(mai_mai_n204_), .B(k), .Y(mai_mai_n371_));
  NA3        m0343(.A(m), .B(mai_mai_n112_), .C(mai_mai_n209_), .Y(mai_mai_n372_));
  NA4        m0344(.A(mai_mai_n201_), .B(mai_mai_n89_), .C(m), .D(mai_mai_n209_), .Y(mai_mai_n373_));
  NO2        m0345(.A(mai_mai_n372_), .B(mai_mai_n371_), .Y(mai_mai_n374_));
  NAi41      m0346(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n375_));
  NA2        m0347(.A(mai_mai_n51_), .B(mai_mai_n113_), .Y(mai_mai_n376_));
  NO2        m0348(.A(mai_mai_n376_), .B(mai_mai_n375_), .Y(mai_mai_n377_));
  AOI220     m0349(.A0(mai_mai_n377_), .A1(b), .B0(mai_mai_n374_), .B1(mai_mai_n370_), .Y(mai_mai_n378_));
  NA4        m0350(.A(mai_mai_n378_), .B(mai_mai_n369_), .C(mai_mai_n363_), .D(mai_mai_n360_), .Y(mai_mai_n379_));
  NO4        m0351(.A(mai_mai_n379_), .B(mai_mai_n354_), .C(mai_mai_n338_), .D(mai_mai_n331_), .Y(mai_mai_n380_));
  NA4        m0352(.A(mai_mai_n380_), .B(mai_mai_n315_), .C(mai_mai_n265_), .D(mai_mai_n197_), .Y(mai10));
  NA3        m0353(.A(m), .B(k), .C(i), .Y(mai_mai_n382_));
  NO3        m0354(.A(mai_mai_n382_), .B(j), .C(mai_mai_n210_), .Y(mai_mai_n383_));
  NOi21      m0355(.An(e), .B(f), .Y(mai_mai_n384_));
  NO4        m0356(.A(mai_mai_n148_), .B(mai_mai_n384_), .C(n), .D(mai_mai_n110_), .Y(mai_mai_n385_));
  NAi31      m0357(.An(b), .B(f), .C(c), .Y(mai_mai_n386_));
  INV        m0358(.A(mai_mai_n386_), .Y(mai_mai_n387_));
  NOi32      m0359(.An(k), .Bn(h), .C(j), .Y(mai_mai_n388_));
  NA2        m0360(.A(mai_mai_n388_), .B(mai_mai_n217_), .Y(mai_mai_n389_));
  NA2        m0361(.A(mai_mai_n157_), .B(mai_mai_n389_), .Y(mai_mai_n390_));
  AOI220     m0362(.A0(mai_mai_n390_), .A1(mai_mai_n387_), .B0(mai_mai_n385_), .B1(mai_mai_n383_), .Y(mai_mai_n391_));
  AN2        m0363(.A(j), .B(h), .Y(mai_mai_n392_));
  NO3        m0364(.A(n), .B(m), .C(k), .Y(mai_mai_n393_));
  NA2        m0365(.A(mai_mai_n393_), .B(mai_mai_n392_), .Y(mai_mai_n394_));
  NO3        m0366(.A(mai_mai_n394_), .B(mai_mai_n148_), .C(mai_mai_n209_), .Y(mai_mai_n395_));
  OR2        m0367(.A(m), .B(k), .Y(mai_mai_n396_));
  NO2        m0368(.A(mai_mai_n170_), .B(mai_mai_n396_), .Y(mai_mai_n397_));
  NA4        m0369(.A(n), .B(f), .C(c), .D(mai_mai_n116_), .Y(mai_mai_n398_));
  NOi21      m0370(.An(mai_mai_n397_), .B(mai_mai_n398_), .Y(mai_mai_n399_));
  NOi32      m0371(.An(d), .Bn(a), .C(c), .Y(mai_mai_n400_));
  NA2        m0372(.A(mai_mai_n400_), .B(mai_mai_n178_), .Y(mai_mai_n401_));
  NAi21      m0373(.An(i), .B(m), .Y(mai_mai_n402_));
  NAi31      m0374(.An(k), .B(m), .C(j), .Y(mai_mai_n403_));
  NO2        m0375(.A(mai_mai_n399_), .B(mai_mai_n395_), .Y(mai_mai_n404_));
  NO2        m0376(.A(mai_mai_n398_), .B(mai_mai_n298_), .Y(mai_mai_n405_));
  NOi32      m0377(.An(f), .Bn(d), .C(c), .Y(mai_mai_n406_));
  AOI220     m0378(.A0(mai_mai_n406_), .A1(mai_mai_n307_), .B0(mai_mai_n405_), .B1(mai_mai_n211_), .Y(mai_mai_n407_));
  NA3        m0379(.A(mai_mai_n407_), .B(mai_mai_n404_), .C(mai_mai_n391_), .Y(mai_mai_n408_));
  NO2        m0380(.A(mai_mai_n59_), .B(mai_mai_n116_), .Y(mai_mai_n409_));
  NA2        m0381(.A(mai_mai_n246_), .B(mai_mai_n409_), .Y(mai_mai_n410_));
  INV        m0382(.A(e), .Y(mai_mai_n411_));
  NA2        m0383(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n412_));
  OAI220     m0384(.A0(mai_mai_n412_), .A1(mai_mai_n198_), .B0(mai_mai_n202_), .B1(mai_mai_n411_), .Y(mai_mai_n413_));
  AN2        m0385(.A(m), .B(e), .Y(mai_mai_n414_));
  NA3        m0386(.A(mai_mai_n414_), .B(mai_mai_n201_), .C(i), .Y(mai_mai_n415_));
  NO2        m0387(.A(mai_mai_n101_), .B(mai_mai_n411_), .Y(mai_mai_n416_));
  NO2        m0388(.A(mai_mai_n416_), .B(mai_mai_n413_), .Y(mai_mai_n417_));
  NOi32      m0389(.An(h), .Bn(e), .C(m), .Y(mai_mai_n418_));
  NA3        m0390(.A(mai_mai_n418_), .B(mai_mai_n291_), .C(m), .Y(mai_mai_n419_));
  NOi21      m0391(.An(m), .B(h), .Y(mai_mai_n420_));
  AN3        m0392(.A(m), .B(l), .C(i), .Y(mai_mai_n421_));
  NA3        m0393(.A(mai_mai_n421_), .B(mai_mai_n420_), .C(e), .Y(mai_mai_n422_));
  AN3        m0394(.A(h), .B(m), .C(e), .Y(mai_mai_n423_));
  NA2        m0395(.A(mai_mai_n423_), .B(mai_mai_n98_), .Y(mai_mai_n424_));
  AN3        m0396(.A(mai_mai_n424_), .B(mai_mai_n422_), .C(mai_mai_n419_), .Y(mai_mai_n425_));
  AOI210     m0397(.A0(mai_mai_n425_), .A1(mai_mai_n417_), .B0(mai_mai_n410_), .Y(mai_mai_n426_));
  NA3        m0398(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n427_));
  NO2        m0399(.A(mai_mai_n427_), .B(mai_mai_n410_), .Y(mai_mai_n428_));
  NA3        m0400(.A(mai_mai_n400_), .B(mai_mai_n178_), .C(mai_mai_n86_), .Y(mai_mai_n429_));
  NAi31      m0401(.An(b), .B(c), .C(a), .Y(mai_mai_n430_));
  NO2        m0402(.A(mai_mai_n430_), .B(n), .Y(mai_mai_n431_));
  OAI210     m0403(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n432_));
  NO2        m0404(.A(mai_mai_n432_), .B(mai_mai_n144_), .Y(mai_mai_n433_));
  NA2        m0405(.A(mai_mai_n433_), .B(mai_mai_n431_), .Y(mai_mai_n434_));
  INV        m0406(.A(mai_mai_n434_), .Y(mai_mai_n435_));
  NO4        m0407(.A(mai_mai_n435_), .B(mai_mai_n428_), .C(mai_mai_n426_), .D(mai_mai_n408_), .Y(mai_mai_n436_));
  NA2        m0408(.A(i), .B(m), .Y(mai_mai_n437_));
  NO3        m0409(.A(mai_mai_n275_), .B(mai_mai_n437_), .C(c), .Y(mai_mai_n438_));
  NOi21      m0410(.An(a), .B(n), .Y(mai_mai_n439_));
  NOi21      m0411(.An(d), .B(c), .Y(mai_mai_n440_));
  NA2        m0412(.A(mai_mai_n440_), .B(mai_mai_n439_), .Y(mai_mai_n441_));
  NA3        m0413(.A(i), .B(m), .C(f), .Y(mai_mai_n442_));
  OR2        m0414(.A(mai_mai_n442_), .B(mai_mai_n71_), .Y(mai_mai_n443_));
  NA3        m0415(.A(mai_mai_n421_), .B(mai_mai_n420_), .C(mai_mai_n178_), .Y(mai_mai_n444_));
  AOI210     m0416(.A0(mai_mai_n444_), .A1(mai_mai_n443_), .B0(mai_mai_n441_), .Y(mai_mai_n445_));
  AOI210     m0417(.A0(mai_mai_n438_), .A1(mai_mai_n290_), .B0(mai_mai_n445_), .Y(mai_mai_n446_));
  OR2        m0418(.A(n), .B(m), .Y(mai_mai_n447_));
  NO2        m0419(.A(mai_mai_n447_), .B(mai_mai_n149_), .Y(mai_mai_n448_));
  NO2        m0420(.A(mai_mai_n179_), .B(mai_mai_n144_), .Y(mai_mai_n449_));
  OAI210     m0421(.A0(mai_mai_n448_), .A1(mai_mai_n172_), .B0(mai_mai_n449_), .Y(mai_mai_n450_));
  INV        m0422(.A(mai_mai_n376_), .Y(mai_mai_n451_));
  NA3        m0423(.A(mai_mai_n451_), .B(mai_mai_n364_), .C(d), .Y(mai_mai_n452_));
  NO2        m0424(.A(mai_mai_n430_), .B(mai_mai_n49_), .Y(mai_mai_n453_));
  NAi21      m0425(.An(k), .B(j), .Y(mai_mai_n454_));
  NAi21      m0426(.An(e), .B(d), .Y(mai_mai_n455_));
  NO2        m0427(.A(mai_mai_n455_), .B(mai_mai_n56_), .Y(mai_mai_n456_));
  NO2        m0428(.A(mai_mai_n249_), .B(mai_mai_n209_), .Y(mai_mai_n457_));
  NA3        m0429(.A(mai_mai_n457_), .B(mai_mai_n456_), .C(mai_mai_n223_), .Y(mai_mai_n458_));
  NA3        m0430(.A(mai_mai_n458_), .B(mai_mai_n452_), .C(mai_mai_n450_), .Y(mai_mai_n459_));
  NO2        m0431(.A(mai_mai_n336_), .B(mai_mai_n209_), .Y(mai_mai_n460_));
  NA2        m0432(.A(mai_mai_n460_), .B(mai_mai_n456_), .Y(mai_mai_n461_));
  NOi31      m0433(.An(n), .B(m), .C(k), .Y(mai_mai_n462_));
  AOI220     m0434(.A0(mai_mai_n462_), .A1(mai_mai_n392_), .B0(mai_mai_n217_), .B1(mai_mai_n50_), .Y(mai_mai_n463_));
  NAi31      m0435(.An(m), .B(f), .C(c), .Y(mai_mai_n464_));
  OR3        m0436(.A(mai_mai_n464_), .B(mai_mai_n463_), .C(e), .Y(mai_mai_n465_));
  NA3        m0437(.A(mai_mai_n465_), .B(mai_mai_n461_), .C(mai_mai_n308_), .Y(mai_mai_n466_));
  NOi41      m0438(.An(mai_mai_n446_), .B(mai_mai_n466_), .C(mai_mai_n459_), .D(mai_mai_n263_), .Y(mai_mai_n467_));
  NOi32      m0439(.An(c), .Bn(a), .C(b), .Y(mai_mai_n468_));
  NA2        m0440(.A(mai_mai_n468_), .B(mai_mai_n113_), .Y(mai_mai_n469_));
  NA2        m0441(.A(mai_mai_n273_), .B(mai_mai_n149_), .Y(mai_mai_n470_));
  AN2        m0442(.A(e), .B(d), .Y(mai_mai_n471_));
  NA2        m0443(.A(mai_mai_n471_), .B(mai_mai_n470_), .Y(mai_mai_n472_));
  INV        m0444(.A(mai_mai_n144_), .Y(mai_mai_n473_));
  NO2        m0445(.A(mai_mai_n129_), .B(mai_mai_n41_), .Y(mai_mai_n474_));
  NO2        m0446(.A(mai_mai_n66_), .B(e), .Y(mai_mai_n475_));
  NOi31      m0447(.An(j), .B(k), .C(i), .Y(mai_mai_n476_));
  NOi21      m0448(.An(mai_mai_n162_), .B(mai_mai_n476_), .Y(mai_mai_n477_));
  NA4        m0449(.A(mai_mai_n322_), .B(mai_mai_n477_), .C(mai_mai_n257_), .D(mai_mai_n119_), .Y(mai_mai_n478_));
  AOI220     m0450(.A0(mai_mai_n478_), .A1(mai_mai_n475_), .B0(mai_mai_n474_), .B1(mai_mai_n473_), .Y(mai_mai_n479_));
  AOI210     m0451(.A0(mai_mai_n479_), .A1(mai_mai_n472_), .B0(mai_mai_n469_), .Y(mai_mai_n480_));
  NO2        m0452(.A(mai_mai_n206_), .B(mai_mai_n203_), .Y(mai_mai_n481_));
  NOi21      m0453(.An(a), .B(b), .Y(mai_mai_n482_));
  NA3        m0454(.A(e), .B(d), .C(c), .Y(mai_mai_n483_));
  NAi21      m0455(.An(mai_mai_n483_), .B(mai_mai_n482_), .Y(mai_mai_n484_));
  NO2        m0456(.A(mai_mai_n429_), .B(mai_mai_n202_), .Y(mai_mai_n485_));
  NOi21      m0457(.An(mai_mai_n484_), .B(mai_mai_n485_), .Y(mai_mai_n486_));
  AOI210     m0458(.A0(mai_mai_n266_), .A1(mai_mai_n481_), .B0(mai_mai_n486_), .Y(mai_mai_n487_));
  NO4        m0459(.A(mai_mai_n185_), .B(mai_mai_n102_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n488_));
  NA2        m0460(.A(mai_mai_n387_), .B(mai_mai_n150_), .Y(mai_mai_n489_));
  OR2        m0461(.A(k), .B(j), .Y(mai_mai_n490_));
  NA2        m0462(.A(l), .B(k), .Y(mai_mai_n491_));
  NA3        m0463(.A(mai_mai_n491_), .B(mai_mai_n490_), .C(mai_mai_n217_), .Y(mai_mai_n492_));
  AOI210     m0464(.A0(mai_mai_n230_), .A1(mai_mai_n339_), .B0(mai_mai_n86_), .Y(mai_mai_n493_));
  NOi21      m0465(.An(mai_mai_n492_), .B(mai_mai_n493_), .Y(mai_mai_n494_));
  OR3        m0466(.A(mai_mai_n494_), .B(mai_mai_n141_), .C(mai_mai_n133_), .Y(mai_mai_n495_));
  INV        m0467(.A(mai_mai_n278_), .Y(mai_mai_n496_));
  NA2        m0468(.A(mai_mai_n400_), .B(mai_mai_n113_), .Y(mai_mai_n497_));
  NO4        m0469(.A(mai_mai_n497_), .B(mai_mai_n95_), .C(mai_mai_n112_), .D(e), .Y(mai_mai_n498_));
  NO3        m0470(.A(mai_mai_n429_), .B(mai_mai_n93_), .C(mai_mai_n129_), .Y(mai_mai_n499_));
  NO3        m0471(.A(mai_mai_n499_), .B(mai_mai_n498_), .C(mai_mai_n496_), .Y(mai_mai_n500_));
  NA3        m0472(.A(mai_mai_n500_), .B(mai_mai_n495_), .C(mai_mai_n489_), .Y(mai_mai_n501_));
  NO4        m0473(.A(mai_mai_n501_), .B(mai_mai_n488_), .C(mai_mai_n487_), .D(mai_mai_n480_), .Y(mai_mai_n502_));
  NA2        m0474(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n503_));
  NOi21      m0475(.An(d), .B(e), .Y(mai_mai_n504_));
  NAi31      m0476(.An(j), .B(l), .C(i), .Y(mai_mai_n505_));
  OAI210     m0477(.A0(mai_mai_n505_), .A1(mai_mai_n130_), .B0(mai_mai_n102_), .Y(mai_mai_n506_));
  NO3        m0478(.A(mai_mai_n401_), .B(mai_mai_n347_), .C(mai_mai_n199_), .Y(mai_mai_n507_));
  NO2        m0479(.A(mai_mai_n401_), .B(mai_mai_n376_), .Y(mai_mai_n508_));
  NO4        m0480(.A(mai_mai_n508_), .B(mai_mai_n507_), .C(mai_mai_n181_), .D(mai_mai_n305_), .Y(mai_mai_n509_));
  NA3        m0481(.A(mai_mai_n509_), .B(mai_mai_n503_), .C(mai_mai_n240_), .Y(mai_mai_n510_));
  OAI210     m0482(.A0(mai_mai_n127_), .A1(mai_mai_n126_), .B0(n), .Y(mai_mai_n511_));
  NO2        m0483(.A(mai_mai_n511_), .B(mai_mai_n129_), .Y(mai_mai_n512_));
  AO210      m0484(.A0(mai_mai_n299_), .A1(mai_mai_n210_), .B0(mai_mai_n242_), .Y(mai_mai_n513_));
  OA210      m0485(.A0(mai_mai_n513_), .A1(mai_mai_n512_), .B0(mai_mai_n190_), .Y(mai_mai_n514_));
  XO2        m0486(.A(i), .B(h), .Y(mai_mai_n515_));
  NA3        m0487(.A(mai_mai_n515_), .B(mai_mai_n156_), .C(n), .Y(mai_mai_n516_));
  NAi41      m0488(.An(mai_mai_n299_), .B(mai_mai_n516_), .C(mai_mai_n463_), .D(mai_mai_n389_), .Y(mai_mai_n517_));
  NOi32      m0489(.An(mai_mai_n517_), .Bn(mai_mai_n475_), .C(mai_mai_n268_), .Y(mai_mai_n518_));
  NAi31      m0490(.An(c), .B(f), .C(d), .Y(mai_mai_n519_));
  AOI210     m0491(.A0(mai_mai_n279_), .A1(mai_mai_n193_), .B0(mai_mai_n519_), .Y(mai_mai_n520_));
  NOi21      m0492(.An(mai_mai_n84_), .B(mai_mai_n520_), .Y(mai_mai_n521_));
  NA3        m0493(.A(mai_mai_n385_), .B(mai_mai_n98_), .C(mai_mai_n97_), .Y(mai_mai_n522_));
  NA2        m0494(.A(mai_mai_n224_), .B(mai_mai_n108_), .Y(mai_mai_n523_));
  AOI210     m0495(.A0(mai_mai_n523_), .A1(mai_mai_n177_), .B0(mai_mai_n519_), .Y(mai_mai_n524_));
  AOI210     m0496(.A0(mai_mai_n362_), .A1(mai_mai_n35_), .B0(mai_mai_n484_), .Y(mai_mai_n525_));
  NOi31      m0497(.An(mai_mai_n522_), .B(mai_mai_n525_), .C(mai_mai_n524_), .Y(mai_mai_n526_));
  AN2        m0498(.A(mai_mai_n287_), .B(mai_mai_n260_), .Y(mai_mai_n527_));
  NA3        m0499(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n528_));
  NO2        m0500(.A(mai_mai_n528_), .B(mai_mai_n441_), .Y(mai_mai_n529_));
  NO2        m0501(.A(mai_mai_n529_), .B(mai_mai_n295_), .Y(mai_mai_n530_));
  NAi41      m0502(.An(mai_mai_n527_), .B(mai_mai_n530_), .C(mai_mai_n526_), .D(mai_mai_n521_), .Y(mai_mai_n531_));
  NO4        m0503(.A(mai_mai_n531_), .B(mai_mai_n518_), .C(mai_mai_n514_), .D(mai_mai_n510_), .Y(mai_mai_n532_));
  NA4        m0504(.A(mai_mai_n532_), .B(mai_mai_n502_), .C(mai_mai_n467_), .D(mai_mai_n436_), .Y(mai11));
  NO2        m0505(.A(mai_mai_n73_), .B(f), .Y(mai_mai_n534_));
  NA2        m0506(.A(j), .B(m), .Y(mai_mai_n535_));
  NAi31      m0507(.An(i), .B(m), .C(l), .Y(mai_mai_n536_));
  NA3        m0508(.A(m), .B(k), .C(j), .Y(mai_mai_n537_));
  OAI220     m0509(.A0(mai_mai_n537_), .A1(mai_mai_n129_), .B0(mai_mai_n536_), .B1(mai_mai_n535_), .Y(mai_mai_n538_));
  NA2        m0510(.A(mai_mai_n538_), .B(mai_mai_n534_), .Y(mai_mai_n539_));
  NOi32      m0511(.An(e), .Bn(b), .C(f), .Y(mai_mai_n540_));
  NA2        m0512(.A(mai_mai_n256_), .B(mai_mai_n113_), .Y(mai_mai_n541_));
  NA2        m0513(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n542_));
  NAi31      m0514(.An(d), .B(e), .C(a), .Y(mai_mai_n543_));
  NO2        m0515(.A(mai_mai_n543_), .B(n), .Y(mai_mai_n544_));
  NAi41      m0516(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n545_));
  AN2        m0517(.A(mai_mai_n545_), .B(mai_mai_n375_), .Y(mai_mai_n546_));
  AOI210     m0518(.A0(mai_mai_n546_), .A1(mai_mai_n401_), .B0(mai_mai_n269_), .Y(mai_mai_n547_));
  NA2        m0519(.A(j), .B(i), .Y(mai_mai_n548_));
  NAi31      m0520(.An(n), .B(m), .C(k), .Y(mai_mai_n549_));
  NO3        m0521(.A(mai_mai_n549_), .B(mai_mai_n548_), .C(mai_mai_n112_), .Y(mai_mai_n550_));
  NO4        m0522(.A(n), .B(d), .C(mai_mai_n116_), .D(a), .Y(mai_mai_n551_));
  OR2        m0523(.A(n), .B(c), .Y(mai_mai_n552_));
  NO2        m0524(.A(mai_mai_n552_), .B(mai_mai_n146_), .Y(mai_mai_n553_));
  NO2        m0525(.A(mai_mai_n553_), .B(mai_mai_n551_), .Y(mai_mai_n554_));
  NOi32      m0526(.An(m), .Bn(f), .C(i), .Y(mai_mai_n555_));
  AOI220     m0527(.A0(mai_mai_n555_), .A1(mai_mai_n100_), .B0(mai_mai_n538_), .B1(f), .Y(mai_mai_n556_));
  NO2        m0528(.A(mai_mai_n273_), .B(mai_mai_n49_), .Y(mai_mai_n557_));
  NO2        m0529(.A(mai_mai_n556_), .B(mai_mai_n554_), .Y(mai_mai_n558_));
  AOI210     m0530(.A0(mai_mai_n550_), .A1(mai_mai_n547_), .B0(mai_mai_n558_), .Y(mai_mai_n559_));
  NA2        m0531(.A(mai_mai_n138_), .B(mai_mai_n34_), .Y(mai_mai_n560_));
  OAI220     m0532(.A0(mai_mai_n560_), .A1(m), .B0(mai_mai_n542_), .B1(mai_mai_n230_), .Y(mai_mai_n561_));
  NOi41      m0533(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n562_));
  NAi32      m0534(.An(e), .Bn(b), .C(c), .Y(mai_mai_n563_));
  OR2        m0535(.A(mai_mai_n563_), .B(mai_mai_n86_), .Y(mai_mai_n564_));
  AN2        m0536(.A(mai_mai_n340_), .B(mai_mai_n319_), .Y(mai_mai_n565_));
  NA2        m0537(.A(mai_mai_n565_), .B(mai_mai_n564_), .Y(mai_mai_n566_));
  OA210      m0538(.A0(mai_mai_n566_), .A1(mai_mai_n562_), .B0(mai_mai_n561_), .Y(mai_mai_n567_));
  OAI220     m0539(.A0(mai_mai_n403_), .A1(mai_mai_n402_), .B0(mai_mai_n536_), .B1(mai_mai_n535_), .Y(mai_mai_n568_));
  NAi31      m0540(.An(d), .B(c), .C(a), .Y(mai_mai_n569_));
  NO2        m0541(.A(mai_mai_n569_), .B(n), .Y(mai_mai_n570_));
  NA3        m0542(.A(mai_mai_n570_), .B(mai_mai_n568_), .C(e), .Y(mai_mai_n571_));
  NO3        m0543(.A(mai_mai_n62_), .B(mai_mai_n49_), .C(mai_mai_n210_), .Y(mai_mai_n572_));
  NO2        m0544(.A(mai_mai_n227_), .B(mai_mai_n110_), .Y(mai_mai_n573_));
  NA2        m0545(.A(mai_mai_n572_), .B(mai_mai_n573_), .Y(mai_mai_n574_));
  NA2        m0546(.A(mai_mai_n574_), .B(mai_mai_n571_), .Y(mai_mai_n575_));
  NO2        m0547(.A(mai_mai_n275_), .B(n), .Y(mai_mai_n576_));
  NO2        m0548(.A(mai_mai_n431_), .B(mai_mai_n576_), .Y(mai_mai_n577_));
  NA2        m0549(.A(mai_mai_n568_), .B(f), .Y(mai_mai_n578_));
  NAi32      m0550(.An(d), .Bn(a), .C(b), .Y(mai_mai_n579_));
  NO2        m0551(.A(mai_mai_n579_), .B(mai_mai_n49_), .Y(mai_mai_n580_));
  NA2        m0552(.A(h), .B(f), .Y(mai_mai_n581_));
  NO2        m0553(.A(mai_mai_n581_), .B(mai_mai_n95_), .Y(mai_mai_n582_));
  NO3        m0554(.A(mai_mai_n173_), .B(mai_mai_n170_), .C(m), .Y(mai_mai_n583_));
  AOI220     m0555(.A0(mai_mai_n583_), .A1(mai_mai_n58_), .B0(mai_mai_n582_), .B1(mai_mai_n580_), .Y(mai_mai_n584_));
  OAI210     m0556(.A0(mai_mai_n578_), .A1(mai_mai_n577_), .B0(mai_mai_n584_), .Y(mai_mai_n585_));
  AN3        m0557(.A(j), .B(h), .C(m), .Y(mai_mai_n586_));
  NO2        m0558(.A(mai_mai_n143_), .B(c), .Y(mai_mai_n587_));
  NA3        m0559(.A(mai_mai_n587_), .B(mai_mai_n586_), .C(mai_mai_n462_), .Y(mai_mai_n588_));
  NA3        m0560(.A(f), .B(d), .C(b), .Y(mai_mai_n589_));
  NO4        m0561(.A(mai_mai_n589_), .B(mai_mai_n173_), .C(mai_mai_n170_), .D(m), .Y(mai_mai_n590_));
  INV        m0562(.A(mai_mai_n588_), .Y(mai_mai_n591_));
  NO4        m0563(.A(mai_mai_n591_), .B(mai_mai_n585_), .C(mai_mai_n575_), .D(mai_mai_n567_), .Y(mai_mai_n592_));
  AN3        m0564(.A(mai_mai_n592_), .B(mai_mai_n559_), .C(mai_mai_n539_), .Y(mai_mai_n593_));
  INV        m0565(.A(k), .Y(mai_mai_n594_));
  NA3        m0566(.A(l), .B(mai_mai_n594_), .C(i), .Y(mai_mai_n595_));
  INV        m0567(.A(mai_mai_n595_), .Y(mai_mai_n596_));
  NA4        m0568(.A(mai_mai_n400_), .B(mai_mai_n420_), .C(mai_mai_n178_), .D(mai_mai_n113_), .Y(mai_mai_n597_));
  NAi32      m0569(.An(h), .Bn(f), .C(m), .Y(mai_mai_n598_));
  NAi41      m0570(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n599_));
  OAI210     m0571(.A0(mai_mai_n543_), .A1(n), .B0(mai_mai_n599_), .Y(mai_mai_n600_));
  NA2        m0572(.A(mai_mai_n600_), .B(m), .Y(mai_mai_n601_));
  NAi31      m0573(.An(h), .B(m), .C(f), .Y(mai_mai_n602_));
  OR3        m0574(.A(mai_mai_n602_), .B(mai_mai_n275_), .C(mai_mai_n49_), .Y(mai_mai_n603_));
  NA4        m0575(.A(mai_mai_n420_), .B(mai_mai_n121_), .C(mai_mai_n113_), .D(e), .Y(mai_mai_n604_));
  AN2        m0576(.A(mai_mai_n604_), .B(mai_mai_n603_), .Y(mai_mai_n605_));
  OA210      m0577(.A0(mai_mai_n601_), .A1(mai_mai_n598_), .B0(mai_mai_n605_), .Y(mai_mai_n606_));
  NO3        m0578(.A(mai_mai_n598_), .B(mai_mai_n73_), .C(mai_mai_n75_), .Y(mai_mai_n607_));
  NO4        m0579(.A(mai_mai_n602_), .B(mai_mai_n552_), .C(mai_mai_n146_), .D(mai_mai_n75_), .Y(mai_mai_n608_));
  OR2        m0580(.A(mai_mai_n608_), .B(mai_mai_n607_), .Y(mai_mai_n609_));
  NAi31      m0581(.An(mai_mai_n609_), .B(mai_mai_n606_), .C(mai_mai_n597_), .Y(mai_mai_n610_));
  NAi31      m0582(.An(f), .B(h), .C(m), .Y(mai_mai_n611_));
  NO4        m0583(.A(mai_mai_n310_), .B(mai_mai_n611_), .C(mai_mai_n73_), .D(mai_mai_n75_), .Y(mai_mai_n612_));
  NOi32      m0584(.An(b), .Bn(a), .C(c), .Y(mai_mai_n613_));
  NOi41      m0585(.An(mai_mai_n613_), .B(mai_mai_n355_), .C(mai_mai_n69_), .D(mai_mai_n117_), .Y(mai_mai_n614_));
  OR2        m0586(.A(mai_mai_n614_), .B(mai_mai_n612_), .Y(mai_mai_n615_));
  NOi32      m0587(.An(d), .Bn(a), .C(e), .Y(mai_mai_n616_));
  NA2        m0588(.A(mai_mai_n616_), .B(mai_mai_n113_), .Y(mai_mai_n617_));
  NO2        m0589(.A(n), .B(c), .Y(mai_mai_n618_));
  NA3        m0590(.A(mai_mai_n618_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n619_));
  NAi32      m0591(.An(n), .Bn(f), .C(m), .Y(mai_mai_n620_));
  NA3        m0592(.A(mai_mai_n620_), .B(mai_mai_n619_), .C(mai_mai_n617_), .Y(mai_mai_n621_));
  NOi32      m0593(.An(e), .Bn(a), .C(d), .Y(mai_mai_n622_));
  AOI210     m0594(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n622_), .Y(mai_mai_n623_));
  AOI210     m0595(.A0(mai_mai_n623_), .A1(mai_mai_n209_), .B0(mai_mai_n560_), .Y(mai_mai_n624_));
  AOI210     m0596(.A0(mai_mai_n624_), .A1(mai_mai_n621_), .B0(mai_mai_n615_), .Y(mai_mai_n625_));
  INV        m0597(.A(mai_mai_n625_), .Y(mai_mai_n626_));
  AOI210     m0598(.A0(mai_mai_n610_), .A1(mai_mai_n596_), .B0(mai_mai_n626_), .Y(mai_mai_n627_));
  NO3        m0599(.A(mai_mai_n317_), .B(mai_mai_n61_), .C(n), .Y(mai_mai_n628_));
  NA3        m0600(.A(mai_mai_n519_), .B(mai_mai_n168_), .C(mai_mai_n167_), .Y(mai_mai_n629_));
  NA2        m0601(.A(mai_mai_n464_), .B(mai_mai_n227_), .Y(mai_mai_n630_));
  OR2        m0602(.A(mai_mai_n630_), .B(mai_mai_n629_), .Y(mai_mai_n631_));
  NA2        m0603(.A(mai_mai_n76_), .B(mai_mai_n113_), .Y(mai_mai_n632_));
  NO2        m0604(.A(mai_mai_n632_), .B(mai_mai_n45_), .Y(mai_mai_n633_));
  AOI220     m0605(.A0(mai_mai_n633_), .A1(mai_mai_n547_), .B0(mai_mai_n631_), .B1(mai_mai_n628_), .Y(mai_mai_n634_));
  NO2        m0606(.A(mai_mai_n634_), .B(mai_mai_n89_), .Y(mai_mai_n635_));
  NA3        m0607(.A(mai_mai_n562_), .B(mai_mai_n342_), .C(mai_mai_n46_), .Y(mai_mai_n636_));
  NOi32      m0608(.An(e), .Bn(c), .C(f), .Y(mai_mai_n637_));
  NOi21      m0609(.An(f), .B(m), .Y(mai_mai_n638_));
  NO2        m0610(.A(mai_mai_n638_), .B(mai_mai_n207_), .Y(mai_mai_n639_));
  AOI220     m0611(.A0(mai_mai_n639_), .A1(mai_mai_n397_), .B0(mai_mai_n637_), .B1(mai_mai_n172_), .Y(mai_mai_n640_));
  NA3        m0612(.A(mai_mai_n640_), .B(mai_mai_n636_), .C(mai_mai_n175_), .Y(mai_mai_n641_));
  AOI210     m0613(.A0(mai_mai_n546_), .A1(mai_mai_n401_), .B0(mai_mai_n300_), .Y(mai_mai_n642_));
  NA2        m0614(.A(mai_mai_n642_), .B(mai_mai_n261_), .Y(mai_mai_n643_));
  NOi21      m0615(.An(j), .B(l), .Y(mai_mai_n644_));
  NAi21      m0616(.An(k), .B(h), .Y(mai_mai_n645_));
  NO2        m0617(.A(mai_mai_n645_), .B(mai_mai_n259_), .Y(mai_mai_n646_));
  NOi31      m0618(.An(m), .B(n), .C(k), .Y(mai_mai_n647_));
  NA2        m0619(.A(mai_mai_n644_), .B(mai_mai_n647_), .Y(mai_mai_n648_));
  AOI210     m0620(.A0(mai_mai_n401_), .A1(mai_mai_n375_), .B0(mai_mai_n300_), .Y(mai_mai_n649_));
  NAi21      m0621(.An(mai_mai_n648_), .B(mai_mai_n649_), .Y(mai_mai_n650_));
  NO2        m0622(.A(mai_mai_n543_), .B(mai_mai_n49_), .Y(mai_mai_n651_));
  NA2        m0623(.A(mai_mai_n650_), .B(mai_mai_n643_), .Y(mai_mai_n652_));
  NA2        m0624(.A(mai_mai_n108_), .B(mai_mai_n36_), .Y(mai_mai_n653_));
  NO2        m0625(.A(k), .B(mai_mai_n210_), .Y(mai_mai_n654_));
  INV        m0626(.A(mai_mai_n364_), .Y(mai_mai_n655_));
  NO2        m0627(.A(mai_mai_n655_), .B(n), .Y(mai_mai_n656_));
  NAi31      m0628(.An(mai_mai_n653_), .B(mai_mai_n656_), .C(mai_mai_n654_), .Y(mai_mai_n657_));
  NO2        m0629(.A(mai_mai_n542_), .B(mai_mai_n173_), .Y(mai_mai_n658_));
  NA3        m0630(.A(mai_mai_n563_), .B(mai_mai_n268_), .C(mai_mai_n142_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n515_), .B(mai_mai_n156_), .Y(mai_mai_n660_));
  NO3        m0632(.A(mai_mai_n398_), .B(mai_mai_n660_), .C(mai_mai_n89_), .Y(mai_mai_n661_));
  AOI210     m0633(.A0(mai_mai_n659_), .A1(mai_mai_n658_), .B0(mai_mai_n661_), .Y(mai_mai_n662_));
  AN3        m0634(.A(f), .B(d), .C(b), .Y(mai_mai_n663_));
  OAI210     m0635(.A0(mai_mai_n663_), .A1(mai_mai_n128_), .B0(n), .Y(mai_mai_n664_));
  NA3        m0636(.A(mai_mai_n515_), .B(mai_mai_n156_), .C(mai_mai_n210_), .Y(mai_mai_n665_));
  AOI210     m0637(.A0(mai_mai_n664_), .A1(mai_mai_n229_), .B0(mai_mai_n665_), .Y(mai_mai_n666_));
  NAi31      m0638(.An(m), .B(n), .C(k), .Y(mai_mai_n667_));
  INV        m0639(.A(mai_mai_n247_), .Y(mai_mai_n668_));
  OAI210     m0640(.A0(mai_mai_n668_), .A1(mai_mai_n666_), .B0(j), .Y(mai_mai_n669_));
  NA3        m0641(.A(mai_mai_n669_), .B(mai_mai_n662_), .C(mai_mai_n657_), .Y(mai_mai_n670_));
  NO4        m0642(.A(mai_mai_n670_), .B(mai_mai_n652_), .C(mai_mai_n641_), .D(mai_mai_n635_), .Y(mai_mai_n671_));
  NA2        m0643(.A(mai_mai_n385_), .B(mai_mai_n159_), .Y(mai_mai_n672_));
  NAi31      m0644(.An(m), .B(h), .C(f), .Y(mai_mai_n673_));
  OR3        m0645(.A(mai_mai_n673_), .B(mai_mai_n275_), .C(n), .Y(mai_mai_n674_));
  OA210      m0646(.A0(mai_mai_n543_), .A1(n), .B0(mai_mai_n599_), .Y(mai_mai_n675_));
  NA3        m0647(.A(mai_mai_n418_), .B(mai_mai_n121_), .C(mai_mai_n86_), .Y(mai_mai_n676_));
  OAI210     m0648(.A0(mai_mai_n675_), .A1(mai_mai_n92_), .B0(mai_mai_n676_), .Y(mai_mai_n677_));
  NOi21      m0649(.An(mai_mai_n674_), .B(mai_mai_n677_), .Y(mai_mai_n678_));
  AOI210     m0650(.A0(mai_mai_n678_), .A1(mai_mai_n672_), .B0(mai_mai_n537_), .Y(mai_mai_n679_));
  NO3        m0651(.A(m), .B(mai_mai_n209_), .C(mai_mai_n56_), .Y(mai_mai_n680_));
  NAi21      m0652(.An(h), .B(j), .Y(mai_mai_n681_));
  NO2        m0653(.A(mai_mai_n523_), .B(mai_mai_n89_), .Y(mai_mai_n682_));
  OAI210     m0654(.A0(mai_mai_n682_), .A1(mai_mai_n397_), .B0(mai_mai_n680_), .Y(mai_mai_n683_));
  OR2        m0655(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n684_));
  NA3        m0656(.A(mai_mai_n534_), .B(mai_mai_n100_), .C(mai_mai_n99_), .Y(mai_mai_n685_));
  AN2        m0657(.A(h), .B(f), .Y(mai_mai_n686_));
  NA2        m0658(.A(mai_mai_n686_), .B(mai_mai_n37_), .Y(mai_mai_n687_));
  NA2        m0659(.A(mai_mai_n100_), .B(mai_mai_n46_), .Y(mai_mai_n688_));
  OAI220     m0660(.A0(mai_mai_n688_), .A1(mai_mai_n333_), .B0(mai_mai_n687_), .B1(mai_mai_n469_), .Y(mai_mai_n689_));
  AOI210     m0661(.A0(mai_mai_n579_), .A1(mai_mai_n430_), .B0(mai_mai_n49_), .Y(mai_mai_n690_));
  OAI220     m0662(.A0(mai_mai_n602_), .A1(mai_mai_n595_), .B0(mai_mai_n326_), .B1(mai_mai_n535_), .Y(mai_mai_n691_));
  AOI210     m0663(.A0(mai_mai_n691_), .A1(mai_mai_n690_), .B0(mai_mai_n689_), .Y(mai_mai_n692_));
  NA3        m0664(.A(mai_mai_n692_), .B(mai_mai_n685_), .C(mai_mai_n683_), .Y(mai_mai_n693_));
  NO2        m0665(.A(mai_mai_n248_), .B(f), .Y(mai_mai_n694_));
  NO2        m0666(.A(mai_mai_n638_), .B(mai_mai_n61_), .Y(mai_mai_n695_));
  NO3        m0667(.A(mai_mai_n695_), .B(mai_mai_n694_), .C(mai_mai_n34_), .Y(mai_mai_n696_));
  NA2        m0668(.A(mai_mai_n329_), .B(mai_mai_n138_), .Y(mai_mai_n697_));
  NA2        m0669(.A(mai_mai_n130_), .B(mai_mai_n49_), .Y(mai_mai_n698_));
  AOI220     m0670(.A0(mai_mai_n698_), .A1(mai_mai_n540_), .B0(mai_mai_n364_), .B1(mai_mai_n113_), .Y(mai_mai_n699_));
  OA220      m0671(.A0(mai_mai_n699_), .A1(mai_mai_n560_), .B0(mai_mai_n362_), .B1(mai_mai_n111_), .Y(mai_mai_n700_));
  OAI210     m0672(.A0(mai_mai_n697_), .A1(mai_mai_n696_), .B0(mai_mai_n700_), .Y(mai_mai_n701_));
  NO3        m0673(.A(mai_mai_n406_), .B(mai_mai_n190_), .C(mai_mai_n189_), .Y(mai_mai_n702_));
  NA2        m0674(.A(mai_mai_n702_), .B(mai_mai_n227_), .Y(mai_mai_n703_));
  NA3        m0675(.A(mai_mai_n703_), .B(mai_mai_n250_), .C(j), .Y(mai_mai_n704_));
  NO3        m0676(.A(mai_mai_n464_), .B(mai_mai_n170_), .C(i), .Y(mai_mai_n705_));
  NA2        m0677(.A(mai_mai_n468_), .B(mai_mai_n86_), .Y(mai_mai_n706_));
  NA3        m0678(.A(mai_mai_n704_), .B(mai_mai_n522_), .C(mai_mai_n404_), .Y(mai_mai_n707_));
  NO4        m0679(.A(mai_mai_n707_), .B(mai_mai_n701_), .C(mai_mai_n693_), .D(mai_mai_n679_), .Y(mai_mai_n708_));
  NA4        m0680(.A(mai_mai_n708_), .B(mai_mai_n671_), .C(mai_mai_n627_), .D(mai_mai_n593_), .Y(mai08));
  NO2        m0681(.A(k), .B(h), .Y(mai_mai_n710_));
  AO210      m0682(.A0(mai_mai_n248_), .A1(mai_mai_n454_), .B0(mai_mai_n710_), .Y(mai_mai_n711_));
  NO2        m0683(.A(mai_mai_n711_), .B(mai_mai_n298_), .Y(mai_mai_n712_));
  NA2        m0684(.A(mai_mai_n637_), .B(mai_mai_n86_), .Y(mai_mai_n713_));
  NA2        m0685(.A(mai_mai_n713_), .B(mai_mai_n464_), .Y(mai_mai_n714_));
  AOI210     m0686(.A0(mai_mai_n714_), .A1(mai_mai_n712_), .B0(mai_mai_n499_), .Y(mai_mai_n715_));
  NA2        m0687(.A(mai_mai_n86_), .B(mai_mai_n110_), .Y(mai_mai_n716_));
  NO2        m0688(.A(mai_mai_n716_), .B(mai_mai_n57_), .Y(mai_mai_n717_));
  NO4        m0689(.A(mai_mai_n382_), .B(mai_mai_n112_), .C(j), .D(mai_mai_n210_), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n589_), .B(mai_mai_n229_), .Y(mai_mai_n719_));
  AOI220     m0691(.A0(mai_mai_n719_), .A1(mai_mai_n349_), .B0(mai_mai_n718_), .B1(mai_mai_n717_), .Y(mai_mai_n720_));
  AOI210     m0692(.A0(mai_mai_n589_), .A1(mai_mai_n152_), .B0(mai_mai_n86_), .Y(mai_mai_n721_));
  NA4        m0693(.A(mai_mai_n212_), .B(mai_mai_n138_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n722_));
  AN2        m0694(.A(l), .B(k), .Y(mai_mai_n723_));
  NA4        m0695(.A(mai_mai_n723_), .B(mai_mai_n108_), .C(mai_mai_n75_), .D(mai_mai_n210_), .Y(mai_mai_n724_));
  OAI210     m0696(.A0(mai_mai_n722_), .A1(m), .B0(mai_mai_n724_), .Y(mai_mai_n725_));
  NA2        m0697(.A(mai_mai_n725_), .B(mai_mai_n721_), .Y(mai_mai_n726_));
  NA4        m0698(.A(mai_mai_n726_), .B(mai_mai_n720_), .C(mai_mai_n715_), .D(mai_mai_n351_), .Y(mai_mai_n727_));
  NO4        m0699(.A(mai_mai_n170_), .B(mai_mai_n396_), .C(mai_mai_n112_), .D(m), .Y(mai_mai_n728_));
  AOI210     m0700(.A0(mai_mai_n728_), .A1(mai_mai_n719_), .B0(mai_mai_n529_), .Y(mai_mai_n729_));
  NA2        m0701(.A(mai_mai_n639_), .B(mai_mai_n348_), .Y(mai_mai_n730_));
  NA2        m0702(.A(mai_mai_n730_), .B(mai_mai_n729_), .Y(mai_mai_n731_));
  NO2        m0703(.A(mai_mai_n546_), .B(mai_mai_n35_), .Y(mai_mai_n732_));
  INV        m0704(.A(mai_mai_n732_), .Y(mai_mai_n733_));
  NO3        m0705(.A(mai_mai_n317_), .B(mai_mai_n129_), .C(mai_mai_n41_), .Y(mai_mai_n734_));
  NA2        m0706(.A(mai_mai_n711_), .B(mai_mai_n134_), .Y(mai_mai_n735_));
  AOI220     m0707(.A0(mai_mai_n735_), .A1(mai_mai_n405_), .B0(mai_mai_n734_), .B1(mai_mai_n78_), .Y(mai_mai_n736_));
  OAI210     m0708(.A0(mai_mai_n733_), .A1(mai_mai_n89_), .B0(mai_mai_n736_), .Y(mai_mai_n737_));
  NA2        m0709(.A(mai_mai_n364_), .B(mai_mai_n43_), .Y(mai_mai_n738_));
  NA3        m0710(.A(mai_mai_n703_), .B(mai_mai_n335_), .C(mai_mai_n388_), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n723_), .B(mai_mai_n217_), .Y(mai_mai_n740_));
  NO2        m0712(.A(mai_mai_n740_), .B(mai_mai_n328_), .Y(mai_mai_n741_));
  AOI210     m0713(.A0(mai_mai_n741_), .A1(mai_mai_n694_), .B0(mai_mai_n498_), .Y(mai_mai_n742_));
  NA3        m0714(.A(m), .B(l), .C(k), .Y(mai_mai_n743_));
  AOI210     m0715(.A0(mai_mai_n676_), .A1(mai_mai_n674_), .B0(mai_mai_n743_), .Y(mai_mai_n744_));
  NO2        m0716(.A(mai_mai_n545_), .B(mai_mai_n269_), .Y(mai_mai_n745_));
  NOi21      m0717(.An(mai_mai_n745_), .B(mai_mai_n541_), .Y(mai_mai_n746_));
  NA4        m0718(.A(mai_mai_n113_), .B(l), .C(k), .D(mai_mai_n89_), .Y(mai_mai_n747_));
  NA3        m0719(.A(mai_mai_n121_), .B(mai_mai_n414_), .C(i), .Y(mai_mai_n748_));
  NO2        m0720(.A(mai_mai_n748_), .B(mai_mai_n747_), .Y(mai_mai_n749_));
  NO3        m0721(.A(mai_mai_n749_), .B(mai_mai_n746_), .C(mai_mai_n744_), .Y(mai_mai_n750_));
  NA4        m0722(.A(mai_mai_n750_), .B(mai_mai_n742_), .C(mai_mai_n739_), .D(mai_mai_n738_), .Y(mai_mai_n751_));
  NO4        m0723(.A(mai_mai_n751_), .B(mai_mai_n737_), .C(mai_mai_n731_), .D(mai_mai_n727_), .Y(mai_mai_n752_));
  NA2        m0724(.A(mai_mai_n639_), .B(mai_mai_n397_), .Y(mai_mai_n753_));
  NOi31      m0725(.An(m), .B(h), .C(f), .Y(mai_mai_n754_));
  NA2        m0726(.A(mai_mai_n651_), .B(mai_mai_n754_), .Y(mai_mai_n755_));
  AO210      m0727(.A0(mai_mai_n755_), .A1(mai_mai_n603_), .B0(mai_mai_n548_), .Y(mai_mai_n756_));
  INV        m0728(.A(mai_mai_n508_), .Y(mai_mai_n757_));
  NA4        m0729(.A(mai_mai_n757_), .B(mai_mai_n756_), .C(mai_mai_n753_), .D(mai_mai_n247_), .Y(mai_mai_n758_));
  NA2        m0730(.A(mai_mai_n723_), .B(mai_mai_n75_), .Y(mai_mai_n759_));
  NO4        m0731(.A(mai_mai_n702_), .B(mai_mai_n170_), .C(n), .D(i), .Y(mai_mai_n760_));
  NOi21      m0732(.An(h), .B(j), .Y(mai_mai_n761_));
  NA2        m0733(.A(mai_mai_n761_), .B(f), .Y(mai_mai_n762_));
  NO2        m0734(.A(mai_mai_n762_), .B(mai_mai_n244_), .Y(mai_mai_n763_));
  NO3        m0735(.A(mai_mai_n763_), .B(mai_mai_n760_), .C(mai_mai_n705_), .Y(mai_mai_n764_));
  OAI220     m0736(.A0(mai_mai_n764_), .A1(mai_mai_n759_), .B0(mai_mai_n605_), .B1(mai_mai_n62_), .Y(mai_mai_n765_));
  AOI210     m0737(.A0(mai_mai_n758_), .A1(l), .B0(mai_mai_n765_), .Y(mai_mai_n766_));
  NO2        m0738(.A(j), .B(i), .Y(mai_mai_n767_));
  NA2        m0739(.A(mai_mai_n767_), .B(mai_mai_n33_), .Y(mai_mai_n768_));
  NA2        m0740(.A(mai_mai_n423_), .B(mai_mai_n121_), .Y(mai_mai_n769_));
  OR2        m0741(.A(mai_mai_n769_), .B(mai_mai_n768_), .Y(mai_mai_n770_));
  NO3        m0742(.A(mai_mai_n148_), .B(mai_mai_n49_), .C(mai_mai_n110_), .Y(mai_mai_n771_));
  NO3        m0743(.A(mai_mai_n552_), .B(mai_mai_n146_), .C(mai_mai_n75_), .Y(mai_mai_n772_));
  NO3        m0744(.A(mai_mai_n491_), .B(mai_mai_n442_), .C(j), .Y(mai_mai_n773_));
  OAI210     m0745(.A0(mai_mai_n772_), .A1(mai_mai_n771_), .B0(mai_mai_n773_), .Y(mai_mai_n774_));
  OAI210     m0746(.A0(mai_mai_n755_), .A1(mai_mai_n62_), .B0(mai_mai_n774_), .Y(mai_mai_n775_));
  NA2        m0747(.A(k), .B(j), .Y(mai_mai_n776_));
  NO3        m0748(.A(mai_mai_n298_), .B(mai_mai_n776_), .C(mai_mai_n40_), .Y(mai_mai_n777_));
  AOI210     m0749(.A0(mai_mai_n540_), .A1(n), .B0(mai_mai_n562_), .Y(mai_mai_n778_));
  NA2        m0750(.A(mai_mai_n778_), .B(mai_mai_n565_), .Y(mai_mai_n779_));
  AN3        m0751(.A(mai_mai_n779_), .B(mai_mai_n777_), .C(mai_mai_n99_), .Y(mai_mai_n780_));
  NA2        m0752(.A(mai_mai_n630_), .B(mai_mai_n307_), .Y(mai_mai_n781_));
  INV        m0753(.A(mai_mai_n781_), .Y(mai_mai_n782_));
  NO2        m0754(.A(mai_mai_n298_), .B(mai_mai_n134_), .Y(mai_mai_n783_));
  AOI220     m0755(.A0(mai_mai_n783_), .A1(mai_mai_n639_), .B0(mai_mai_n734_), .B1(mai_mai_n721_), .Y(mai_mai_n784_));
  NO2        m0756(.A(mai_mai_n743_), .B(mai_mai_n92_), .Y(mai_mai_n785_));
  NA2        m0757(.A(mai_mai_n785_), .B(mai_mai_n600_), .Y(mai_mai_n786_));
  NO2        m0758(.A(mai_mai_n602_), .B(mai_mai_n117_), .Y(mai_mai_n787_));
  OAI210     m0759(.A0(mai_mai_n787_), .A1(mai_mai_n773_), .B0(mai_mai_n690_), .Y(mai_mai_n788_));
  NA3        m0760(.A(mai_mai_n788_), .B(mai_mai_n786_), .C(mai_mai_n784_), .Y(mai_mai_n789_));
  OR4        m0761(.A(mai_mai_n789_), .B(mai_mai_n782_), .C(mai_mai_n780_), .D(mai_mai_n775_), .Y(mai_mai_n790_));
  NA3        m0762(.A(mai_mai_n778_), .B(mai_mai_n565_), .C(mai_mai_n564_), .Y(mai_mai_n791_));
  NA4        m0763(.A(mai_mai_n791_), .B(mai_mai_n212_), .C(mai_mai_n454_), .D(mai_mai_n34_), .Y(mai_mai_n792_));
  NO4        m0764(.A(mai_mai_n491_), .B(mai_mai_n437_), .C(j), .D(f), .Y(mai_mai_n793_));
  OAI220     m0765(.A0(mai_mai_n722_), .A1(mai_mai_n713_), .B0(mai_mai_n333_), .B1(mai_mai_n38_), .Y(mai_mai_n794_));
  AOI210     m0766(.A0(mai_mai_n793_), .A1(mai_mai_n254_), .B0(mai_mai_n794_), .Y(mai_mai_n795_));
  NA3        m0767(.A(mai_mai_n555_), .B(mai_mai_n291_), .C(h), .Y(mai_mai_n796_));
  NOi21      m0768(.An(mai_mai_n690_), .B(mai_mai_n796_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n93_), .B(mai_mai_n47_), .Y(mai_mai_n798_));
  NO2        m0770(.A(mai_mai_n796_), .B(mai_mai_n619_), .Y(mai_mai_n799_));
  AOI210     m0771(.A0(mai_mai_n798_), .A1(mai_mai_n656_), .B0(mai_mai_n799_), .Y(mai_mai_n800_));
  NAi41      m0772(.An(mai_mai_n797_), .B(mai_mai_n800_), .C(mai_mai_n795_), .D(mai_mai_n792_), .Y(mai_mai_n801_));
  OR2        m0773(.A(mai_mai_n785_), .B(mai_mai_n96_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n802_), .B(mai_mai_n235_), .Y(mai_mai_n803_));
  INV        m0775(.A(mai_mai_n337_), .Y(mai_mai_n804_));
  OAI210     m0776(.A0(mai_mai_n743_), .A1(mai_mai_n673_), .B0(mai_mai_n528_), .Y(mai_mai_n805_));
  NA3        m0777(.A(mai_mai_n246_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n806_));
  AOI220     m0778(.A0(mai_mai_n618_), .A1(mai_mai_n29_), .B0(mai_mai_n468_), .B1(mai_mai_n86_), .Y(mai_mai_n807_));
  NA2        m0779(.A(mai_mai_n807_), .B(mai_mai_n806_), .Y(mai_mai_n808_));
  NO2        m0780(.A(mai_mai_n796_), .B(mai_mai_n497_), .Y(mai_mai_n809_));
  AOI210     m0781(.A0(mai_mai_n808_), .A1(mai_mai_n805_), .B0(mai_mai_n809_), .Y(mai_mai_n810_));
  NA3        m0782(.A(mai_mai_n810_), .B(mai_mai_n804_), .C(mai_mai_n803_), .Y(mai_mai_n811_));
  NOi41      m0783(.An(mai_mai_n770_), .B(mai_mai_n811_), .C(mai_mai_n801_), .D(mai_mai_n790_), .Y(mai_mai_n812_));
  OR3        m0784(.A(mai_mai_n722_), .B(mai_mai_n229_), .C(m), .Y(mai_mai_n813_));
  NO3        m0785(.A(mai_mai_n343_), .B(mai_mai_n300_), .C(mai_mai_n112_), .Y(mai_mai_n814_));
  NA2        m0786(.A(mai_mai_n814_), .B(mai_mai_n779_), .Y(mai_mai_n815_));
  NA2        m0787(.A(mai_mai_n46_), .B(mai_mai_n56_), .Y(mai_mai_n816_));
  NO3        m0788(.A(mai_mai_n816_), .B(mai_mai_n768_), .C(mai_mai_n275_), .Y(mai_mai_n817_));
  NO3        m0789(.A(mai_mai_n535_), .B(mai_mai_n94_), .C(h), .Y(mai_mai_n818_));
  AOI210     m0790(.A0(mai_mai_n818_), .A1(mai_mai_n717_), .B0(mai_mai_n817_), .Y(mai_mai_n819_));
  NA4        m0791(.A(mai_mai_n819_), .B(mai_mai_n815_), .C(mai_mai_n813_), .D(mai_mai_n407_), .Y(mai_mai_n820_));
  OR2        m0792(.A(mai_mai_n673_), .B(mai_mai_n93_), .Y(mai_mai_n821_));
  NOi31      m0793(.An(b), .B(d), .C(a), .Y(mai_mai_n822_));
  NO2        m0794(.A(mai_mai_n822_), .B(mai_mai_n616_), .Y(mai_mai_n823_));
  NO2        m0795(.A(mai_mai_n823_), .B(n), .Y(mai_mai_n824_));
  NOi21      m0796(.An(mai_mai_n807_), .B(mai_mai_n824_), .Y(mai_mai_n825_));
  NO2        m0797(.A(mai_mai_n825_), .B(mai_mai_n821_), .Y(mai_mai_n826_));
  NO2        m0798(.A(mai_mai_n563_), .B(mai_mai_n86_), .Y(mai_mai_n827_));
  NO3        m0799(.A(mai_mai_n638_), .B(mai_mai_n328_), .C(mai_mai_n117_), .Y(mai_mai_n828_));
  NOi21      m0800(.An(mai_mai_n828_), .B(mai_mai_n157_), .Y(mai_mai_n829_));
  AOI210     m0801(.A0(mai_mai_n814_), .A1(mai_mai_n827_), .B0(mai_mai_n829_), .Y(mai_mai_n830_));
  OAI210     m0802(.A0(mai_mai_n722_), .A1(mai_mai_n398_), .B0(mai_mai_n830_), .Y(mai_mai_n831_));
  NO2        m0803(.A(mai_mai_n702_), .B(n), .Y(mai_mai_n832_));
  AOI220     m0804(.A0(mai_mai_n783_), .A1(mai_mai_n680_), .B0(mai_mai_n832_), .B1(mai_mai_n712_), .Y(mai_mai_n833_));
  NO2        m0805(.A(mai_mai_n323_), .B(mai_mai_n234_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n121_), .B(mai_mai_n86_), .Y(mai_mai_n835_));
  AOI210     m0807(.A0(mai_mai_n427_), .A1(mai_mai_n419_), .B0(mai_mai_n835_), .Y(mai_mai_n836_));
  NA2        m0808(.A(mai_mai_n741_), .B(mai_mai_n34_), .Y(mai_mai_n837_));
  NAi21      m0809(.An(mai_mai_n747_), .B(mai_mai_n438_), .Y(mai_mai_n838_));
  NO2        m0810(.A(mai_mai_n269_), .B(i), .Y(mai_mai_n839_));
  NA2        m0811(.A(mai_mai_n728_), .B(mai_mai_n350_), .Y(mai_mai_n840_));
  OAI210     m0812(.A0(mai_mai_n608_), .A1(mai_mai_n607_), .B0(mai_mai_n365_), .Y(mai_mai_n841_));
  AN3        m0813(.A(mai_mai_n841_), .B(mai_mai_n840_), .C(mai_mai_n838_), .Y(mai_mai_n842_));
  NAi41      m0814(.An(mai_mai_n836_), .B(mai_mai_n842_), .C(mai_mai_n837_), .D(mai_mai_n833_), .Y(mai_mai_n843_));
  NO4        m0815(.A(mai_mai_n843_), .B(mai_mai_n831_), .C(mai_mai_n826_), .D(mai_mai_n820_), .Y(mai_mai_n844_));
  NA4        m0816(.A(mai_mai_n844_), .B(mai_mai_n812_), .C(mai_mai_n766_), .D(mai_mai_n752_), .Y(mai09));
  INV        m0817(.A(mai_mai_n122_), .Y(mai_mai_n846_));
  NA2        m0818(.A(f), .B(e), .Y(mai_mai_n847_));
  NO2        m0819(.A(mai_mai_n222_), .B(mai_mai_n112_), .Y(mai_mai_n848_));
  NA2        m0820(.A(mai_mai_n848_), .B(m), .Y(mai_mai_n849_));
  NA4        m0821(.A(mai_mai_n310_), .B(mai_mai_n477_), .C(mai_mai_n257_), .D(mai_mai_n119_), .Y(mai_mai_n850_));
  AOI210     m0822(.A0(mai_mai_n850_), .A1(m), .B0(mai_mai_n474_), .Y(mai_mai_n851_));
  AOI210     m0823(.A0(mai_mai_n851_), .A1(mai_mai_n849_), .B0(mai_mai_n847_), .Y(mai_mai_n852_));
  NA2        m0824(.A(mai_mai_n448_), .B(e), .Y(mai_mai_n853_));
  NO2        m0825(.A(mai_mai_n853_), .B(mai_mai_n519_), .Y(mai_mai_n854_));
  AOI210     m0826(.A0(mai_mai_n852_), .A1(mai_mai_n846_), .B0(mai_mai_n854_), .Y(mai_mai_n855_));
  NA3        m0827(.A(m), .B(l), .C(i), .Y(mai_mai_n856_));
  OAI220     m0828(.A0(mai_mai_n602_), .A1(mai_mai_n856_), .B0(mai_mai_n355_), .B1(mai_mai_n536_), .Y(mai_mai_n857_));
  NA4        m0829(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(m), .D(f), .Y(mai_mai_n858_));
  NAi31      m0830(.An(mai_mai_n857_), .B(mai_mai_n858_), .C(mai_mai_n443_), .Y(mai_mai_n859_));
  NA3        m0831(.A(mai_mai_n821_), .B(mai_mai_n578_), .C(mai_mai_n528_), .Y(mai_mai_n860_));
  OA210      m0832(.A0(mai_mai_n860_), .A1(mai_mai_n859_), .B0(mai_mai_n824_), .Y(mai_mai_n861_));
  INV        m0833(.A(mai_mai_n340_), .Y(mai_mai_n862_));
  NO2        m0834(.A(mai_mai_n127_), .B(mai_mai_n126_), .Y(mai_mai_n863_));
  NOi31      m0835(.An(k), .B(m), .C(l), .Y(mai_mai_n864_));
  NO2        m0836(.A(mai_mai_n342_), .B(mai_mai_n864_), .Y(mai_mai_n865_));
  AOI210     m0837(.A0(mai_mai_n865_), .A1(mai_mai_n863_), .B0(mai_mai_n611_), .Y(mai_mai_n866_));
  NA2        m0838(.A(mai_mai_n806_), .B(mai_mai_n333_), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n344_), .B(mai_mai_n346_), .Y(mai_mai_n868_));
  OAI210     m0840(.A0(mai_mai_n202_), .A1(mai_mai_n209_), .B0(mai_mai_n868_), .Y(mai_mai_n869_));
  AOI220     m0841(.A0(mai_mai_n869_), .A1(mai_mai_n867_), .B0(mai_mai_n866_), .B1(mai_mai_n862_), .Y(mai_mai_n870_));
  NA2        m0842(.A(mai_mai_n164_), .B(mai_mai_n114_), .Y(mai_mai_n871_));
  NA3        m0843(.A(mai_mai_n871_), .B(mai_mai_n711_), .C(mai_mai_n134_), .Y(mai_mai_n872_));
  NA3        m0844(.A(mai_mai_n872_), .B(mai_mai_n187_), .C(mai_mai_n31_), .Y(mai_mai_n873_));
  NA4        m0845(.A(mai_mai_n873_), .B(mai_mai_n870_), .C(mai_mai_n640_), .D(mai_mai_n84_), .Y(mai_mai_n874_));
  NO2        m0846(.A(mai_mai_n598_), .B(mai_mai_n505_), .Y(mai_mai_n875_));
  NA2        m0847(.A(mai_mai_n875_), .B(mai_mai_n187_), .Y(mai_mai_n876_));
  NOi21      m0848(.An(f), .B(d), .Y(mai_mai_n877_));
  NA2        m0849(.A(mai_mai_n877_), .B(m), .Y(mai_mai_n878_));
  NO2        m0850(.A(mai_mai_n878_), .B(mai_mai_n52_), .Y(mai_mai_n879_));
  NOi32      m0851(.An(m), .Bn(f), .C(d), .Y(mai_mai_n880_));
  NA4        m0852(.A(mai_mai_n880_), .B(mai_mai_n618_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n881_));
  NA2        m0853(.A(mai_mai_n879_), .B(mai_mai_n553_), .Y(mai_mai_n882_));
  NA3        m0854(.A(mai_mai_n310_), .B(mai_mai_n257_), .C(mai_mai_n119_), .Y(mai_mai_n883_));
  AN2        m0855(.A(f), .B(d), .Y(mai_mai_n884_));
  NA3        m0856(.A(mai_mai_n482_), .B(mai_mai_n884_), .C(mai_mai_n86_), .Y(mai_mai_n885_));
  NO3        m0857(.A(mai_mai_n885_), .B(mai_mai_n75_), .C(mai_mai_n210_), .Y(mai_mai_n886_));
  NO2        m0858(.A(mai_mai_n284_), .B(mai_mai_n56_), .Y(mai_mai_n887_));
  NA2        m0859(.A(mai_mai_n883_), .B(mai_mai_n886_), .Y(mai_mai_n888_));
  NAi41      m0860(.An(mai_mai_n496_), .B(mai_mai_n888_), .C(mai_mai_n882_), .D(mai_mai_n876_), .Y(mai_mai_n889_));
  NO4        m0861(.A(mai_mai_n638_), .B(mai_mai_n130_), .C(mai_mai_n328_), .D(mai_mai_n149_), .Y(mai_mai_n890_));
  NO2        m0862(.A(mai_mai_n667_), .B(mai_mai_n328_), .Y(mai_mai_n891_));
  AN2        m0863(.A(mai_mai_n891_), .B(mai_mai_n694_), .Y(mai_mai_n892_));
  NO3        m0864(.A(mai_mai_n892_), .B(mai_mai_n890_), .C(mai_mai_n231_), .Y(mai_mai_n893_));
  NA2        m0865(.A(mai_mai_n616_), .B(mai_mai_n86_), .Y(mai_mai_n894_));
  NA3        m0866(.A(mai_mai_n156_), .B(mai_mai_n108_), .C(mai_mai_n107_), .Y(mai_mai_n895_));
  OAI220     m0867(.A0(mai_mai_n885_), .A1(mai_mai_n432_), .B0(mai_mai_n340_), .B1(mai_mai_n895_), .Y(mai_mai_n896_));
  NOi31      m0868(.An(mai_mai_n220_), .B(mai_mai_n896_), .C(mai_mai_n305_), .Y(mai_mai_n897_));
  NA2        m0869(.A(c), .B(mai_mai_n116_), .Y(mai_mai_n898_));
  NO2        m0870(.A(mai_mai_n898_), .B(mai_mai_n411_), .Y(mai_mai_n899_));
  NA3        m0871(.A(mai_mai_n899_), .B(mai_mai_n517_), .C(f), .Y(mai_mai_n900_));
  OR2        m0872(.A(mai_mai_n673_), .B(mai_mai_n549_), .Y(mai_mai_n901_));
  INV        m0873(.A(mai_mai_n901_), .Y(mai_mai_n902_));
  NA2        m0874(.A(mai_mai_n823_), .B(mai_mai_n111_), .Y(mai_mai_n903_));
  NA2        m0875(.A(mai_mai_n903_), .B(mai_mai_n902_), .Y(mai_mai_n904_));
  NA4        m0876(.A(mai_mai_n904_), .B(mai_mai_n900_), .C(mai_mai_n897_), .D(mai_mai_n893_), .Y(mai_mai_n905_));
  NO4        m0877(.A(mai_mai_n905_), .B(mai_mai_n889_), .C(mai_mai_n874_), .D(mai_mai_n861_), .Y(mai_mai_n906_));
  OR2        m0878(.A(mai_mai_n885_), .B(mai_mai_n75_), .Y(mai_mai_n907_));
  NA2        m0879(.A(mai_mai_n112_), .B(j), .Y(mai_mai_n908_));
  NA2        m0880(.A(mai_mai_n848_), .B(m), .Y(mai_mai_n909_));
  AOI210     m0881(.A0(mai_mai_n909_), .A1(mai_mai_n292_), .B0(mai_mai_n907_), .Y(mai_mai_n910_));
  NO2        m0882(.A(mai_mai_n134_), .B(mai_mai_n130_), .Y(mai_mai_n911_));
  NO2        m0883(.A(mai_mai_n227_), .B(mai_mai_n221_), .Y(mai_mai_n912_));
  AOI220     m0884(.A0(mai_mai_n912_), .A1(mai_mai_n224_), .B0(mai_mai_n303_), .B1(mai_mai_n911_), .Y(mai_mai_n913_));
  NO2        m0885(.A(mai_mai_n432_), .B(mai_mai_n847_), .Y(mai_mai_n914_));
  NA2        m0886(.A(mai_mai_n914_), .B(mai_mai_n570_), .Y(mai_mai_n915_));
  NA2        m0887(.A(mai_mai_n915_), .B(mai_mai_n913_), .Y(mai_mai_n916_));
  NA2        m0888(.A(e), .B(d), .Y(mai_mai_n917_));
  OAI220     m0889(.A0(mai_mai_n917_), .A1(c), .B0(mai_mai_n323_), .B1(d), .Y(mai_mai_n918_));
  NA3        m0890(.A(mai_mai_n918_), .B(mai_mai_n457_), .C(mai_mai_n515_), .Y(mai_mai_n919_));
  AOI210     m0891(.A0(mai_mai_n523_), .A1(mai_mai_n177_), .B0(mai_mai_n227_), .Y(mai_mai_n920_));
  AOI210     m0892(.A0(mai_mai_n639_), .A1(mai_mai_n348_), .B0(mai_mai_n920_), .Y(mai_mai_n921_));
  NA2        m0893(.A(mai_mai_n284_), .B(mai_mai_n162_), .Y(mai_mai_n922_));
  NA2        m0894(.A(mai_mai_n886_), .B(mai_mai_n922_), .Y(mai_mai_n923_));
  NA3        m0895(.A(mai_mai_n163_), .B(mai_mai_n87_), .C(mai_mai_n34_), .Y(mai_mai_n924_));
  NA4        m0896(.A(mai_mai_n924_), .B(mai_mai_n923_), .C(mai_mai_n921_), .D(mai_mai_n919_), .Y(mai_mai_n925_));
  NO3        m0897(.A(mai_mai_n925_), .B(mai_mai_n916_), .C(mai_mai_n910_), .Y(mai_mai_n926_));
  NA2        m0898(.A(mai_mai_n862_), .B(mai_mai_n31_), .Y(mai_mai_n927_));
  AO210      m0899(.A0(mai_mai_n927_), .A1(mai_mai_n713_), .B0(mai_mai_n213_), .Y(mai_mai_n928_));
  OAI220     m0900(.A0(mai_mai_n638_), .A1(mai_mai_n61_), .B0(mai_mai_n300_), .B1(j), .Y(mai_mai_n929_));
  AOI220     m0901(.A0(mai_mai_n929_), .A1(mai_mai_n891_), .B0(mai_mai_n628_), .B1(mai_mai_n637_), .Y(mai_mai_n930_));
  OAI210     m0902(.A0(mai_mai_n853_), .A1(mai_mai_n167_), .B0(mai_mai_n930_), .Y(mai_mai_n931_));
  OAI210     m0903(.A0(mai_mai_n848_), .A1(mai_mai_n922_), .B0(mai_mai_n880_), .Y(mai_mai_n932_));
  NO2        m0904(.A(mai_mai_n932_), .B(mai_mai_n619_), .Y(mai_mai_n933_));
  AOI210     m0905(.A0(mai_mai_n118_), .A1(mai_mai_n117_), .B0(mai_mai_n256_), .Y(mai_mai_n934_));
  AN2        m0906(.A(mai_mai_n867_), .B(mai_mai_n857_), .Y(mai_mai_n935_));
  NO3        m0907(.A(mai_mai_n935_), .B(mai_mai_n933_), .C(mai_mai_n931_), .Y(mai_mai_n936_));
  AO220      m0908(.A0(mai_mai_n457_), .A1(mai_mai_n761_), .B0(mai_mai_n172_), .B1(f), .Y(mai_mai_n937_));
  OAI210     m0909(.A0(mai_mai_n937_), .A1(mai_mai_n460_), .B0(mai_mai_n918_), .Y(mai_mai_n938_));
  NA2        m0910(.A(mai_mai_n860_), .B(mai_mai_n717_), .Y(mai_mai_n939_));
  AN4        m0911(.A(mai_mai_n939_), .B(mai_mai_n938_), .C(mai_mai_n936_), .D(mai_mai_n928_), .Y(mai_mai_n940_));
  NA4        m0912(.A(mai_mai_n940_), .B(mai_mai_n926_), .C(mai_mai_n906_), .D(mai_mai_n855_), .Y(mai12));
  NO2        m0913(.A(mai_mai_n455_), .B(c), .Y(mai_mai_n942_));
  NO4        m0914(.A(mai_mai_n447_), .B(mai_mai_n248_), .C(mai_mai_n594_), .D(mai_mai_n210_), .Y(mai_mai_n943_));
  NA2        m0915(.A(mai_mai_n943_), .B(mai_mai_n942_), .Y(mai_mai_n944_));
  NO2        m0916(.A(mai_mai_n455_), .B(mai_mai_n116_), .Y(mai_mai_n945_));
  NO2        m0917(.A(mai_mai_n863_), .B(mai_mai_n355_), .Y(mai_mai_n946_));
  NO2        m0918(.A(mai_mai_n673_), .B(mai_mai_n382_), .Y(mai_mai_n947_));
  AOI220     m0919(.A0(mai_mai_n947_), .A1(mai_mai_n551_), .B0(mai_mai_n946_), .B1(mai_mai_n945_), .Y(mai_mai_n948_));
  NA3        m0920(.A(mai_mai_n948_), .B(mai_mai_n944_), .C(mai_mai_n446_), .Y(mai_mai_n949_));
  AOI210     m0921(.A0(mai_mai_n230_), .A1(mai_mai_n339_), .B0(mai_mai_n199_), .Y(mai_mai_n950_));
  OR2        m0922(.A(mai_mai_n950_), .B(mai_mai_n943_), .Y(mai_mai_n951_));
  AOI210     m0923(.A0(mai_mai_n336_), .A1(mai_mai_n394_), .B0(mai_mai_n210_), .Y(mai_mai_n952_));
  OAI210     m0924(.A0(mai_mai_n952_), .A1(mai_mai_n951_), .B0(mai_mai_n406_), .Y(mai_mai_n953_));
  NO2        m0925(.A(mai_mai_n653_), .B(mai_mai_n259_), .Y(mai_mai_n954_));
  NO2        m0926(.A(mai_mai_n602_), .B(mai_mai_n856_), .Y(mai_mai_n955_));
  AOI220     m0927(.A0(mai_mai_n955_), .A1(mai_mai_n576_), .B0(mai_mai_n834_), .B1(mai_mai_n954_), .Y(mai_mai_n956_));
  NO2        m0928(.A(mai_mai_n148_), .B(mai_mai_n234_), .Y(mai_mai_n957_));
  NA2        m0929(.A(mai_mai_n956_), .B(mai_mai_n953_), .Y(mai_mai_n958_));
  OR2        m0930(.A(mai_mai_n324_), .B(mai_mai_n945_), .Y(mai_mai_n959_));
  NA2        m0931(.A(mai_mai_n959_), .B(mai_mai_n356_), .Y(mai_mai_n960_));
  NO3        m0932(.A(mai_mai_n130_), .B(mai_mai_n149_), .C(mai_mai_n210_), .Y(mai_mai_n961_));
  NA2        m0933(.A(mai_mai_n961_), .B(mai_mai_n540_), .Y(mai_mai_n962_));
  NA4        m0934(.A(mai_mai_n448_), .B(mai_mai_n440_), .C(mai_mai_n178_), .D(m), .Y(mai_mai_n963_));
  NA3        m0935(.A(mai_mai_n963_), .B(mai_mai_n962_), .C(mai_mai_n960_), .Y(mai_mai_n964_));
  NO3        m0936(.A(mai_mai_n678_), .B(mai_mai_n93_), .C(mai_mai_n45_), .Y(mai_mai_n965_));
  NO4        m0937(.A(mai_mai_n965_), .B(mai_mai_n964_), .C(mai_mai_n958_), .D(mai_mai_n949_), .Y(mai_mai_n966_));
  NO2        m0938(.A(mai_mai_n372_), .B(mai_mai_n371_), .Y(mai_mai_n967_));
  NA2        m0939(.A(mai_mai_n599_), .B(mai_mai_n73_), .Y(mai_mai_n968_));
  NA2        m0940(.A(mai_mai_n563_), .B(mai_mai_n142_), .Y(mai_mai_n969_));
  NOi21      m0941(.An(mai_mai_n34_), .B(mai_mai_n667_), .Y(mai_mai_n970_));
  AOI220     m0942(.A0(mai_mai_n970_), .A1(mai_mai_n969_), .B0(mai_mai_n968_), .B1(mai_mai_n967_), .Y(mai_mai_n971_));
  OAI210     m0943(.A0(mai_mai_n247_), .A1(mai_mai_n45_), .B0(mai_mai_n971_), .Y(mai_mai_n972_));
  NA2        m0944(.A(mai_mai_n438_), .B(mai_mai_n261_), .Y(mai_mai_n973_));
  NO3        m0945(.A(mai_mai_n835_), .B(mai_mai_n91_), .C(mai_mai_n411_), .Y(mai_mai_n974_));
  NAi31      m0946(.An(mai_mai_n974_), .B(mai_mai_n973_), .C(mai_mai_n321_), .Y(mai_mai_n975_));
  NO2        m0947(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n976_));
  NO2        m0948(.A(mai_mai_n511_), .B(mai_mai_n300_), .Y(mai_mai_n977_));
  INV        m0949(.A(mai_mai_n977_), .Y(mai_mai_n978_));
  NO2        m0950(.A(mai_mai_n978_), .B(mai_mai_n142_), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n647_), .B(mai_mai_n365_), .Y(mai_mai_n980_));
  OAI210     m0952(.A0(mai_mai_n748_), .A1(mai_mai_n980_), .B0(mai_mai_n369_), .Y(mai_mai_n981_));
  NO4        m0953(.A(mai_mai_n981_), .B(mai_mai_n979_), .C(mai_mai_n975_), .D(mai_mai_n972_), .Y(mai_mai_n982_));
  NA2        m0954(.A(mai_mai_n348_), .B(m), .Y(mai_mai_n983_));
  NA2        m0955(.A(mai_mai_n159_), .B(i), .Y(mai_mai_n984_));
  NA2        m0956(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n985_));
  OAI220     m0957(.A0(mai_mai_n985_), .A1(mai_mai_n198_), .B0(mai_mai_n984_), .B1(mai_mai_n93_), .Y(mai_mai_n986_));
  AOI210     m0958(.A0(mai_mai_n421_), .A1(mai_mai_n37_), .B0(mai_mai_n986_), .Y(mai_mai_n987_));
  NO2        m0959(.A(mai_mai_n142_), .B(mai_mai_n86_), .Y(mai_mai_n988_));
  OR2        m0960(.A(mai_mai_n988_), .B(mai_mai_n562_), .Y(mai_mai_n989_));
  NA2        m0961(.A(mai_mai_n563_), .B(mai_mai_n386_), .Y(mai_mai_n990_));
  AOI210     m0962(.A0(mai_mai_n990_), .A1(n), .B0(mai_mai_n989_), .Y(mai_mai_n991_));
  OAI220     m0963(.A0(mai_mai_n991_), .A1(mai_mai_n983_), .B0(mai_mai_n987_), .B1(mai_mai_n333_), .Y(mai_mai_n992_));
  NO2        m0964(.A(mai_mai_n673_), .B(mai_mai_n505_), .Y(mai_mai_n993_));
  NA3        m0965(.A(mai_mai_n344_), .B(mai_mai_n644_), .C(i), .Y(mai_mai_n994_));
  OAI210     m0966(.A0(mai_mai_n442_), .A1(mai_mai_n310_), .B0(mai_mai_n994_), .Y(mai_mai_n995_));
  OAI220     m0967(.A0(mai_mai_n995_), .A1(mai_mai_n993_), .B0(mai_mai_n690_), .B1(mai_mai_n772_), .Y(mai_mai_n996_));
  NA2        m0968(.A(mai_mai_n622_), .B(mai_mai_n113_), .Y(mai_mai_n997_));
  OR3        m0969(.A(mai_mai_n310_), .B(mai_mai_n437_), .C(f), .Y(mai_mai_n998_));
  NA3        m0970(.A(mai_mai_n325_), .B(mai_mai_n118_), .C(m), .Y(mai_mai_n999_));
  AOI210     m0971(.A0(mai_mai_n687_), .A1(mai_mai_n999_), .B0(m), .Y(mai_mai_n1000_));
  OAI210     m0972(.A0(mai_mai_n1000_), .A1(mai_mai_n946_), .B0(mai_mai_n324_), .Y(mai_mai_n1001_));
  NA2        m0973(.A(mai_mai_n706_), .B(mai_mai_n894_), .Y(mai_mai_n1002_));
  NA2        m0974(.A(mai_mai_n858_), .B(mai_mai_n443_), .Y(mai_mai_n1003_));
  INV        m0975(.A(mai_mai_n998_), .Y(mai_mai_n1004_));
  AOI220     m0976(.A0(mai_mai_n1004_), .A1(mai_mai_n254_), .B0(mai_mai_n1003_), .B1(mai_mai_n1002_), .Y(mai_mai_n1005_));
  NA3        m0977(.A(mai_mai_n1005_), .B(mai_mai_n1001_), .C(mai_mai_n996_), .Y(mai_mai_n1006_));
  NO2        m0978(.A(mai_mai_n382_), .B(mai_mai_n92_), .Y(mai_mai_n1007_));
  OAI210     m0979(.A0(mai_mai_n1007_), .A1(mai_mai_n954_), .B0(mai_mai_n235_), .Y(mai_mai_n1008_));
  NA2        m0980(.A(mai_mai_n677_), .B(mai_mai_n90_), .Y(mai_mai_n1009_));
  NO2        m0981(.A(mai_mai_n463_), .B(mai_mai_n210_), .Y(mai_mai_n1010_));
  AOI220     m0982(.A0(mai_mai_n1010_), .A1(mai_mai_n387_), .B0(mai_mai_n959_), .B1(mai_mai_n214_), .Y(mai_mai_n1011_));
  NA2        m0983(.A(mai_mai_n947_), .B(mai_mai_n957_), .Y(mai_mai_n1012_));
  NA4        m0984(.A(mai_mai_n1012_), .B(mai_mai_n1011_), .C(mai_mai_n1009_), .D(mai_mai_n1008_), .Y(mai_mai_n1013_));
  OAI210     m0985(.A0(mai_mai_n1003_), .A1(mai_mai_n955_), .B0(mai_mai_n551_), .Y(mai_mai_n1014_));
  AOI210     m0986(.A0(mai_mai_n422_), .A1(mai_mai_n415_), .B0(mai_mai_n835_), .Y(mai_mai_n1015_));
  OAI210     m0987(.A0(mai_mai_n372_), .A1(mai_mai_n371_), .B0(mai_mai_n109_), .Y(mai_mai_n1016_));
  AOI210     m0988(.A0(mai_mai_n1016_), .A1(mai_mai_n544_), .B0(mai_mai_n1015_), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n1000_), .B(mai_mai_n945_), .Y(mai_mai_n1018_));
  NO3        m0990(.A(mai_mai_n908_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n1019_));
  AOI220     m0991(.A0(mai_mai_n1019_), .A1(mai_mai_n642_), .B0(mai_mai_n658_), .B1(mai_mai_n540_), .Y(mai_mai_n1020_));
  NA4        m0992(.A(mai_mai_n1020_), .B(mai_mai_n1018_), .C(mai_mai_n1017_), .D(mai_mai_n1014_), .Y(mai_mai_n1021_));
  NO4        m0993(.A(mai_mai_n1021_), .B(mai_mai_n1013_), .C(mai_mai_n1006_), .D(mai_mai_n992_), .Y(mai_mai_n1022_));
  NAi31      m0994(.An(mai_mai_n139_), .B(mai_mai_n423_), .C(n), .Y(mai_mai_n1023_));
  NO3        m0995(.A(mai_mai_n126_), .B(mai_mai_n342_), .C(mai_mai_n864_), .Y(mai_mai_n1024_));
  NO2        m0996(.A(mai_mai_n1024_), .B(mai_mai_n1023_), .Y(mai_mai_n1025_));
  NO3        m0997(.A(mai_mai_n269_), .B(mai_mai_n139_), .C(mai_mai_n411_), .Y(mai_mai_n1026_));
  AOI210     m0998(.A0(mai_mai_n1026_), .A1(mai_mai_n506_), .B0(mai_mai_n1025_), .Y(mai_mai_n1027_));
  NA2        m0999(.A(mai_mai_n499_), .B(i), .Y(mai_mai_n1028_));
  NA2        m1000(.A(mai_mai_n1028_), .B(mai_mai_n1027_), .Y(mai_mai_n1029_));
  NA2        m1001(.A(mai_mai_n227_), .B(mai_mai_n168_), .Y(mai_mai_n1030_));
  NO3        m1002(.A(mai_mai_n307_), .B(mai_mai_n448_), .C(mai_mai_n172_), .Y(mai_mai_n1031_));
  NOi31      m1003(.An(mai_mai_n1030_), .B(mai_mai_n1031_), .C(mai_mai_n210_), .Y(mai_mai_n1032_));
  NAi21      m1004(.An(mai_mai_n563_), .B(mai_mai_n1010_), .Y(mai_mai_n1033_));
  NA2        m1005(.A(mai_mai_n441_), .B(mai_mai_n894_), .Y(mai_mai_n1034_));
  NO3        m1006(.A(mai_mai_n442_), .B(mai_mai_n310_), .C(mai_mai_n75_), .Y(mai_mai_n1035_));
  AOI220     m1007(.A0(mai_mai_n1035_), .A1(mai_mai_n1034_), .B0(mai_mai_n488_), .B1(m), .Y(mai_mai_n1036_));
  NA2        m1008(.A(mai_mai_n1036_), .B(mai_mai_n1033_), .Y(mai_mai_n1037_));
  OAI220     m1009(.A0(mai_mai_n1023_), .A1(mai_mai_n230_), .B0(mai_mai_n994_), .B1(mai_mai_n617_), .Y(mai_mai_n1038_));
  NO2        m1010(.A(mai_mai_n674_), .B(mai_mai_n382_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n950_), .B(mai_mai_n942_), .Y(mai_mai_n1040_));
  NO3        m1012(.A(mai_mai_n552_), .B(mai_mai_n146_), .C(mai_mai_n209_), .Y(mai_mai_n1041_));
  OAI210     m1013(.A0(mai_mai_n1041_), .A1(mai_mai_n534_), .B0(mai_mai_n383_), .Y(mai_mai_n1042_));
  OAI220     m1014(.A0(mai_mai_n947_), .A1(mai_mai_n955_), .B0(mai_mai_n553_), .B1(mai_mai_n431_), .Y(mai_mai_n1043_));
  NA4        m1015(.A(mai_mai_n1043_), .B(mai_mai_n1042_), .C(mai_mai_n1040_), .D(mai_mai_n636_), .Y(mai_mai_n1044_));
  OAI210     m1016(.A0(mai_mai_n950_), .A1(mai_mai_n943_), .B0(mai_mai_n1030_), .Y(mai_mai_n1045_));
  NA3        m1017(.A(mai_mai_n990_), .B(mai_mai_n493_), .C(mai_mai_n46_), .Y(mai_mai_n1046_));
  INV        m1018(.A(mai_mai_n332_), .Y(mai_mai_n1047_));
  NA4        m1019(.A(mai_mai_n1047_), .B(mai_mai_n1046_), .C(mai_mai_n1045_), .D(mai_mai_n270_), .Y(mai_mai_n1048_));
  OR4        m1020(.A(mai_mai_n1048_), .B(mai_mai_n1044_), .C(mai_mai_n1039_), .D(mai_mai_n1038_), .Y(mai_mai_n1049_));
  NO4        m1021(.A(mai_mai_n1049_), .B(mai_mai_n1037_), .C(mai_mai_n1032_), .D(mai_mai_n1029_), .Y(mai_mai_n1050_));
  NA4        m1022(.A(mai_mai_n1050_), .B(mai_mai_n1022_), .C(mai_mai_n982_), .D(mai_mai_n966_), .Y(mai13));
  NA2        m1023(.A(mai_mai_n46_), .B(mai_mai_n89_), .Y(mai_mai_n1052_));
  AN2        m1024(.A(c), .B(b), .Y(mai_mai_n1053_));
  NA3        m1025(.A(mai_mai_n246_), .B(mai_mai_n1053_), .C(m), .Y(mai_mai_n1054_));
  NA2        m1026(.A(mai_mai_n504_), .B(f), .Y(mai_mai_n1055_));
  NO4        m1027(.A(mai_mai_n1055_), .B(mai_mai_n1054_), .C(mai_mai_n1052_), .D(mai_mai_n595_), .Y(mai_mai_n1056_));
  NA2        m1028(.A(mai_mai_n261_), .B(mai_mai_n1053_), .Y(mai_mai_n1057_));
  NO4        m1029(.A(mai_mai_n1057_), .B(mai_mai_n1055_), .C(mai_mai_n984_), .D(a), .Y(mai_mai_n1058_));
  NAi32      m1030(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1059_));
  NA2        m1031(.A(mai_mai_n138_), .B(mai_mai_n45_), .Y(mai_mai_n1060_));
  NO4        m1032(.A(mai_mai_n1060_), .B(mai_mai_n1059_), .C(mai_mai_n602_), .D(mai_mai_n306_), .Y(mai_mai_n1061_));
  NA2        m1033(.A(mai_mai_n681_), .B(mai_mai_n221_), .Y(mai_mai_n1062_));
  NA2        m1034(.A(mai_mai_n414_), .B(mai_mai_n209_), .Y(mai_mai_n1063_));
  AN2        m1035(.A(d), .B(c), .Y(mai_mai_n1064_));
  NA2        m1036(.A(mai_mai_n1064_), .B(mai_mai_n116_), .Y(mai_mai_n1065_));
  NO4        m1037(.A(mai_mai_n1065_), .B(mai_mai_n1063_), .C(mai_mai_n173_), .D(mai_mai_n164_), .Y(mai_mai_n1066_));
  NA2        m1038(.A(mai_mai_n504_), .B(c), .Y(mai_mai_n1067_));
  NO4        m1039(.A(mai_mai_n1060_), .B(mai_mai_n598_), .C(mai_mai_n1067_), .D(mai_mai_n306_), .Y(mai_mai_n1068_));
  AO210      m1040(.A0(mai_mai_n1066_), .A1(mai_mai_n1062_), .B0(mai_mai_n1068_), .Y(mai_mai_n1069_));
  OR4        m1041(.A(mai_mai_n1069_), .B(mai_mai_n1061_), .C(mai_mai_n1058_), .D(mai_mai_n1056_), .Y(mai_mai_n1070_));
  NAi32      m1042(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1071_));
  NO2        m1043(.A(mai_mai_n1071_), .B(mai_mai_n143_), .Y(mai_mai_n1072_));
  NA2        m1044(.A(mai_mai_n1072_), .B(m), .Y(mai_mai_n1073_));
  OR3        m1045(.A(mai_mai_n221_), .B(mai_mai_n173_), .C(mai_mai_n164_), .Y(mai_mai_n1074_));
  NO2        m1046(.A(mai_mai_n1074_), .B(mai_mai_n1073_), .Y(mai_mai_n1075_));
  NO2        m1047(.A(mai_mai_n1067_), .B(mai_mai_n306_), .Y(mai_mai_n1076_));
  NO2        m1048(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1077_));
  NA2        m1049(.A(mai_mai_n646_), .B(mai_mai_n1077_), .Y(mai_mai_n1078_));
  NOi21      m1050(.An(mai_mai_n1076_), .B(mai_mai_n1078_), .Y(mai_mai_n1079_));
  NO2        m1051(.A(mai_mai_n776_), .B(mai_mai_n112_), .Y(mai_mai_n1080_));
  NOi41      m1052(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1081_));
  NA2        m1053(.A(mai_mai_n1081_), .B(mai_mai_n1080_), .Y(mai_mai_n1082_));
  NO2        m1054(.A(mai_mai_n1082_), .B(mai_mai_n1073_), .Y(mai_mai_n1083_));
  OR3        m1055(.A(e), .B(d), .C(c), .Y(mai_mai_n1084_));
  NA3        m1056(.A(k), .B(j), .C(i), .Y(mai_mai_n1085_));
  NO3        m1057(.A(mai_mai_n1085_), .B(mai_mai_n306_), .C(mai_mai_n92_), .Y(mai_mai_n1086_));
  NOi21      m1058(.An(mai_mai_n1086_), .B(mai_mai_n1084_), .Y(mai_mai_n1087_));
  OR4        m1059(.A(mai_mai_n1087_), .B(mai_mai_n1083_), .C(mai_mai_n1079_), .D(mai_mai_n1075_), .Y(mai_mai_n1088_));
  NA3        m1060(.A(mai_mai_n471_), .B(mai_mai_n335_), .C(mai_mai_n56_), .Y(mai_mai_n1089_));
  NO2        m1061(.A(mai_mai_n1089_), .B(mai_mai_n1078_), .Y(mai_mai_n1090_));
  NO4        m1062(.A(mai_mai_n1089_), .B(mai_mai_n598_), .C(mai_mai_n454_), .D(mai_mai_n45_), .Y(mai_mai_n1091_));
  NO2        m1063(.A(f), .B(c), .Y(mai_mai_n1092_));
  NOi21      m1064(.An(mai_mai_n1092_), .B(mai_mai_n447_), .Y(mai_mai_n1093_));
  NA2        m1065(.A(mai_mai_n1093_), .B(mai_mai_n59_), .Y(mai_mai_n1094_));
  OR2        m1066(.A(k), .B(i), .Y(mai_mai_n1095_));
  NO3        m1067(.A(mai_mai_n1095_), .B(mai_mai_n241_), .C(l), .Y(mai_mai_n1096_));
  NOi31      m1068(.An(mai_mai_n1096_), .B(mai_mai_n1094_), .C(j), .Y(mai_mai_n1097_));
  OR3        m1069(.A(mai_mai_n1097_), .B(mai_mai_n1091_), .C(mai_mai_n1090_), .Y(mai_mai_n1098_));
  OR3        m1070(.A(mai_mai_n1098_), .B(mai_mai_n1088_), .C(mai_mai_n1070_), .Y(mai02));
  OR2        m1071(.A(l), .B(k), .Y(mai_mai_n1100_));
  OR3        m1072(.A(h), .B(m), .C(f), .Y(mai_mai_n1101_));
  OR3        m1073(.A(n), .B(m), .C(i), .Y(mai_mai_n1102_));
  NO4        m1074(.A(mai_mai_n1102_), .B(mai_mai_n1101_), .C(mai_mai_n1100_), .D(mai_mai_n1084_), .Y(mai_mai_n1103_));
  NOi31      m1075(.An(e), .B(d), .C(c), .Y(mai_mai_n1104_));
  AOI210     m1076(.A0(mai_mai_n1086_), .A1(mai_mai_n1104_), .B0(mai_mai_n1061_), .Y(mai_mai_n1105_));
  AN3        m1077(.A(m), .B(f), .C(c), .Y(mai_mai_n1106_));
  NA3        m1078(.A(mai_mai_n1106_), .B(mai_mai_n471_), .C(h), .Y(mai_mai_n1107_));
  OR2        m1079(.A(mai_mai_n1085_), .B(mai_mai_n306_), .Y(mai_mai_n1108_));
  OR2        m1080(.A(mai_mai_n1108_), .B(mai_mai_n1107_), .Y(mai_mai_n1109_));
  NO3        m1081(.A(mai_mai_n1089_), .B(mai_mai_n1060_), .C(mai_mai_n598_), .Y(mai_mai_n1110_));
  NO2        m1082(.A(mai_mai_n1110_), .B(mai_mai_n1075_), .Y(mai_mai_n1111_));
  NA3        m1083(.A(l), .B(k), .C(j), .Y(mai_mai_n1112_));
  NA2        m1084(.A(i), .B(h), .Y(mai_mai_n1113_));
  NO3        m1085(.A(mai_mai_n1113_), .B(mai_mai_n1112_), .C(mai_mai_n130_), .Y(mai_mai_n1114_));
  NO3        m1086(.A(mai_mai_n140_), .B(mai_mai_n282_), .C(mai_mai_n210_), .Y(mai_mai_n1115_));
  AOI210     m1087(.A0(mai_mai_n1115_), .A1(mai_mai_n1114_), .B0(mai_mai_n1079_), .Y(mai_mai_n1116_));
  NA3        m1088(.A(c), .B(b), .C(a), .Y(mai_mai_n1117_));
  NO3        m1089(.A(mai_mai_n1117_), .B(mai_mai_n917_), .C(mai_mai_n209_), .Y(mai_mai_n1118_));
  NO4        m1090(.A(mai_mai_n1085_), .B(mai_mai_n300_), .C(mai_mai_n49_), .D(mai_mai_n112_), .Y(mai_mai_n1119_));
  AOI210     m1091(.A0(mai_mai_n1119_), .A1(mai_mai_n1118_), .B0(mai_mai_n1090_), .Y(mai_mai_n1120_));
  AN4        m1092(.A(mai_mai_n1120_), .B(mai_mai_n1116_), .C(mai_mai_n1111_), .D(mai_mai_n1109_), .Y(mai_mai_n1121_));
  NO2        m1093(.A(mai_mai_n1065_), .B(mai_mai_n1063_), .Y(mai_mai_n1122_));
  NA2        m1094(.A(mai_mai_n1082_), .B(mai_mai_n1074_), .Y(mai_mai_n1123_));
  AOI210     m1095(.A0(mai_mai_n1123_), .A1(mai_mai_n1122_), .B0(mai_mai_n1056_), .Y(mai_mai_n1124_));
  NAi41      m1096(.An(mai_mai_n1103_), .B(mai_mai_n1124_), .C(mai_mai_n1121_), .D(mai_mai_n1105_), .Y(mai03));
  INV        m1097(.A(mai_mai_n373_), .Y(mai_mai_n1126_));
  NO2        m1098(.A(mai_mai_n1126_), .B(mai_mai_n1016_), .Y(mai_mai_n1127_));
  NOi31      m1099(.An(mai_mai_n821_), .B(mai_mai_n869_), .C(mai_mai_n859_), .Y(mai_mai_n1128_));
  OAI220     m1100(.A0(mai_mai_n1128_), .A1(mai_mai_n706_), .B0(mai_mai_n1127_), .B1(mai_mai_n599_), .Y(mai_mai_n1129_));
  NOi31      m1101(.An(i), .B(k), .C(j), .Y(mai_mai_n1130_));
  NA4        m1102(.A(mai_mai_n1130_), .B(mai_mai_n1104_), .C(mai_mai_n344_), .D(mai_mai_n335_), .Y(mai_mai_n1131_));
  OAI210     m1103(.A0(mai_mai_n835_), .A1(mai_mai_n424_), .B0(mai_mai_n1131_), .Y(mai_mai_n1132_));
  NOi31      m1104(.An(m), .B(n), .C(f), .Y(mai_mai_n1133_));
  NA2        m1105(.A(mai_mai_n1133_), .B(mai_mai_n51_), .Y(mai_mai_n1134_));
  AN2        m1106(.A(e), .B(c), .Y(mai_mai_n1135_));
  NA2        m1107(.A(mai_mai_n1135_), .B(a), .Y(mai_mai_n1136_));
  OAI220     m1108(.A0(mai_mai_n1136_), .A1(mai_mai_n1134_), .B0(mai_mai_n901_), .B1(mai_mai_n430_), .Y(mai_mai_n1137_));
  NA2        m1109(.A(mai_mai_n515_), .B(l), .Y(mai_mai_n1138_));
  NOi31      m1110(.An(mai_mai_n880_), .B(mai_mai_n1054_), .C(mai_mai_n1138_), .Y(mai_mai_n1139_));
  NO4        m1111(.A(mai_mai_n1139_), .B(mai_mai_n1137_), .C(mai_mai_n1132_), .D(mai_mai_n1015_), .Y(mai_mai_n1140_));
  NO2        m1112(.A(mai_mai_n282_), .B(a), .Y(mai_mai_n1141_));
  INV        m1113(.A(mai_mai_n1061_), .Y(mai_mai_n1142_));
  NO2        m1114(.A(mai_mai_n1113_), .B(mai_mai_n491_), .Y(mai_mai_n1143_));
  NO2        m1115(.A(mai_mai_n89_), .B(m), .Y(mai_mai_n1144_));
  AOI210     m1116(.A0(mai_mai_n1144_), .A1(mai_mai_n1143_), .B0(mai_mai_n1096_), .Y(mai_mai_n1145_));
  OR2        m1117(.A(mai_mai_n1145_), .B(mai_mai_n1094_), .Y(mai_mai_n1146_));
  NA3        m1118(.A(mai_mai_n1146_), .B(mai_mai_n1142_), .C(mai_mai_n1140_), .Y(mai_mai_n1147_));
  NO4        m1119(.A(mai_mai_n1147_), .B(mai_mai_n1129_), .C(mai_mai_n836_), .D(mai_mai_n575_), .Y(mai_mai_n1148_));
  NA2        m1120(.A(c), .B(b), .Y(mai_mai_n1149_));
  NO2        m1121(.A(mai_mai_n716_), .B(mai_mai_n1149_), .Y(mai_mai_n1150_));
  OAI210     m1122(.A0(mai_mai_n878_), .A1(mai_mai_n851_), .B0(mai_mai_n417_), .Y(mai_mai_n1151_));
  OAI210     m1123(.A0(mai_mai_n1151_), .A1(mai_mai_n879_), .B0(mai_mai_n1150_), .Y(mai_mai_n1152_));
  NAi21      m1124(.An(mai_mai_n425_), .B(mai_mai_n1150_), .Y(mai_mai_n1153_));
  NA3        m1125(.A(mai_mai_n431_), .B(mai_mai_n568_), .C(f), .Y(mai_mai_n1154_));
  OAI210     m1126(.A0(mai_mai_n557_), .A1(mai_mai_n39_), .B0(mai_mai_n1141_), .Y(mai_mai_n1155_));
  NA3        m1127(.A(mai_mai_n1155_), .B(mai_mai_n1154_), .C(mai_mai_n1153_), .Y(mai_mai_n1156_));
  NA2        m1128(.A(mai_mai_n257_), .B(mai_mai_n119_), .Y(mai_mai_n1157_));
  OAI210     m1129(.A0(mai_mai_n1157_), .A1(mai_mai_n286_), .B0(m), .Y(mai_mai_n1158_));
  NAi21      m1130(.An(f), .B(d), .Y(mai_mai_n1159_));
  NO2        m1131(.A(mai_mai_n1159_), .B(mai_mai_n1117_), .Y(mai_mai_n1160_));
  INV        m1132(.A(mai_mai_n1160_), .Y(mai_mai_n1161_));
  NO2        m1133(.A(mai_mai_n1158_), .B(mai_mai_n1161_), .Y(mai_mai_n1162_));
  AOI210     m1134(.A0(mai_mai_n1162_), .A1(mai_mai_n113_), .B0(mai_mai_n1156_), .Y(mai_mai_n1163_));
  NO2        m1135(.A(mai_mai_n179_), .B(mai_mai_n234_), .Y(mai_mai_n1164_));
  NA2        m1136(.A(mai_mai_n1164_), .B(m), .Y(mai_mai_n1165_));
  NA3        m1137(.A(mai_mai_n934_), .B(mai_mai_n1138_), .C(mai_mai_n477_), .Y(mai_mai_n1166_));
  NA2        m1138(.A(mai_mai_n1166_), .B(mai_mai_n475_), .Y(mai_mai_n1167_));
  NO2        m1139(.A(mai_mai_n1167_), .B(mai_mai_n1165_), .Y(mai_mai_n1168_));
  NA2        m1140(.A(mai_mai_n570_), .B(mai_mai_n413_), .Y(mai_mai_n1169_));
  NA2        m1141(.A(mai_mai_n155_), .B(mai_mai_n33_), .Y(mai_mai_n1170_));
  AOI210     m1142(.A0(mai_mai_n980_), .A1(mai_mai_n1170_), .B0(mai_mai_n210_), .Y(mai_mai_n1171_));
  OAI210     m1143(.A0(mai_mai_n1171_), .A1(mai_mai_n451_), .B0(mai_mai_n1160_), .Y(mai_mai_n1172_));
  NO2        m1144(.A(mai_mai_n376_), .B(mai_mai_n375_), .Y(mai_mai_n1173_));
  AOI210     m1145(.A0(mai_mai_n1164_), .A1(mai_mai_n433_), .B0(mai_mai_n974_), .Y(mai_mai_n1174_));
  NAi41      m1146(.An(mai_mai_n1173_), .B(mai_mai_n1174_), .C(mai_mai_n1172_), .D(mai_mai_n1169_), .Y(mai_mai_n1175_));
  NO2        m1147(.A(mai_mai_n1175_), .B(mai_mai_n1168_), .Y(mai_mai_n1176_));
  NA4        m1148(.A(mai_mai_n1176_), .B(mai_mai_n1163_), .C(mai_mai_n1152_), .D(mai_mai_n1148_), .Y(mai00));
  AOI210     m1149(.A0(mai_mai_n299_), .A1(mai_mai_n210_), .B0(mai_mai_n274_), .Y(mai_mai_n1178_));
  NO2        m1150(.A(mai_mai_n1178_), .B(mai_mai_n589_), .Y(mai_mai_n1179_));
  AOI210     m1151(.A0(mai_mai_n914_), .A1(mai_mai_n957_), .B0(mai_mai_n1132_), .Y(mai_mai_n1180_));
  NO2        m1152(.A(mai_mai_n1110_), .B(mai_mai_n974_), .Y(mai_mai_n1181_));
  NA3        m1153(.A(mai_mai_n1181_), .B(mai_mai_n1180_), .C(mai_mai_n1017_), .Y(mai_mai_n1182_));
  NA2        m1154(.A(mai_mai_n517_), .B(f), .Y(mai_mai_n1183_));
  OAI210     m1155(.A0(mai_mai_n1024_), .A1(mai_mai_n40_), .B0(mai_mai_n660_), .Y(mai_mai_n1184_));
  NA3        m1156(.A(mai_mai_n1184_), .B(mai_mai_n253_), .C(n), .Y(mai_mai_n1185_));
  AOI210     m1157(.A0(mai_mai_n1185_), .A1(mai_mai_n1183_), .B0(mai_mai_n1065_), .Y(mai_mai_n1186_));
  NO4        m1158(.A(mai_mai_n1186_), .B(mai_mai_n1182_), .C(mai_mai_n1179_), .D(mai_mai_n1088_), .Y(mai_mai_n1187_));
  NA3        m1159(.A(mai_mai_n163_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1188_));
  NA3        m1160(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1189_));
  NOi31      m1161(.An(n), .B(m), .C(i), .Y(mai_mai_n1190_));
  NA3        m1162(.A(mai_mai_n1190_), .B(mai_mai_n663_), .C(mai_mai_n51_), .Y(mai_mai_n1191_));
  OAI210     m1163(.A0(mai_mai_n1189_), .A1(mai_mai_n1188_), .B0(mai_mai_n1191_), .Y(mai_mai_n1192_));
  INV        m1164(.A(mai_mai_n588_), .Y(mai_mai_n1193_));
  NO3        m1165(.A(mai_mai_n1193_), .B(mai_mai_n1192_), .C(mai_mai_n1173_), .Y(mai_mai_n1194_));
  NO4        m1166(.A(mai_mai_n494_), .B(mai_mai_n358_), .C(mai_mai_n1149_), .D(mai_mai_n59_), .Y(mai_mai_n1195_));
  NA3        m1167(.A(mai_mai_n388_), .B(mai_mai_n217_), .C(m), .Y(mai_mai_n1196_));
  OA220      m1168(.A0(mai_mai_n1196_), .A1(mai_mai_n1189_), .B0(mai_mai_n389_), .B1(mai_mai_n133_), .Y(mai_mai_n1197_));
  NO2        m1169(.A(h), .B(m), .Y(mai_mai_n1198_));
  NA4        m1170(.A(mai_mai_n506_), .B(mai_mai_n471_), .C(mai_mai_n1198_), .D(mai_mai_n1053_), .Y(mai_mai_n1199_));
  NA2        m1171(.A(mai_mai_n961_), .B(mai_mai_n587_), .Y(mai_mai_n1200_));
  NA3        m1172(.A(mai_mai_n1200_), .B(mai_mai_n1199_), .C(mai_mai_n1197_), .Y(mai_mai_n1201_));
  NO3        m1173(.A(mai_mai_n1201_), .B(mai_mai_n1195_), .C(mai_mai_n263_), .Y(mai_mai_n1202_));
  NO2        m1174(.A(mai_mai_n236_), .B(mai_mai_n178_), .Y(mai_mai_n1203_));
  NA2        m1175(.A(mai_mai_n1203_), .B(mai_mai_n431_), .Y(mai_mai_n1204_));
  NA3        m1176(.A(mai_mai_n176_), .B(mai_mai_n112_), .C(m), .Y(mai_mai_n1205_));
  NA3        m1177(.A(mai_mai_n471_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1206_));
  NOi31      m1178(.An(mai_mai_n887_), .B(mai_mai_n1206_), .C(mai_mai_n1205_), .Y(mai_mai_n1207_));
  NAi31      m1179(.An(mai_mai_n183_), .B(mai_mai_n875_), .C(mai_mai_n471_), .Y(mai_mai_n1208_));
  NAi31      m1180(.An(mai_mai_n1207_), .B(mai_mai_n1208_), .C(mai_mai_n1204_), .Y(mai_mai_n1209_));
  INV        m1181(.A(mai_mai_n1103_), .Y(mai_mai_n1210_));
  NAi31      m1182(.An(mai_mai_n1068_), .B(mai_mai_n1210_), .C(mai_mai_n74_), .Y(mai_mai_n1211_));
  NO4        m1183(.A(mai_mai_n1211_), .B(mai_mai_n1209_), .C(mai_mai_n590_), .D(mai_mai_n527_), .Y(mai_mai_n1212_));
  AN3        m1184(.A(mai_mai_n1212_), .B(mai_mai_n1202_), .C(mai_mai_n1194_), .Y(mai_mai_n1213_));
  NA3        m1185(.A(mai_mai_n1133_), .B(mai_mai_n622_), .C(mai_mai_n470_), .Y(mai_mai_n1214_));
  NA3        m1186(.A(mai_mai_n1214_), .B(mai_mai_n571_), .C(mai_mai_n239_), .Y(mai_mai_n1215_));
  OAI210     m1187(.A0(mai_mai_n469_), .A1(mai_mai_n120_), .B0(mai_mai_n881_), .Y(mai_mai_n1216_));
  AOI220     m1188(.A0(mai_mai_n1216_), .A1(mai_mai_n1166_), .B0(mai_mai_n570_), .B1(mai_mai_n413_), .Y(mai_mai_n1217_));
  OR4        m1189(.A(mai_mai_n1065_), .B(mai_mai_n269_), .C(mai_mai_n219_), .D(e), .Y(mai_mai_n1218_));
  NO2        m1190(.A(mai_mai_n213_), .B(mai_mai_n210_), .Y(mai_mai_n1219_));
  NA2        m1191(.A(n), .B(e), .Y(mai_mai_n1220_));
  NO2        m1192(.A(mai_mai_n1220_), .B(mai_mai_n143_), .Y(mai_mai_n1221_));
  AOI220     m1193(.A0(mai_mai_n1221_), .A1(mai_mai_n271_), .B0(mai_mai_n862_), .B1(mai_mai_n1219_), .Y(mai_mai_n1222_));
  OAI210     m1194(.A0(mai_mai_n359_), .A1(mai_mai_n312_), .B0(mai_mai_n453_), .Y(mai_mai_n1223_));
  NA4        m1195(.A(mai_mai_n1223_), .B(mai_mai_n1222_), .C(mai_mai_n1218_), .D(mai_mai_n1217_), .Y(mai_mai_n1224_));
  AOI210     m1196(.A0(mai_mai_n1221_), .A1(mai_mai_n866_), .B0(mai_mai_n836_), .Y(mai_mai_n1225_));
  AOI220     m1197(.A0(mai_mai_n970_), .A1(mai_mai_n587_), .B0(mai_mai_n663_), .B1(mai_mai_n242_), .Y(mai_mai_n1226_));
  NO2        m1198(.A(mai_mai_n68_), .B(h), .Y(mai_mai_n1227_));
  NO3        m1199(.A(mai_mai_n1065_), .B(mai_mai_n1063_), .C(mai_mai_n740_), .Y(mai_mai_n1228_));
  NO2        m1200(.A(mai_mai_n1100_), .B(mai_mai_n130_), .Y(mai_mai_n1229_));
  AN2        m1201(.A(mai_mai_n1229_), .B(mai_mai_n1115_), .Y(mai_mai_n1230_));
  OAI210     m1202(.A0(mai_mai_n1230_), .A1(mai_mai_n1228_), .B0(mai_mai_n1227_), .Y(mai_mai_n1231_));
  NA4        m1203(.A(mai_mai_n1231_), .B(mai_mai_n1226_), .C(mai_mai_n1225_), .D(mai_mai_n882_), .Y(mai_mai_n1232_));
  NO4        m1204(.A(mai_mai_n1232_), .B(mai_mai_n1224_), .C(mai_mai_n295_), .D(mai_mai_n1215_), .Y(mai_mai_n1233_));
  NA2        m1205(.A(mai_mai_n852_), .B(mai_mai_n771_), .Y(mai_mai_n1234_));
  NA4        m1206(.A(mai_mai_n1234_), .B(mai_mai_n1233_), .C(mai_mai_n1213_), .D(mai_mai_n1187_), .Y(mai01));
  AN2        m1207(.A(mai_mai_n1042_), .B(mai_mai_n1040_), .Y(mai_mai_n1236_));
  NO4        m1208(.A(mai_mai_n817_), .B(mai_mai_n809_), .C(mai_mai_n485_), .D(mai_mai_n280_), .Y(mai_mai_n1237_));
  NO2        m1209(.A(mai_mai_n604_), .B(mai_mai_n289_), .Y(mai_mai_n1238_));
  OAI210     m1210(.A0(mai_mai_n1238_), .A1(mai_mai_n399_), .B0(i), .Y(mai_mai_n1239_));
  NA3        m1211(.A(mai_mai_n1239_), .B(mai_mai_n1237_), .C(mai_mai_n1236_), .Y(mai_mai_n1240_));
  NA2        m1212(.A(mai_mai_n563_), .B(mai_mai_n268_), .Y(mai_mai_n1241_));
  NA2        m1213(.A(mai_mai_n977_), .B(mai_mai_n1241_), .Y(mai_mai_n1242_));
  NA3        m1214(.A(mai_mai_n1242_), .B(mai_mai_n930_), .C(mai_mai_n334_), .Y(mai_mai_n1243_));
  NA2        m1215(.A(mai_mai_n45_), .B(f), .Y(mai_mai_n1244_));
  NA2        m1216(.A(mai_mai_n723_), .B(mai_mai_n97_), .Y(mai_mai_n1245_));
  OAI220     m1217(.A0(mai_mai_n1245_), .A1(mai_mai_n1244_), .B0(mai_mai_n355_), .B1(mai_mai_n284_), .Y(mai_mai_n1246_));
  NA2        m1218(.A(mai_mai_n118_), .B(l), .Y(mai_mai_n1247_));
  OA220      m1219(.A0(mai_mai_n1247_), .A1(mai_mai_n597_), .B0(mai_mai_n675_), .B1(mai_mai_n373_), .Y(mai_mai_n1248_));
  NAi31      m1220(.An(mai_mai_n158_), .B(mai_mai_n1248_), .C(mai_mai_n913_), .Y(mai_mai_n1249_));
  NO3        m1221(.A(mai_mai_n797_), .B(mai_mai_n689_), .C(mai_mai_n520_), .Y(mai_mai_n1250_));
  NA4        m1222(.A(mai_mai_n723_), .B(mai_mai_n97_), .C(mai_mai_n45_), .D(mai_mai_n209_), .Y(mai_mai_n1251_));
  OA220      m1223(.A0(mai_mai_n1251_), .A1(mai_mai_n684_), .B0(mai_mai_n193_), .B1(mai_mai_n191_), .Y(mai_mai_n1252_));
  NA3        m1224(.A(mai_mai_n1252_), .B(mai_mai_n1250_), .C(mai_mai_n136_), .Y(mai_mai_n1253_));
  NO4        m1225(.A(mai_mai_n1253_), .B(mai_mai_n1249_), .C(mai_mai_n1243_), .D(mai_mai_n1240_), .Y(mai_mai_n1254_));
  INV        m1226(.A(mai_mai_n1196_), .Y(mai_mai_n1255_));
  NA2        m1227(.A(mai_mai_n1255_), .B(mai_mai_n540_), .Y(mai_mai_n1256_));
  NA2        m1228(.A(mai_mai_n546_), .B(mai_mai_n401_), .Y(mai_mai_n1257_));
  NA2        m1229(.A(mai_mai_n76_), .B(i), .Y(mai_mai_n1258_));
  AOI210     m1230(.A0(mai_mai_n603_), .A1(mai_mai_n597_), .B0(mai_mai_n1258_), .Y(mai_mai_n1259_));
  NOi21      m1231(.An(mai_mai_n572_), .B(mai_mai_n594_), .Y(mai_mai_n1260_));
  AOI210     m1232(.A0(mai_mai_n1260_), .A1(mai_mai_n1257_), .B0(mai_mai_n1259_), .Y(mai_mai_n1261_));
  AOI210     m1233(.A0(mai_mai_n202_), .A1(mai_mai_n91_), .B0(mai_mai_n209_), .Y(mai_mai_n1262_));
  OAI210     m1234(.A0(mai_mai_n824_), .A1(mai_mai_n431_), .B0(mai_mai_n1262_), .Y(mai_mai_n1263_));
  AN3        m1235(.A(m), .B(l), .C(k), .Y(mai_mai_n1264_));
  OAI210     m1236(.A0(mai_mai_n361_), .A1(mai_mai_n34_), .B0(mai_mai_n1264_), .Y(mai_mai_n1265_));
  OR2        m1237(.A(mai_mai_n1265_), .B(mai_mai_n333_), .Y(mai_mai_n1266_));
  NA4        m1238(.A(mai_mai_n1266_), .B(mai_mai_n1263_), .C(mai_mai_n1261_), .D(mai_mai_n1256_), .Y(mai_mai_n1267_));
  AOI210     m1239(.A0(mai_mai_n609_), .A1(mai_mai_n118_), .B0(mai_mai_n615_), .Y(mai_mai_n1268_));
  OAI210     m1240(.A0(mai_mai_n1247_), .A1(mai_mai_n606_), .B0(mai_mai_n1268_), .Y(mai_mai_n1269_));
  NA2        m1241(.A(mai_mai_n279_), .B(mai_mai_n193_), .Y(mai_mai_n1270_));
  OAI210     m1242(.A0(mai_mai_n1270_), .A1(mai_mai_n390_), .B0(mai_mai_n680_), .Y(mai_mai_n1271_));
  NO3        m1243(.A(mai_mai_n835_), .B(mai_mai_n202_), .C(mai_mai_n411_), .Y(mai_mai_n1272_));
  NO2        m1244(.A(mai_mai_n1272_), .B(mai_mai_n974_), .Y(mai_mai_n1273_));
  OAI210     m1245(.A0(mai_mai_n1246_), .A1(mai_mai_n327_), .B0(mai_mai_n690_), .Y(mai_mai_n1274_));
  NA4        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1273_), .C(mai_mai_n1271_), .D(mai_mai_n800_), .Y(mai_mai_n1275_));
  NO3        m1247(.A(mai_mai_n1275_), .B(mai_mai_n1269_), .C(mai_mai_n1267_), .Y(mai_mai_n1276_));
  NA2        m1248(.A(mai_mai_n512_), .B(mai_mai_n58_), .Y(mai_mai_n1277_));
  NA3        m1249(.A(mai_mai_n754_), .B(mai_mai_n76_), .C(i), .Y(mai_mai_n1278_));
  AOI210     m1250(.A0(mai_mai_n1278_), .A1(mai_mai_n1251_), .B0(mai_mai_n997_), .Y(mai_mai_n1279_));
  NO2        m1251(.A(mai_mai_n1279_), .B(mai_mai_n1192_), .Y(mai_mai_n1280_));
  NA3        m1252(.A(mai_mai_n1280_), .B(mai_mai_n1277_), .C(mai_mai_n770_), .Y(mai_mai_n1281_));
  NO2        m1253(.A(mai_mai_n984_), .B(mai_mai_n229_), .Y(mai_mai_n1282_));
  NO2        m1254(.A(mai_mai_n985_), .B(mai_mai_n565_), .Y(mai_mai_n1283_));
  OAI210     m1255(.A0(mai_mai_n1283_), .A1(mai_mai_n1282_), .B0(mai_mai_n342_), .Y(mai_mai_n1284_));
  NA2        m1256(.A(mai_mai_n582_), .B(mai_mai_n580_), .Y(mai_mai_n1285_));
  NO3        m1257(.A(mai_mai_n81_), .B(mai_mai_n300_), .C(mai_mai_n45_), .Y(mai_mai_n1286_));
  NA2        m1258(.A(mai_mai_n1286_), .B(mai_mai_n562_), .Y(mai_mai_n1287_));
  NA2        m1259(.A(mai_mai_n1287_), .B(mai_mai_n1285_), .Y(mai_mai_n1288_));
  OR2        m1260(.A(mai_mai_n1196_), .B(mai_mai_n1189_), .Y(mai_mai_n1289_));
  NO2        m1261(.A(mai_mai_n373_), .B(mai_mai_n73_), .Y(mai_mai_n1290_));
  AOI210     m1262(.A0(mai_mai_n745_), .A1(mai_mai_n633_), .B0(mai_mai_n1290_), .Y(mai_mai_n1291_));
  NA2        m1263(.A(mai_mai_n1286_), .B(mai_mai_n827_), .Y(mai_mai_n1292_));
  NA4        m1264(.A(mai_mai_n1292_), .B(mai_mai_n1291_), .C(mai_mai_n1289_), .D(mai_mai_n391_), .Y(mai_mai_n1293_));
  NOi41      m1265(.An(mai_mai_n1284_), .B(mai_mai_n1293_), .C(mai_mai_n1288_), .D(mai_mai_n1281_), .Y(mai_mai_n1294_));
  NO2        m1266(.A(mai_mai_n129_), .B(mai_mai_n45_), .Y(mai_mai_n1295_));
  NO2        m1267(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1296_));
  AO220      m1268(.A0(mai_mai_n1296_), .A1(mai_mai_n639_), .B0(mai_mai_n1295_), .B1(mai_mai_n721_), .Y(mai_mai_n1297_));
  NA2        m1269(.A(mai_mai_n1297_), .B(mai_mai_n342_), .Y(mai_mai_n1298_));
  NO3        m1270(.A(mai_mai_n1113_), .B(mai_mai_n173_), .C(mai_mai_n89_), .Y(mai_mai_n1299_));
  NA2        m1271(.A(mai_mai_n1286_), .B(mai_mai_n988_), .Y(mai_mai_n1300_));
  NA2        m1272(.A(mai_mai_n1300_), .B(mai_mai_n1298_), .Y(mai_mai_n1301_));
  NO2        m1273(.A(mai_mai_n630_), .B(mai_mai_n629_), .Y(mai_mai_n1302_));
  NO4        m1274(.A(mai_mai_n1113_), .B(mai_mai_n1302_), .C(mai_mai_n171_), .D(mai_mai_n89_), .Y(mai_mai_n1303_));
  NO3        m1275(.A(mai_mai_n1303_), .B(mai_mai_n1301_), .C(mai_mai_n652_), .Y(mai_mai_n1304_));
  NA4        m1276(.A(mai_mai_n1304_), .B(mai_mai_n1294_), .C(mai_mai_n1276_), .D(mai_mai_n1254_), .Y(mai06));
  NO2        m1277(.A(mai_mai_n412_), .B(mai_mai_n569_), .Y(mai_mai_n1306_));
  NO2        m1278(.A(mai_mai_n747_), .B(i), .Y(mai_mai_n1307_));
  OAI210     m1279(.A0(mai_mai_n1307_), .A1(mai_mai_n264_), .B0(mai_mai_n1306_), .Y(mai_mai_n1308_));
  NO2        m1280(.A(mai_mai_n221_), .B(mai_mai_n102_), .Y(mai_mai_n1309_));
  OAI210     m1281(.A0(mai_mai_n1309_), .A1(mai_mai_n1299_), .B0(mai_mai_n387_), .Y(mai_mai_n1310_));
  NO3        m1282(.A(mai_mai_n613_), .B(mai_mai_n822_), .C(mai_mai_n616_), .Y(mai_mai_n1311_));
  OR2        m1283(.A(mai_mai_n1311_), .B(mai_mai_n901_), .Y(mai_mai_n1312_));
  NA4        m1284(.A(mai_mai_n1312_), .B(mai_mai_n1310_), .C(mai_mai_n1308_), .D(mai_mai_n1284_), .Y(mai_mai_n1313_));
  NO3        m1285(.A(mai_mai_n1313_), .B(mai_mai_n1288_), .C(mai_mai_n252_), .Y(mai_mai_n1314_));
  NO2        m1286(.A(mai_mai_n300_), .B(mai_mai_n45_), .Y(mai_mai_n1315_));
  AOI210     m1287(.A0(mai_mai_n1315_), .A1(mai_mai_n989_), .B0(mai_mai_n1282_), .Y(mai_mai_n1316_));
  AOI210     m1288(.A0(mai_mai_n1315_), .A1(mai_mai_n566_), .B0(mai_mai_n1297_), .Y(mai_mai_n1317_));
  AOI210     m1289(.A0(mai_mai_n1317_), .A1(mai_mai_n1316_), .B0(mai_mai_n339_), .Y(mai_mai_n1318_));
  OAI210     m1290(.A0(mai_mai_n91_), .A1(mai_mai_n40_), .B0(mai_mai_n688_), .Y(mai_mai_n1319_));
  NA2        m1291(.A(mai_mai_n1319_), .B(mai_mai_n656_), .Y(mai_mai_n1320_));
  NO2        m1292(.A(mai_mai_n523_), .B(mai_mai_n168_), .Y(mai_mai_n1321_));
  NOi21      m1293(.An(mai_mai_n135_), .B(mai_mai_n45_), .Y(mai_mai_n1322_));
  NO2        m1294(.A(mai_mai_n623_), .B(mai_mai_n1134_), .Y(mai_mai_n1323_));
  OAI210     m1295(.A0(mai_mai_n464_), .A1(mai_mai_n245_), .B0(mai_mai_n924_), .Y(mai_mai_n1324_));
  NO4        m1296(.A(mai_mai_n1324_), .B(mai_mai_n1323_), .C(mai_mai_n1322_), .D(mai_mai_n1321_), .Y(mai_mai_n1325_));
  OR2        m1297(.A(mai_mai_n614_), .B(mai_mai_n612_), .Y(mai_mai_n1326_));
  NO2        m1298(.A(mai_mai_n372_), .B(mai_mai_n134_), .Y(mai_mai_n1327_));
  AOI210     m1299(.A0(mai_mai_n1327_), .A1(mai_mai_n600_), .B0(mai_mai_n1326_), .Y(mai_mai_n1328_));
  NA3        m1300(.A(mai_mai_n1328_), .B(mai_mai_n1325_), .C(mai_mai_n1320_), .Y(mai_mai_n1329_));
  NO2        m1301(.A(mai_mai_n762_), .B(mai_mai_n371_), .Y(mai_mai_n1330_));
  NO2        m1302(.A(mai_mai_n690_), .B(mai_mai_n772_), .Y(mai_mai_n1331_));
  NOi21      m1303(.An(mai_mai_n1330_), .B(mai_mai_n1331_), .Y(mai_mai_n1332_));
  AN2        m1304(.A(mai_mai_n970_), .B(mai_mai_n659_), .Y(mai_mai_n1333_));
  NO4        m1305(.A(mai_mai_n1333_), .B(mai_mai_n1332_), .C(mai_mai_n1329_), .D(mai_mai_n1318_), .Y(mai_mai_n1334_));
  NO2        m1306(.A(mai_mai_n816_), .B(mai_mai_n275_), .Y(mai_mai_n1335_));
  OAI220     m1307(.A0(mai_mai_n747_), .A1(mai_mai_n47_), .B0(mai_mai_n221_), .B1(mai_mai_n632_), .Y(mai_mai_n1336_));
  AOI220     m1308(.A0(mai_mai_n364_), .A1(mai_mai_n1336_), .B0(mai_mai_n1335_), .B1(mai_mai_n264_), .Y(mai_mai_n1337_));
  NO3        m1309(.A(mai_mai_n241_), .B(mai_mai_n102_), .C(mai_mai_n282_), .Y(mai_mai_n1338_));
  OAI220     m1310(.A0(mai_mai_n713_), .A1(mai_mai_n245_), .B0(mai_mai_n519_), .B1(mai_mai_n523_), .Y(mai_mai_n1339_));
  OAI210     m1311(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1340_));
  NO3        m1312(.A(mai_mai_n1340_), .B(mai_mai_n611_), .C(j), .Y(mai_mai_n1341_));
  NOi21      m1313(.An(mai_mai_n1341_), .B(mai_mai_n684_), .Y(mai_mai_n1342_));
  NO4        m1314(.A(mai_mai_n1342_), .B(mai_mai_n1339_), .C(mai_mai_n1338_), .D(mai_mai_n1137_), .Y(mai_mai_n1343_));
  NA4        m1315(.A(mai_mai_n807_), .B(mai_mai_n806_), .C(mai_mai_n441_), .D(mai_mai_n894_), .Y(mai_mai_n1344_));
  NAi31      m1316(.An(mai_mai_n762_), .B(mai_mai_n1344_), .C(mai_mai_n201_), .Y(mai_mai_n1345_));
  NA4        m1317(.A(mai_mai_n1345_), .B(mai_mai_n1343_), .C(mai_mai_n1337_), .D(mai_mai_n1226_), .Y(mai_mai_n1346_));
  NOi31      m1318(.An(mai_mai_n1311_), .B(mai_mai_n468_), .C(mai_mai_n400_), .Y(mai_mai_n1347_));
  OR3        m1319(.A(mai_mai_n1347_), .B(mai_mai_n796_), .C(mai_mai_n549_), .Y(mai_mai_n1348_));
  OR3        m1320(.A(mai_mai_n375_), .B(mai_mai_n221_), .C(mai_mai_n632_), .Y(mai_mai_n1349_));
  AOI210     m1321(.A0(mai_mai_n582_), .A1(mai_mai_n453_), .B0(mai_mai_n377_), .Y(mai_mai_n1350_));
  NA3        m1322(.A(mai_mai_n1350_), .B(mai_mai_n1349_), .C(mai_mai_n1348_), .Y(mai_mai_n1351_));
  NA2        m1323(.A(mai_mai_n1327_), .B(mai_mai_n235_), .Y(mai_mai_n1352_));
  AN2        m1324(.A(mai_mai_n943_), .B(mai_mai_n942_), .Y(mai_mai_n1353_));
  NO4        m1325(.A(mai_mai_n1353_), .B(mai_mai_n892_), .C(mai_mai_n508_), .D(mai_mai_n488_), .Y(mai_mai_n1354_));
  NA3        m1326(.A(mai_mai_n1354_), .B(mai_mai_n1352_), .C(mai_mai_n1292_), .Y(mai_mai_n1355_));
  NAi21      m1327(.An(j), .B(i), .Y(mai_mai_n1356_));
  NO4        m1328(.A(mai_mai_n1302_), .B(mai_mai_n1356_), .C(mai_mai_n447_), .D(mai_mai_n232_), .Y(mai_mai_n1357_));
  NO4        m1329(.A(mai_mai_n1357_), .B(mai_mai_n1355_), .C(mai_mai_n1351_), .D(mai_mai_n1346_), .Y(mai_mai_n1358_));
  NA4        m1330(.A(mai_mai_n1358_), .B(mai_mai_n1334_), .C(mai_mai_n1314_), .D(mai_mai_n1304_), .Y(mai07));
  NAi32      m1331(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1360_));
  NO3        m1332(.A(mai_mai_n1360_), .B(m), .C(f), .Y(mai_mai_n1361_));
  OAI210     m1333(.A0(mai_mai_n322_), .A1(mai_mai_n490_), .B0(mai_mai_n1361_), .Y(mai_mai_n1362_));
  NAi21      m1334(.An(f), .B(c), .Y(mai_mai_n1363_));
  OR2        m1335(.A(e), .B(d), .Y(mai_mai_n1364_));
  OAI220     m1336(.A0(mai_mai_n1364_), .A1(mai_mai_n1363_), .B0(mai_mai_n645_), .B1(mai_mai_n323_), .Y(mai_mai_n1365_));
  NA3        m1337(.A(mai_mai_n1365_), .B(mai_mai_n1077_), .C(mai_mai_n176_), .Y(mai_mai_n1366_));
  NOi31      m1338(.An(n), .B(m), .C(b), .Y(mai_mai_n1367_));
  NO3        m1339(.A(mai_mai_n130_), .B(mai_mai_n454_), .C(h), .Y(mai_mai_n1368_));
  NA2        m1340(.A(mai_mai_n1366_), .B(mai_mai_n1362_), .Y(mai_mai_n1369_));
  NOi41      m1341(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1370_));
  NOi21      m1342(.An(h), .B(k), .Y(mai_mai_n1371_));
  NO2        m1343(.A(k), .B(i), .Y(mai_mai_n1372_));
  NA3        m1344(.A(mai_mai_n1372_), .B(mai_mai_n912_), .C(mai_mai_n176_), .Y(mai_mai_n1373_));
  NA2        m1345(.A(mai_mai_n89_), .B(mai_mai_n45_), .Y(mai_mai_n1374_));
  NO2        m1346(.A(mai_mai_n1071_), .B(mai_mai_n447_), .Y(mai_mai_n1375_));
  NA3        m1347(.A(mai_mai_n1375_), .B(mai_mai_n1374_), .C(mai_mai_n210_), .Y(mai_mai_n1376_));
  NO2        m1348(.A(mai_mai_n1085_), .B(mai_mai_n306_), .Y(mai_mai_n1377_));
  NA2        m1349(.A(mai_mai_n550_), .B(mai_mai_n82_), .Y(mai_mai_n1378_));
  NA2        m1350(.A(mai_mai_n1227_), .B(mai_mai_n290_), .Y(mai_mai_n1379_));
  NA4        m1351(.A(mai_mai_n1379_), .B(mai_mai_n1378_), .C(mai_mai_n1376_), .D(mai_mai_n1373_), .Y(mai_mai_n1380_));
  NO2        m1352(.A(mai_mai_n1380_), .B(mai_mai_n1369_), .Y(mai_mai_n1381_));
  NO3        m1353(.A(e), .B(d), .C(c), .Y(mai_mai_n1382_));
  NA2        m1354(.A(mai_mai_n1566_), .B(mai_mai_n1382_), .Y(mai_mai_n1383_));
  NO2        m1355(.A(mai_mai_n1383_), .B(mai_mai_n210_), .Y(mai_mai_n1384_));
  OR2        m1356(.A(h), .B(f), .Y(mai_mai_n1385_));
  NO3        m1357(.A(n), .B(m), .C(i), .Y(mai_mai_n1386_));
  OAI210     m1358(.A0(mai_mai_n1135_), .A1(mai_mai_n153_), .B0(mai_mai_n1386_), .Y(mai_mai_n1387_));
  NO2        m1359(.A(mai_mai_n1387_), .B(mai_mai_n1385_), .Y(mai_mai_n1388_));
  NA3        m1360(.A(mai_mai_n710_), .B(mai_mai_n698_), .C(mai_mai_n112_), .Y(mai_mai_n1389_));
  NO2        m1361(.A(mai_mai_n1389_), .B(mai_mai_n45_), .Y(mai_mai_n1390_));
  NA2        m1362(.A(mai_mai_n1386_), .B(mai_mai_n654_), .Y(mai_mai_n1391_));
  NO2        m1363(.A(l), .B(k), .Y(mai_mai_n1392_));
  NOi41      m1364(.An(mai_mai_n555_), .B(mai_mai_n1392_), .C(mai_mai_n483_), .D(mai_mai_n447_), .Y(mai_mai_n1393_));
  NO3        m1365(.A(mai_mai_n447_), .B(d), .C(c), .Y(mai_mai_n1394_));
  NO4        m1366(.A(mai_mai_n1393_), .B(mai_mai_n1390_), .C(mai_mai_n1388_), .D(mai_mai_n1384_), .Y(mai_mai_n1395_));
  NO2        m1367(.A(mai_mai_n144_), .B(h), .Y(mai_mai_n1396_));
  NO2        m1368(.A(mai_mai_n1095_), .B(l), .Y(mai_mai_n1397_));
  NO2        m1369(.A(m), .B(c), .Y(mai_mai_n1398_));
  NA3        m1370(.A(mai_mai_n1398_), .B(mai_mai_n140_), .C(mai_mai_n184_), .Y(mai_mai_n1399_));
  NO2        m1371(.A(mai_mai_n1399_), .B(mai_mai_n1397_), .Y(mai_mai_n1400_));
  NA2        m1372(.A(mai_mai_n1400_), .B(mai_mai_n176_), .Y(mai_mai_n1401_));
  OAI210     m1373(.A0(mai_mai_n1371_), .A1(mai_mai_n209_), .B0(mai_mai_n1095_), .Y(mai_mai_n1402_));
  NO2        m1374(.A(mai_mai_n455_), .B(a), .Y(mai_mai_n1403_));
  NA3        m1375(.A(mai_mai_n1403_), .B(mai_mai_n1402_), .C(mai_mai_n113_), .Y(mai_mai_n1404_));
  NO2        m1376(.A(i), .B(h), .Y(mai_mai_n1405_));
  AOI210     m1377(.A0(mai_mai_n1159_), .A1(h), .B0(mai_mai_n418_), .Y(mai_mai_n1406_));
  NA2        m1378(.A(mai_mai_n137_), .B(mai_mai_n217_), .Y(mai_mai_n1407_));
  NO2        m1379(.A(mai_mai_n1407_), .B(mai_mai_n1406_), .Y(mai_mai_n1408_));
  NO2        m1380(.A(mai_mai_n768_), .B(mai_mai_n185_), .Y(mai_mai_n1409_));
  NOi31      m1381(.An(m), .B(n), .C(b), .Y(mai_mai_n1410_));
  NOi31      m1382(.An(f), .B(d), .C(c), .Y(mai_mai_n1411_));
  NA2        m1383(.A(mai_mai_n1411_), .B(mai_mai_n1410_), .Y(mai_mai_n1412_));
  INV        m1384(.A(mai_mai_n1412_), .Y(mai_mai_n1413_));
  NO3        m1385(.A(mai_mai_n1413_), .B(mai_mai_n1409_), .C(mai_mai_n1408_), .Y(mai_mai_n1414_));
  NA2        m1386(.A(mai_mai_n1106_), .B(mai_mai_n471_), .Y(mai_mai_n1415_));
  NO4        m1387(.A(mai_mai_n1415_), .B(mai_mai_n1080_), .C(mai_mai_n447_), .D(mai_mai_n45_), .Y(mai_mai_n1416_));
  OAI210     m1388(.A0(mai_mai_n179_), .A1(mai_mai_n535_), .B0(mai_mai_n1081_), .Y(mai_mai_n1417_));
  NO3        m1389(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1418_));
  INV        m1390(.A(mai_mai_n1417_), .Y(mai_mai_n1419_));
  NO2        m1391(.A(mai_mai_n1419_), .B(mai_mai_n1416_), .Y(mai_mai_n1420_));
  AN4        m1392(.A(mai_mai_n1420_), .B(mai_mai_n1414_), .C(mai_mai_n1404_), .D(mai_mai_n1401_), .Y(mai_mai_n1421_));
  NA2        m1393(.A(mai_mai_n1367_), .B(mai_mai_n384_), .Y(mai_mai_n1422_));
  NO2        m1394(.A(mai_mai_n1422_), .B(mai_mai_n1062_), .Y(mai_mai_n1423_));
  NA2        m1395(.A(mai_mai_n1394_), .B(mai_mai_n211_), .Y(mai_mai_n1424_));
  NO2        m1396(.A(mai_mai_n185_), .B(b), .Y(mai_mai_n1425_));
  AOI220     m1397(.A0(mai_mai_n1190_), .A1(mai_mai_n1425_), .B0(mai_mai_n1114_), .B1(mai_mai_n1415_), .Y(mai_mai_n1426_));
  NAi31      m1398(.An(mai_mai_n1423_), .B(mai_mai_n1426_), .C(mai_mai_n1424_), .Y(mai_mai_n1427_));
  NO4        m1399(.A(mai_mai_n130_), .B(m), .C(f), .D(e), .Y(mai_mai_n1428_));
  NA3        m1400(.A(mai_mai_n1372_), .B(mai_mai_n291_), .C(h), .Y(mai_mai_n1429_));
  NA2        m1401(.A(mai_mai_n192_), .B(mai_mai_n99_), .Y(mai_mai_n1430_));
  OR2        m1402(.A(e), .B(a), .Y(mai_mai_n1431_));
  NO2        m1403(.A(mai_mai_n1364_), .B(mai_mai_n1363_), .Y(mai_mai_n1432_));
  AOI210     m1404(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1432_), .Y(mai_mai_n1433_));
  NO2        m1405(.A(mai_mai_n1433_), .B(mai_mai_n1102_), .Y(mai_mai_n1434_));
  NOi41      m1406(.An(h), .B(f), .C(e), .D(a), .Y(mai_mai_n1435_));
  NA2        m1407(.A(mai_mai_n1435_), .B(mai_mai_n113_), .Y(mai_mai_n1436_));
  NA2        m1408(.A(mai_mai_n1370_), .B(mai_mai_n1392_), .Y(mai_mai_n1437_));
  NA2        m1409(.A(mai_mai_n1437_), .B(mai_mai_n1436_), .Y(mai_mai_n1438_));
  OR3        m1410(.A(mai_mai_n549_), .B(mai_mai_n548_), .C(mai_mai_n112_), .Y(mai_mai_n1439_));
  NA2        m1411(.A(mai_mai_n1133_), .B(mai_mai_n411_), .Y(mai_mai_n1440_));
  OAI220     m1412(.A0(mai_mai_n1440_), .A1(mai_mai_n440_), .B0(mai_mai_n1439_), .B1(mai_mai_n300_), .Y(mai_mai_n1441_));
  AO210      m1413(.A0(mai_mai_n1441_), .A1(mai_mai_n116_), .B0(mai_mai_n1438_), .Y(mai_mai_n1442_));
  NO3        m1414(.A(mai_mai_n1442_), .B(mai_mai_n1434_), .C(mai_mai_n1427_), .Y(mai_mai_n1443_));
  NA4        m1415(.A(mai_mai_n1443_), .B(mai_mai_n1421_), .C(mai_mai_n1395_), .D(mai_mai_n1381_), .Y(mai_mai_n1444_));
  NO2        m1416(.A(mai_mai_n1149_), .B(mai_mai_n110_), .Y(mai_mai_n1445_));
  NA2        m1417(.A(mai_mai_n384_), .B(mai_mai_n56_), .Y(mai_mai_n1446_));
  AOI210     m1418(.A0(mai_mai_n1446_), .A1(mai_mai_n1071_), .B0(mai_mai_n1391_), .Y(mai_mai_n1447_));
  NA2        m1419(.A(mai_mai_n211_), .B(mai_mai_n176_), .Y(mai_mai_n1448_));
  AOI210     m1420(.A0(mai_mai_n1448_), .A1(mai_mai_n1205_), .B0(mai_mai_n1446_), .Y(mai_mai_n1449_));
  NO2        m1421(.A(mai_mai_n1107_), .B(mai_mai_n1102_), .Y(mai_mai_n1450_));
  NO3        m1422(.A(mai_mai_n1450_), .B(mai_mai_n1449_), .C(mai_mai_n1447_), .Y(mai_mai_n1451_));
  NO2        m1423(.A(mai_mai_n396_), .B(j), .Y(mai_mai_n1452_));
  NA3        m1424(.A(mai_mai_n1418_), .B(mai_mai_n1364_), .C(mai_mai_n1133_), .Y(mai_mai_n1453_));
  NAi41      m1425(.An(mai_mai_n1405_), .B(mai_mai_n1093_), .C(mai_mai_n164_), .D(mai_mai_n147_), .Y(mai_mai_n1454_));
  NA2        m1426(.A(mai_mai_n1454_), .B(mai_mai_n1453_), .Y(mai_mai_n1455_));
  NA3        m1427(.A(m), .B(mai_mai_n1452_), .C(mai_mai_n155_), .Y(mai_mai_n1456_));
  INV        m1428(.A(mai_mai_n1456_), .Y(mai_mai_n1457_));
  NO3        m1429(.A(mai_mai_n762_), .B(mai_mai_n171_), .C(mai_mai_n414_), .Y(mai_mai_n1458_));
  NO3        m1430(.A(mai_mai_n1458_), .B(mai_mai_n1457_), .C(mai_mai_n1455_), .Y(mai_mai_n1459_));
  AOI210     m1431(.A0(mai_mai_n1448_), .A1(mai_mai_n1430_), .B0(mai_mai_n1071_), .Y(mai_mai_n1460_));
  OR2        m1432(.A(n), .B(i), .Y(mai_mai_n1461_));
  OAI210     m1433(.A0(mai_mai_n1461_), .A1(mai_mai_n1092_), .B0(mai_mai_n49_), .Y(mai_mai_n1462_));
  AOI220     m1434(.A0(mai_mai_n1462_), .A1(mai_mai_n1198_), .B0(mai_mai_n839_), .B1(mai_mai_n192_), .Y(mai_mai_n1463_));
  INV        m1435(.A(mai_mai_n1463_), .Y(mai_mai_n1464_));
  OAI220     m1436(.A0(mai_mai_n681_), .A1(m), .B0(mai_mai_n221_), .B1(c), .Y(mai_mai_n1465_));
  AOI210     m1437(.A0(mai_mai_n1425_), .A1(mai_mai_n41_), .B0(mai_mai_n1465_), .Y(mai_mai_n1466_));
  NO2        m1438(.A(mai_mai_n130_), .B(l), .Y(mai_mai_n1467_));
  NO2        m1439(.A(mai_mai_n221_), .B(k), .Y(mai_mai_n1468_));
  OAI210     m1440(.A0(mai_mai_n1468_), .A1(mai_mai_n1405_), .B0(mai_mai_n1467_), .Y(mai_mai_n1469_));
  OAI220     m1441(.A0(mai_mai_n1469_), .A1(mai_mai_n31_), .B0(mai_mai_n1466_), .B1(mai_mai_n173_), .Y(mai_mai_n1470_));
  NO3        m1442(.A(mai_mai_n1439_), .B(mai_mai_n471_), .C(mai_mai_n355_), .Y(mai_mai_n1471_));
  NO4        m1443(.A(mai_mai_n1471_), .B(mai_mai_n1470_), .C(mai_mai_n1464_), .D(mai_mai_n1460_), .Y(mai_mai_n1472_));
  NO3        m1444(.A(mai_mai_n1117_), .B(mai_mai_n1364_), .C(mai_mai_n49_), .Y(mai_mai_n1473_));
  NO2        m1445(.A(mai_mai_n1102_), .B(h), .Y(mai_mai_n1474_));
  NA3        m1446(.A(mai_mai_n1474_), .B(d), .C(mai_mai_n1063_), .Y(mai_mai_n1475_));
  NO2        m1447(.A(mai_mai_n1475_), .B(c), .Y(mai_mai_n1476_));
  NA3        m1448(.A(mai_mai_n1445_), .B(mai_mai_n471_), .C(f), .Y(mai_mai_n1477_));
  NA2        m1449(.A(mai_mai_n176_), .B(mai_mai_n112_), .Y(mai_mai_n1478_));
  NO2        m1450(.A(mai_mai_n42_), .B(mai_mai_n1477_), .Y(mai_mai_n1479_));
  NO2        m1451(.A(mai_mai_n1356_), .B(mai_mai_n171_), .Y(mai_mai_n1480_));
  NOi21      m1452(.An(d), .B(f), .Y(mai_mai_n1481_));
  NO3        m1453(.A(mai_mai_n1411_), .B(mai_mai_n1481_), .C(mai_mai_n40_), .Y(mai_mai_n1482_));
  NA2        m1454(.A(mai_mai_n1482_), .B(mai_mai_n1480_), .Y(mai_mai_n1483_));
  NO2        m1455(.A(mai_mai_n1364_), .B(f), .Y(mai_mai_n1484_));
  INV        m1456(.A(mai_mai_n1483_), .Y(mai_mai_n1485_));
  NO3        m1457(.A(mai_mai_n1485_), .B(mai_mai_n1479_), .C(mai_mai_n1476_), .Y(mai_mai_n1486_));
  NA4        m1458(.A(mai_mai_n1486_), .B(mai_mai_n1472_), .C(mai_mai_n1459_), .D(mai_mai_n1451_), .Y(mai_mai_n1487_));
  NO3        m1459(.A(mai_mai_n1106_), .B(mai_mai_n1092_), .C(mai_mai_n40_), .Y(mai_mai_n1488_));
  NO2        m1460(.A(mai_mai_n471_), .B(mai_mai_n300_), .Y(mai_mai_n1489_));
  OAI210     m1461(.A0(mai_mai_n1489_), .A1(mai_mai_n1488_), .B0(mai_mai_n1377_), .Y(mai_mai_n1490_));
  OAI210     m1462(.A0(mai_mai_n1428_), .A1(mai_mai_n1367_), .B0(mai_mai_n898_), .Y(mai_mai_n1491_));
  OAI220     m1463(.A0(mai_mai_n1059_), .A1(mai_mai_n130_), .B0(mai_mai_n681_), .B1(mai_mai_n171_), .Y(mai_mai_n1492_));
  NA2        m1464(.A(mai_mai_n1492_), .B(mai_mai_n638_), .Y(mai_mai_n1493_));
  NA3        m1465(.A(mai_mai_n1493_), .B(mai_mai_n1491_), .C(mai_mai_n1490_), .Y(mai_mai_n1494_));
  NA2        m1466(.A(mai_mai_n1398_), .B(mai_mai_n1481_), .Y(mai_mai_n1495_));
  NO2        m1467(.A(mai_mai_n1495_), .B(m), .Y(mai_mai_n1496_));
  NO2        m1468(.A(mai_mai_n148_), .B(mai_mai_n178_), .Y(mai_mai_n1497_));
  OAI210     m1469(.A0(mai_mai_n1497_), .A1(mai_mai_n110_), .B0(mai_mai_n1410_), .Y(mai_mai_n1498_));
  INV        m1470(.A(mai_mai_n1498_), .Y(mai_mai_n1499_));
  NO3        m1471(.A(mai_mai_n1499_), .B(mai_mai_n1496_), .C(mai_mai_n1494_), .Y(mai_mai_n1500_));
  NO2        m1472(.A(mai_mai_n1363_), .B(e), .Y(mai_mai_n1501_));
  NA2        m1473(.A(mai_mai_n1501_), .B(mai_mai_n409_), .Y(mai_mai_n1502_));
  OAI210     m1474(.A0(mai_mai_n1484_), .A1(mai_mai_n1144_), .B0(mai_mai_n647_), .Y(mai_mai_n1503_));
  OR3        m1475(.A(mai_mai_n1468_), .B(mai_mai_n1227_), .C(mai_mai_n130_), .Y(mai_mai_n1504_));
  OAI220     m1476(.A0(mai_mai_n1504_), .A1(mai_mai_n1502_), .B0(mai_mai_n1503_), .B1(mai_mai_n449_), .Y(mai_mai_n1505_));
  INV        m1477(.A(mai_mai_n1505_), .Y(mai_mai_n1506_));
  NO2        m1478(.A(mai_mai_n178_), .B(c), .Y(mai_mai_n1507_));
  OAI210     m1479(.A0(mai_mai_n1507_), .A1(mai_mai_n1501_), .B0(mai_mai_n176_), .Y(mai_mai_n1508_));
  AOI220     m1480(.A0(mai_mai_n1508_), .A1(mai_mai_n1094_), .B0(mai_mai_n542_), .B1(mai_mai_n371_), .Y(mai_mai_n1509_));
  NA2        m1481(.A(mai_mai_n548_), .B(m), .Y(mai_mai_n1510_));
  AOI210     m1482(.A0(mai_mai_n1510_), .A1(mai_mai_n1394_), .B0(mai_mai_n1473_), .Y(mai_mai_n1511_));
  NO2        m1483(.A(mai_mai_n1431_), .B(f), .Y(mai_mai_n1512_));
  NA2        m1484(.A(mai_mai_n1144_), .B(a), .Y(mai_mai_n1513_));
  OAI220     m1485(.A0(mai_mai_n1513_), .A1(mai_mai_n69_), .B0(mai_mai_n1511_), .B1(mai_mai_n209_), .Y(mai_mai_n1514_));
  AOI210     m1486(.A0(mai_mai_n917_), .A1(mai_mai_n420_), .B0(mai_mai_n104_), .Y(mai_mai_n1515_));
  OR2        m1487(.A(mai_mai_n1515_), .B(mai_mai_n548_), .Y(mai_mai_n1516_));
  NA2        m1488(.A(mai_mai_n1512_), .B(mai_mai_n1374_), .Y(mai_mai_n1517_));
  OAI220     m1489(.A0(mai_mai_n1517_), .A1(mai_mai_n49_), .B0(mai_mai_n1516_), .B1(mai_mai_n171_), .Y(mai_mai_n1518_));
  NA4        m1490(.A(mai_mai_n1115_), .B(mai_mai_n1112_), .C(mai_mai_n217_), .D(mai_mai_n68_), .Y(mai_mai_n1519_));
  NA2        m1491(.A(mai_mai_n1368_), .B(mai_mai_n179_), .Y(mai_mai_n1520_));
  NO2        m1492(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1521_));
  OAI210     m1493(.A0(mai_mai_n1431_), .A1(mai_mai_n877_), .B0(mai_mai_n490_), .Y(mai_mai_n1522_));
  OAI210     m1494(.A0(mai_mai_n1522_), .A1(mai_mai_n1118_), .B0(mai_mai_n1521_), .Y(mai_mai_n1523_));
  NO2        m1495(.A(mai_mai_n248_), .B(m), .Y(mai_mai_n1524_));
  NO2        m1496(.A(m), .B(i), .Y(mai_mai_n1525_));
  BUFFER     m1497(.A(mai_mai_n1525_), .Y(mai_mai_n1526_));
  AOI220     m1498(.A0(mai_mai_n1526_), .A1(mai_mai_n1396_), .B0(mai_mai_n1093_), .B1(mai_mai_n1524_), .Y(mai_mai_n1527_));
  NA4        m1499(.A(mai_mai_n1527_), .B(mai_mai_n1523_), .C(mai_mai_n1520_), .D(mai_mai_n1519_), .Y(mai_mai_n1528_));
  NO4        m1500(.A(mai_mai_n1528_), .B(mai_mai_n1518_), .C(mai_mai_n1514_), .D(mai_mai_n1509_), .Y(mai_mai_n1529_));
  NA3        m1501(.A(mai_mai_n1529_), .B(mai_mai_n1506_), .C(mai_mai_n1500_), .Y(mai_mai_n1530_));
  NA3        m1502(.A(mai_mai_n976_), .B(mai_mai_n137_), .C(mai_mai_n46_), .Y(mai_mai_n1531_));
  AOI210     m1503(.A0(mai_mai_n145_), .A1(c), .B0(mai_mai_n1531_), .Y(mai_mai_n1532_));
  INV        m1504(.A(mai_mai_n182_), .Y(mai_mai_n1533_));
  NA2        m1505(.A(mai_mai_n1533_), .B(mai_mai_n1474_), .Y(mai_mai_n1534_));
  AO210      m1506(.A0(mai_mai_n131_), .A1(l), .B0(mai_mai_n1422_), .Y(mai_mai_n1535_));
  NO2        m1507(.A(mai_mai_n72_), .B(c), .Y(mai_mai_n1536_));
  NA2        m1508(.A(mai_mai_n1480_), .B(mai_mai_n1536_), .Y(mai_mai_n1537_));
  NA3        m1509(.A(mai_mai_n1537_), .B(mai_mai_n1535_), .C(mai_mai_n1534_), .Y(mai_mai_n1538_));
  NO2        m1510(.A(mai_mai_n1538_), .B(mai_mai_n1532_), .Y(mai_mai_n1539_));
  AOI210     m1511(.A0(mai_mai_n153_), .A1(mai_mai_n56_), .B0(mai_mai_n1501_), .Y(mai_mai_n1540_));
  NO2        m1512(.A(mai_mai_n1540_), .B(mai_mai_n1478_), .Y(mai_mai_n1541_));
  NOi21      m1513(.An(mai_mai_n1368_), .B(e), .Y(mai_mai_n1542_));
  NO2        m1514(.A(mai_mai_n1542_), .B(mai_mai_n1541_), .Y(mai_mai_n1543_));
  AN2        m1515(.A(mai_mai_n1115_), .B(mai_mai_n1100_), .Y(mai_mai_n1544_));
  AOI220     m1516(.A0(mai_mai_n1525_), .A1(mai_mai_n654_), .B0(mai_mai_n1077_), .B1(mai_mai_n156_), .Y(mai_mai_n1545_));
  NOi31      m1517(.An(mai_mai_n30_), .B(mai_mai_n1545_), .C(n), .Y(mai_mai_n1546_));
  AOI210     m1518(.A0(mai_mai_n1544_), .A1(mai_mai_n1190_), .B0(mai_mai_n1546_), .Y(mai_mai_n1547_));
  NO2        m1519(.A(mai_mai_n1477_), .B(mai_mai_n69_), .Y(mai_mai_n1548_));
  NA2        m1520(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1549_));
  NO2        m1521(.A(mai_mai_n1372_), .B(mai_mai_n118_), .Y(mai_mai_n1550_));
  OAI220     m1522(.A0(mai_mai_n1550_), .A1(mai_mai_n1422_), .B0(mai_mai_n1440_), .B1(mai_mai_n1549_), .Y(mai_mai_n1551_));
  NO2        m1523(.A(mai_mai_n1551_), .B(mai_mai_n1548_), .Y(mai_mai_n1552_));
  NA4        m1524(.A(mai_mai_n1552_), .B(mai_mai_n1547_), .C(mai_mai_n1543_), .D(mai_mai_n1539_), .Y(mai_mai_n1553_));
  OR4        m1525(.A(mai_mai_n1553_), .B(mai_mai_n1530_), .C(mai_mai_n1487_), .D(mai_mai_n1444_), .Y(mai04));
  NOi31      m1526(.An(mai_mai_n1428_), .B(mai_mai_n1429_), .C(mai_mai_n1065_), .Y(mai_mai_n1555_));
  NA2        m1527(.A(mai_mai_n1484_), .B(mai_mai_n839_), .Y(mai_mai_n1556_));
  NO4        m1528(.A(mai_mai_n1556_), .B(mai_mai_n1054_), .C(mai_mai_n491_), .D(j), .Y(mai_mai_n1557_));
  OR3        m1529(.A(mai_mai_n1557_), .B(mai_mai_n1555_), .C(mai_mai_n1083_), .Y(mai_mai_n1558_));
  NO3        m1530(.A(mai_mai_n1374_), .B(mai_mai_n92_), .C(k), .Y(mai_mai_n1559_));
  AOI210     m1531(.A0(mai_mai_n1559_), .A1(mai_mai_n1076_), .B0(mai_mai_n1207_), .Y(mai_mai_n1560_));
  NA2        m1532(.A(mai_mai_n1560_), .B(mai_mai_n1231_), .Y(mai_mai_n1561_));
  NO4        m1533(.A(mai_mai_n1561_), .B(mai_mai_n1558_), .C(mai_mai_n1091_), .D(mai_mai_n1070_), .Y(mai_mai_n1562_));
  NA4        m1534(.A(mai_mai_n1562_), .B(mai_mai_n1146_), .C(mai_mai_n1131_), .D(mai_mai_n1121_), .Y(mai05));
  INV        m1535(.A(m), .Y(mai_mai_n1566_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(u), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(u), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(u), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(u), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(u), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(u), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(u), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(u), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(u), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(u), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(u), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NO2        u0066(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u0067(.A(m), .B(l), .Y(men_men_n96_));
  NAi31      u0068(.An(k), .B(j), .C(u), .Y(men_men_n97_));
  NO3        u0069(.A(men_men_n97_), .B(men_men_n96_), .C(f), .Y(men_men_n98_));
  AN2        u0070(.A(j), .B(u), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(l), .C(i), .Y(men_men_n100_));
  NOi21      u0072(.An(u), .B(i), .Y(men_men_n101_));
  NOi32      u0073(.An(m), .Bn(j), .C(k), .Y(men_men_n102_));
  AOI220     u0074(.A0(men_men_n102_), .A1(men_men_n101_), .B0(men_men_n100_), .B1(men_men_n99_), .Y(men_men_n103_));
  NO2        u0075(.A(men_men_n103_), .B(f), .Y(men_men_n104_));
  NO4        u0076(.A(men_men_n104_), .B(men_men_n98_), .C(men_men_n95_), .D(men_men_n92_), .Y(men_men_n105_));
  NAi41      u0077(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n106_));
  AN2        u0078(.A(e), .B(b), .Y(men_men_n107_));
  NOi31      u0079(.An(c), .B(h), .C(f), .Y(men_men_n108_));
  NA2        u0080(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NO3        u0081(.A(men_men_n109_), .B(men_men_n106_), .C(u), .Y(men_men_n110_));
  NOi21      u0082(.An(u), .B(f), .Y(men_men_n111_));
  NOi21      u0083(.An(i), .B(h), .Y(men_men_n112_));
  NA3        u0084(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n36_), .Y(men_men_n113_));
  INV        u0085(.A(a), .Y(men_men_n114_));
  NA2        u0086(.A(men_men_n107_), .B(men_men_n114_), .Y(men_men_n115_));
  INV        u0087(.A(l), .Y(men_men_n116_));
  NOi21      u0088(.An(m), .B(n), .Y(men_men_n117_));
  AN2        u0089(.A(k), .B(h), .Y(men_men_n118_));
  NO2        u0090(.A(men_men_n113_), .B(men_men_n88_), .Y(men_men_n119_));
  INV        u0091(.A(b), .Y(men_men_n120_));
  NA2        u0092(.A(l), .B(j), .Y(men_men_n121_));
  AN2        u0093(.A(k), .B(i), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n121_), .Y(men_men_n123_));
  NA2        u0095(.A(u), .B(e), .Y(men_men_n124_));
  NOi32      u0096(.An(c), .Bn(a), .C(d), .Y(men_men_n125_));
  NA2        u0097(.A(men_men_n125_), .B(men_men_n117_), .Y(men_men_n126_));
  NO4        u0098(.A(men_men_n126_), .B(men_men_n124_), .C(men_men_n123_), .D(men_men_n120_), .Y(men_men_n127_));
  NO3        u0099(.A(men_men_n127_), .B(men_men_n119_), .C(men_men_n110_), .Y(men_men_n128_));
  OAI210     u0100(.A0(men_men_n105_), .A1(men_men_n88_), .B0(men_men_n128_), .Y(men_men_n129_));
  NOi31      u0101(.An(k), .B(m), .C(j), .Y(men_men_n130_));
  NA3        u0102(.A(men_men_n130_), .B(men_men_n79_), .C(men_men_n78_), .Y(men_men_n131_));
  NOi31      u0103(.An(k), .B(m), .C(i), .Y(men_men_n132_));
  NA3        u0104(.A(men_men_n132_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n133_));
  NA2        u0105(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n134_));
  NOi32      u0106(.An(f), .Bn(b), .C(e), .Y(men_men_n135_));
  NAi21      u0107(.An(u), .B(h), .Y(men_men_n136_));
  NAi21      u0108(.An(m), .B(n), .Y(men_men_n137_));
  NAi21      u0109(.An(j), .B(k), .Y(men_men_n138_));
  NAi41      u0110(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n139_));
  NAi31      u0111(.An(j), .B(k), .C(h), .Y(men_men_n140_));
  NO3        u0112(.A(men_men_n140_), .B(men_men_n139_), .C(men_men_n137_), .Y(men_men_n141_));
  INV        u0113(.A(men_men_n141_), .Y(men_men_n142_));
  NO2        u0114(.A(k), .B(j), .Y(men_men_n143_));
  NO2        u0115(.A(men_men_n143_), .B(men_men_n137_), .Y(men_men_n144_));
  AN2        u0116(.A(k), .B(j), .Y(men_men_n145_));
  NAi21      u0117(.An(c), .B(b), .Y(men_men_n146_));
  NA2        u0118(.A(f), .B(d), .Y(men_men_n147_));
  NO4        u0119(.A(men_men_n147_), .B(men_men_n146_), .C(men_men_n145_), .D(men_men_n136_), .Y(men_men_n148_));
  NA2        u0120(.A(h), .B(c), .Y(men_men_n149_));
  NAi31      u0121(.An(f), .B(e), .C(b), .Y(men_men_n150_));
  NA2        u0122(.A(men_men_n148_), .B(men_men_n144_), .Y(men_men_n151_));
  NA2        u0123(.A(d), .B(b), .Y(men_men_n152_));
  NAi21      u0124(.An(e), .B(f), .Y(men_men_n153_));
  NO2        u0125(.A(men_men_n153_), .B(men_men_n152_), .Y(men_men_n154_));
  NA2        u0126(.A(b), .B(a), .Y(men_men_n155_));
  NAi21      u0127(.An(e), .B(u), .Y(men_men_n156_));
  NAi21      u0128(.An(c), .B(d), .Y(men_men_n157_));
  NAi31      u0129(.An(l), .B(k), .C(h), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n137_), .B(men_men_n158_), .Y(men_men_n159_));
  NA2        u0131(.A(men_men_n159_), .B(men_men_n154_), .Y(men_men_n160_));
  NAi41      u0132(.An(men_men_n134_), .B(men_men_n160_), .C(men_men_n151_), .D(men_men_n142_), .Y(men_men_n161_));
  NAi31      u0133(.An(e), .B(f), .C(b), .Y(men_men_n162_));
  NOi21      u0134(.An(u), .B(d), .Y(men_men_n163_));
  NO2        u0135(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  NOi21      u0136(.An(h), .B(i), .Y(men_men_n165_));
  NOi21      u0137(.An(k), .B(m), .Y(men_men_n166_));
  NA3        u0138(.A(men_men_n166_), .B(men_men_n165_), .C(n), .Y(men_men_n167_));
  NOi21      u0139(.An(men_men_n164_), .B(men_men_n167_), .Y(men_men_n168_));
  NOi21      u0140(.An(h), .B(u), .Y(men_men_n169_));
  NO2        u0141(.A(men_men_n147_), .B(men_men_n146_), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n169_), .Y(men_men_n171_));
  NAi31      u0143(.An(l), .B(j), .C(h), .Y(men_men_n172_));
  NO2        u0144(.A(men_men_n172_), .B(men_men_n49_), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n67_), .Y(men_men_n174_));
  NOi32      u0146(.An(n), .Bn(k), .C(m), .Y(men_men_n175_));
  NA2        u0147(.A(l), .B(i), .Y(men_men_n176_));
  NA2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  OAI210     u0149(.A0(men_men_n177_), .A1(men_men_n171_), .B0(men_men_n174_), .Y(men_men_n178_));
  NAi31      u0150(.An(d), .B(f), .C(c), .Y(men_men_n179_));
  NAi31      u0151(.An(e), .B(f), .C(c), .Y(men_men_n180_));
  NA2        u0152(.A(men_men_n180_), .B(men_men_n179_), .Y(men_men_n181_));
  NA2        u0153(.A(j), .B(h), .Y(men_men_n182_));
  OR3        u0154(.A(n), .B(m), .C(k), .Y(men_men_n183_));
  NO2        u0155(.A(men_men_n183_), .B(men_men_n182_), .Y(men_men_n184_));
  NAi32      u0156(.An(m), .Bn(k), .C(n), .Y(men_men_n185_));
  NO2        u0157(.A(men_men_n185_), .B(men_men_n182_), .Y(men_men_n186_));
  AOI220     u0158(.A0(men_men_n186_), .A1(men_men_n164_), .B0(men_men_n184_), .B1(men_men_n181_), .Y(men_men_n187_));
  NO2        u0159(.A(n), .B(m), .Y(men_men_n188_));
  NA2        u0160(.A(men_men_n188_), .B(men_men_n50_), .Y(men_men_n189_));
  NAi21      u0161(.An(f), .B(e), .Y(men_men_n190_));
  NA2        u0162(.A(d), .B(c), .Y(men_men_n191_));
  NO2        u0163(.A(men_men_n191_), .B(men_men_n190_), .Y(men_men_n192_));
  NOi21      u0164(.An(men_men_n192_), .B(men_men_n189_), .Y(men_men_n193_));
  NAi21      u0165(.An(d), .B(c), .Y(men_men_n194_));
  NAi31      u0166(.An(m), .B(n), .C(b), .Y(men_men_n195_));
  NA2        u0167(.A(k), .B(i), .Y(men_men_n196_));
  NAi21      u0168(.An(h), .B(f), .Y(men_men_n197_));
  NO2        u0169(.A(men_men_n197_), .B(men_men_n196_), .Y(men_men_n198_));
  NO2        u0170(.A(men_men_n195_), .B(men_men_n157_), .Y(men_men_n199_));
  NA2        u0171(.A(men_men_n199_), .B(men_men_n198_), .Y(men_men_n200_));
  NOi32      u0172(.An(f), .Bn(c), .C(d), .Y(men_men_n201_));
  NOi32      u0173(.An(f), .Bn(c), .C(e), .Y(men_men_n202_));
  NO2        u0174(.A(men_men_n202_), .B(men_men_n201_), .Y(men_men_n203_));
  NO3        u0175(.A(n), .B(m), .C(j), .Y(men_men_n204_));
  NA2        u0176(.A(men_men_n204_), .B(men_men_n118_), .Y(men_men_n205_));
  AO210      u0177(.A0(men_men_n205_), .A1(men_men_n189_), .B0(men_men_n203_), .Y(men_men_n206_));
  NAi41      u0178(.An(men_men_n193_), .B(men_men_n206_), .C(men_men_n200_), .D(men_men_n187_), .Y(men_men_n207_));
  OR4        u0179(.A(men_men_n207_), .B(men_men_n178_), .C(men_men_n168_), .D(men_men_n161_), .Y(men_men_n208_));
  NO4        u0180(.A(men_men_n208_), .B(men_men_n129_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n209_));
  NA3        u0181(.A(m), .B(men_men_n116_), .C(j), .Y(men_men_n210_));
  NAi31      u0182(.An(n), .B(h), .C(u), .Y(men_men_n211_));
  NO2        u0183(.A(men_men_n211_), .B(men_men_n210_), .Y(men_men_n212_));
  NOi32      u0184(.An(m), .Bn(k), .C(l), .Y(men_men_n213_));
  NA3        u0185(.A(men_men_n213_), .B(men_men_n89_), .C(u), .Y(men_men_n214_));
  NO2        u0186(.A(men_men_n214_), .B(n), .Y(men_men_n215_));
  NOi21      u0187(.An(k), .B(j), .Y(men_men_n216_));
  NA4        u0188(.A(men_men_n216_), .B(men_men_n117_), .C(i), .D(u), .Y(men_men_n217_));
  AN2        u0189(.A(i), .B(u), .Y(men_men_n218_));
  NA3        u0190(.A(men_men_n76_), .B(men_men_n218_), .C(men_men_n117_), .Y(men_men_n219_));
  NA2        u0191(.A(men_men_n219_), .B(men_men_n217_), .Y(men_men_n220_));
  NO3        u0192(.A(men_men_n220_), .B(men_men_n215_), .C(men_men_n212_), .Y(men_men_n221_));
  NAi41      u0193(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n222_));
  INV        u0194(.A(men_men_n222_), .Y(men_men_n223_));
  INV        u0195(.A(f), .Y(men_men_n224_));
  INV        u0196(.A(u), .Y(men_men_n225_));
  NOi31      u0197(.An(i), .B(j), .C(h), .Y(men_men_n226_));
  NOi21      u0198(.An(l), .B(m), .Y(men_men_n227_));
  NA2        u0199(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n228_));
  NO3        u0200(.A(men_men_n228_), .B(men_men_n225_), .C(men_men_n224_), .Y(men_men_n229_));
  NA2        u0201(.A(men_men_n229_), .B(men_men_n223_), .Y(men_men_n230_));
  OAI210     u0202(.A0(men_men_n221_), .A1(men_men_n32_), .B0(men_men_n230_), .Y(men_men_n231_));
  NOi21      u0203(.An(n), .B(m), .Y(men_men_n232_));
  NOi32      u0204(.An(l), .Bn(i), .C(j), .Y(men_men_n233_));
  NA2        u0205(.A(men_men_n233_), .B(men_men_n232_), .Y(men_men_n234_));
  OA220      u0206(.A0(men_men_n234_), .A1(men_men_n109_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n235_));
  NAi21      u0207(.An(j), .B(h), .Y(men_men_n236_));
  XN2        u0208(.A(i), .B(h), .Y(men_men_n237_));
  NA2        u0209(.A(men_men_n237_), .B(men_men_n236_), .Y(men_men_n238_));
  NOi31      u0210(.An(k), .B(n), .C(m), .Y(men_men_n239_));
  NOi31      u0211(.An(men_men_n239_), .B(men_men_n191_), .C(men_men_n190_), .Y(men_men_n240_));
  NA2        u0212(.A(men_men_n240_), .B(men_men_n238_), .Y(men_men_n241_));
  NAi31      u0213(.An(f), .B(e), .C(c), .Y(men_men_n242_));
  NO4        u0214(.A(men_men_n242_), .B(men_men_n183_), .C(men_men_n182_), .D(men_men_n59_), .Y(men_men_n243_));
  NA4        u0215(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n244_));
  NAi32      u0216(.An(m), .Bn(i), .C(k), .Y(men_men_n245_));
  NO3        u0217(.A(men_men_n245_), .B(men_men_n93_), .C(men_men_n244_), .Y(men_men_n246_));
  NA2        u0218(.A(k), .B(h), .Y(men_men_n247_));
  NO2        u0219(.A(men_men_n246_), .B(men_men_n243_), .Y(men_men_n248_));
  NAi21      u0220(.An(n), .B(a), .Y(men_men_n249_));
  NO2        u0221(.A(men_men_n249_), .B(men_men_n152_), .Y(men_men_n250_));
  NAi41      u0222(.An(u), .B(m), .C(k), .D(h), .Y(men_men_n251_));
  NO2        u0223(.A(men_men_n251_), .B(e), .Y(men_men_n252_));
  NO3        u0224(.A(men_men_n153_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n253_));
  OAI210     u0225(.A0(men_men_n253_), .A1(men_men_n252_), .B0(men_men_n250_), .Y(men_men_n254_));
  AN4        u0226(.A(men_men_n254_), .B(men_men_n248_), .C(men_men_n241_), .D(men_men_n235_), .Y(men_men_n255_));
  OR2        u0227(.A(h), .B(u), .Y(men_men_n256_));
  NO2        u0228(.A(men_men_n256_), .B(men_men_n106_), .Y(men_men_n257_));
  NA2        u0229(.A(men_men_n257_), .B(men_men_n135_), .Y(men_men_n258_));
  NAi41      u0230(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n259_), .B(men_men_n224_), .Y(men_men_n260_));
  NA2        u0232(.A(men_men_n166_), .B(men_men_n112_), .Y(men_men_n261_));
  NAi21      u0233(.An(men_men_n261_), .B(men_men_n260_), .Y(men_men_n262_));
  NO2        u0234(.A(n), .B(a), .Y(men_men_n263_));
  NAi31      u0235(.An(men_men_n251_), .B(men_men_n263_), .C(men_men_n107_), .Y(men_men_n264_));
  AN2        u0236(.A(men_men_n264_), .B(men_men_n262_), .Y(men_men_n265_));
  NAi21      u0237(.An(h), .B(i), .Y(men_men_n266_));
  NA2        u0238(.A(men_men_n188_), .B(k), .Y(men_men_n267_));
  NO2        u0239(.A(men_men_n267_), .B(men_men_n266_), .Y(men_men_n268_));
  NA2        u0240(.A(men_men_n268_), .B(men_men_n201_), .Y(men_men_n269_));
  NA3        u0241(.A(men_men_n269_), .B(men_men_n265_), .C(men_men_n258_), .Y(men_men_n270_));
  NOi21      u0242(.An(u), .B(e), .Y(men_men_n271_));
  NO2        u0243(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n272_));
  NA2        u0244(.A(men_men_n272_), .B(men_men_n271_), .Y(men_men_n273_));
  NOi32      u0245(.An(l), .Bn(j), .C(i), .Y(men_men_n274_));
  AOI210     u0246(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n274_), .Y(men_men_n275_));
  NO2        u0247(.A(men_men_n266_), .B(men_men_n44_), .Y(men_men_n276_));
  NAi21      u0248(.An(f), .B(u), .Y(men_men_n277_));
  NO2        u0249(.A(men_men_n277_), .B(men_men_n65_), .Y(men_men_n278_));
  NO2        u0250(.A(men_men_n69_), .B(men_men_n121_), .Y(men_men_n279_));
  AOI220     u0251(.A0(men_men_n279_), .A1(men_men_n278_), .B0(men_men_n276_), .B1(men_men_n67_), .Y(men_men_n280_));
  OAI210     u0252(.A0(men_men_n275_), .A1(men_men_n273_), .B0(men_men_n280_), .Y(men_men_n281_));
  NO3        u0253(.A(men_men_n138_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n282_));
  NOi41      u0254(.An(men_men_n255_), .B(men_men_n281_), .C(men_men_n270_), .D(men_men_n231_), .Y(men_men_n283_));
  NO4        u0255(.A(men_men_n212_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n284_));
  NO2        u0256(.A(men_men_n284_), .B(men_men_n115_), .Y(men_men_n285_));
  NA3        u0257(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n286_));
  NAi21      u0258(.An(h), .B(u), .Y(men_men_n287_));
  OR4        u0259(.A(men_men_n287_), .B(men_men_n286_), .C(men_men_n234_), .D(e), .Y(men_men_n288_));
  NO2        u0260(.A(men_men_n261_), .B(men_men_n277_), .Y(men_men_n289_));
  NA2        u0261(.A(men_men_n289_), .B(men_men_n78_), .Y(men_men_n290_));
  NAi31      u0262(.An(u), .B(k), .C(h), .Y(men_men_n291_));
  NO3        u0263(.A(men_men_n137_), .B(men_men_n291_), .C(l), .Y(men_men_n292_));
  NAi31      u0264(.An(e), .B(d), .C(a), .Y(men_men_n293_));
  NA2        u0265(.A(men_men_n292_), .B(men_men_n135_), .Y(men_men_n294_));
  NA3        u0266(.A(men_men_n294_), .B(men_men_n290_), .C(men_men_n288_), .Y(men_men_n295_));
  NA3        u0267(.A(men_men_n166_), .B(men_men_n165_), .C(men_men_n86_), .Y(men_men_n296_));
  NO2        u0268(.A(men_men_n296_), .B(men_men_n203_), .Y(men_men_n297_));
  INV        u0269(.A(men_men_n297_), .Y(men_men_n298_));
  NA3        u0270(.A(e), .B(c), .C(b), .Y(men_men_n299_));
  NO2        u0271(.A(men_men_n60_), .B(men_men_n299_), .Y(men_men_n300_));
  NAi32      u0272(.An(k), .Bn(i), .C(j), .Y(men_men_n301_));
  NAi31      u0273(.An(h), .B(l), .C(i), .Y(men_men_n302_));
  NA3        u0274(.A(men_men_n302_), .B(men_men_n301_), .C(men_men_n172_), .Y(men_men_n303_));
  NOi21      u0275(.An(men_men_n303_), .B(men_men_n49_), .Y(men_men_n304_));
  OAI210     u0276(.A0(men_men_n278_), .A1(men_men_n300_), .B0(men_men_n304_), .Y(men_men_n305_));
  NAi21      u0277(.An(l), .B(k), .Y(men_men_n306_));
  NO2        u0278(.A(men_men_n306_), .B(men_men_n49_), .Y(men_men_n307_));
  NOi21      u0279(.An(l), .B(j), .Y(men_men_n308_));
  NA2        u0280(.A(men_men_n169_), .B(men_men_n308_), .Y(men_men_n309_));
  NAi32      u0281(.An(j), .Bn(h), .C(i), .Y(men_men_n310_));
  NAi21      u0282(.An(m), .B(l), .Y(men_men_n311_));
  NO3        u0283(.A(men_men_n311_), .B(men_men_n310_), .C(men_men_n86_), .Y(men_men_n312_));
  NA2        u0284(.A(h), .B(u), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n175_), .B(men_men_n45_), .Y(men_men_n314_));
  NO2        u0286(.A(men_men_n314_), .B(men_men_n313_), .Y(men_men_n315_));
  OAI210     u0287(.A0(men_men_n315_), .A1(men_men_n312_), .B0(men_men_n170_), .Y(men_men_n316_));
  NA3        u0288(.A(men_men_n316_), .B(men_men_n305_), .C(men_men_n298_), .Y(men_men_n317_));
  NO2        u0289(.A(men_men_n150_), .B(d), .Y(men_men_n318_));
  NA2        u0290(.A(men_men_n318_), .B(men_men_n53_), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n109_), .B(men_men_n106_), .Y(men_men_n320_));
  NAi32      u0292(.An(n), .Bn(m), .C(l), .Y(men_men_n321_));
  NO2        u0293(.A(men_men_n321_), .B(men_men_n310_), .Y(men_men_n322_));
  NA2        u0294(.A(men_men_n322_), .B(men_men_n192_), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n126_), .B(men_men_n120_), .Y(men_men_n324_));
  NAi31      u0296(.An(k), .B(l), .C(j), .Y(men_men_n325_));
  OAI210     u0297(.A0(men_men_n306_), .A1(j), .B0(men_men_n325_), .Y(men_men_n326_));
  NOi21      u0298(.An(men_men_n326_), .B(men_men_n124_), .Y(men_men_n327_));
  NA2        u0299(.A(men_men_n327_), .B(men_men_n324_), .Y(men_men_n328_));
  NA3        u0300(.A(men_men_n328_), .B(men_men_n323_), .C(men_men_n319_), .Y(men_men_n329_));
  NO4        u0301(.A(men_men_n329_), .B(men_men_n317_), .C(men_men_n295_), .D(men_men_n285_), .Y(men_men_n330_));
  NA2        u0302(.A(men_men_n268_), .B(men_men_n202_), .Y(men_men_n331_));
  NAi21      u0303(.An(m), .B(k), .Y(men_men_n332_));
  NO2        u0304(.A(men_men_n237_), .B(men_men_n332_), .Y(men_men_n333_));
  NAi41      u0305(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n334_));
  NO2        u0306(.A(men_men_n334_), .B(men_men_n156_), .Y(men_men_n335_));
  NA2        u0307(.A(men_men_n335_), .B(men_men_n333_), .Y(men_men_n336_));
  NAi31      u0308(.An(i), .B(l), .C(h), .Y(men_men_n337_));
  NO4        u0309(.A(men_men_n337_), .B(men_men_n156_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n338_));
  NA2        u0310(.A(e), .B(c), .Y(men_men_n339_));
  NO3        u0311(.A(men_men_n339_), .B(n), .C(d), .Y(men_men_n340_));
  NOi21      u0312(.An(f), .B(h), .Y(men_men_n341_));
  NA2        u0313(.A(men_men_n341_), .B(men_men_n122_), .Y(men_men_n342_));
  NO2        u0314(.A(men_men_n342_), .B(men_men_n225_), .Y(men_men_n343_));
  NAi31      u0315(.An(d), .B(e), .C(b), .Y(men_men_n344_));
  NO2        u0316(.A(men_men_n137_), .B(men_men_n344_), .Y(men_men_n345_));
  NA2        u0317(.A(men_men_n345_), .B(men_men_n343_), .Y(men_men_n346_));
  NAi41      u0318(.An(men_men_n338_), .B(men_men_n346_), .C(men_men_n336_), .D(men_men_n331_), .Y(men_men_n347_));
  NO4        u0319(.A(men_men_n334_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n225_), .Y(men_men_n348_));
  NA2        u0320(.A(men_men_n263_), .B(men_men_n107_), .Y(men_men_n349_));
  OR2        u0321(.A(men_men_n349_), .B(men_men_n214_), .Y(men_men_n350_));
  NOi31      u0322(.An(l), .B(n), .C(m), .Y(men_men_n351_));
  NA2        u0323(.A(men_men_n351_), .B(men_men_n226_), .Y(men_men_n352_));
  NO2        u0324(.A(men_men_n352_), .B(men_men_n203_), .Y(men_men_n353_));
  NAi32      u0325(.An(men_men_n353_), .Bn(men_men_n348_), .C(men_men_n350_), .Y(men_men_n354_));
  NAi32      u0326(.An(m), .Bn(j), .C(k), .Y(men_men_n355_));
  NAi41      u0327(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n356_));
  OAI210     u0328(.A0(men_men_n222_), .A1(men_men_n355_), .B0(men_men_n356_), .Y(men_men_n357_));
  NOi31      u0329(.An(j), .B(m), .C(k), .Y(men_men_n358_));
  NO2        u0330(.A(men_men_n130_), .B(men_men_n358_), .Y(men_men_n359_));
  AN3        u0331(.A(h), .B(u), .C(f), .Y(men_men_n360_));
  NAi31      u0332(.An(men_men_n359_), .B(men_men_n360_), .C(men_men_n357_), .Y(men_men_n361_));
  NOi32      u0333(.An(m), .Bn(j), .C(l), .Y(men_men_n362_));
  NO2        u0334(.A(men_men_n362_), .B(men_men_n100_), .Y(men_men_n363_));
  NAi32      u0335(.An(men_men_n363_), .Bn(men_men_n211_), .C(men_men_n318_), .Y(men_men_n364_));
  NO2        u0336(.A(men_men_n311_), .B(men_men_n310_), .Y(men_men_n365_));
  NO2        u0337(.A(men_men_n228_), .B(u), .Y(men_men_n366_));
  NA2        u0338(.A(men_men_n260_), .B(men_men_n365_), .Y(men_men_n367_));
  NA2        u0339(.A(men_men_n245_), .B(men_men_n81_), .Y(men_men_n368_));
  NA3        u0340(.A(men_men_n368_), .B(men_men_n360_), .C(men_men_n223_), .Y(men_men_n369_));
  NA4        u0341(.A(men_men_n369_), .B(men_men_n367_), .C(men_men_n364_), .D(men_men_n361_), .Y(men_men_n370_));
  NA3        u0342(.A(h), .B(u), .C(f), .Y(men_men_n371_));
  NO2        u0343(.A(men_men_n371_), .B(men_men_n77_), .Y(men_men_n372_));
  INV        u0344(.A(men_men_n222_), .Y(men_men_n373_));
  NA2        u0345(.A(men_men_n169_), .B(e), .Y(men_men_n374_));
  NO2        u0346(.A(men_men_n374_), .B(men_men_n41_), .Y(men_men_n375_));
  AOI220     u0347(.A0(men_men_n375_), .A1(men_men_n324_), .B0(men_men_n373_), .B1(men_men_n372_), .Y(men_men_n376_));
  NOi32      u0348(.An(j), .Bn(u), .C(i), .Y(men_men_n377_));
  NA3        u0349(.A(men_men_n377_), .B(men_men_n306_), .C(men_men_n117_), .Y(men_men_n378_));
  AO210      u0350(.A0(men_men_n115_), .A1(men_men_n32_), .B0(men_men_n378_), .Y(men_men_n379_));
  NOi32      u0351(.An(e), .Bn(b), .C(a), .Y(men_men_n380_));
  AN2        u0352(.A(l), .B(j), .Y(men_men_n381_));
  NO2        u0353(.A(men_men_n332_), .B(men_men_n381_), .Y(men_men_n382_));
  NO3        u0354(.A(men_men_n334_), .B(men_men_n72_), .C(men_men_n225_), .Y(men_men_n383_));
  NA3        u0355(.A(men_men_n219_), .B(men_men_n217_), .C(men_men_n35_), .Y(men_men_n384_));
  AOI220     u0356(.A0(men_men_n384_), .A1(men_men_n380_), .B0(men_men_n383_), .B1(men_men_n382_), .Y(men_men_n385_));
  NO2        u0357(.A(men_men_n344_), .B(n), .Y(men_men_n386_));
  NA2        u0358(.A(men_men_n218_), .B(k), .Y(men_men_n387_));
  NA3        u0359(.A(m), .B(men_men_n116_), .C(men_men_n224_), .Y(men_men_n388_));
  NA4        u0360(.A(men_men_n213_), .B(men_men_n89_), .C(u), .D(men_men_n224_), .Y(men_men_n389_));
  OAI210     u0361(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n389_), .Y(men_men_n390_));
  NAi41      u0362(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n391_));
  NA2        u0363(.A(men_men_n51_), .B(men_men_n117_), .Y(men_men_n392_));
  NO2        u0364(.A(men_men_n392_), .B(men_men_n391_), .Y(men_men_n393_));
  AOI220     u0365(.A0(men_men_n393_), .A1(b), .B0(men_men_n390_), .B1(men_men_n386_), .Y(men_men_n394_));
  NA4        u0366(.A(men_men_n394_), .B(men_men_n385_), .C(men_men_n379_), .D(men_men_n376_), .Y(men_men_n395_));
  NO4        u0367(.A(men_men_n395_), .B(men_men_n370_), .C(men_men_n354_), .D(men_men_n347_), .Y(men_men_n396_));
  NA4        u0368(.A(men_men_n396_), .B(men_men_n330_), .C(men_men_n283_), .D(men_men_n209_), .Y(men10));
  NA3        u0369(.A(m), .B(k), .C(i), .Y(men_men_n398_));
  NO3        u0370(.A(men_men_n398_), .B(j), .C(men_men_n225_), .Y(men_men_n399_));
  NOi21      u0371(.An(e), .B(f), .Y(men_men_n400_));
  NO4        u0372(.A(men_men_n157_), .B(men_men_n400_), .C(n), .D(men_men_n114_), .Y(men_men_n401_));
  NAi31      u0373(.An(b), .B(f), .C(c), .Y(men_men_n402_));
  INV        u0374(.A(men_men_n402_), .Y(men_men_n403_));
  NOi32      u0375(.An(k), .Bn(h), .C(j), .Y(men_men_n404_));
  NA2        u0376(.A(men_men_n404_), .B(men_men_n232_), .Y(men_men_n405_));
  NA2        u0377(.A(men_men_n167_), .B(men_men_n405_), .Y(men_men_n406_));
  AOI220     u0378(.A0(men_men_n406_), .A1(men_men_n403_), .B0(men_men_n401_), .B1(men_men_n399_), .Y(men_men_n407_));
  AN2        u0379(.A(j), .B(h), .Y(men_men_n408_));
  NO3        u0380(.A(n), .B(m), .C(k), .Y(men_men_n409_));
  NA2        u0381(.A(men_men_n409_), .B(men_men_n408_), .Y(men_men_n410_));
  NO3        u0382(.A(men_men_n410_), .B(men_men_n157_), .C(men_men_n224_), .Y(men_men_n411_));
  OR2        u0383(.A(m), .B(k), .Y(men_men_n412_));
  NO2        u0384(.A(men_men_n182_), .B(men_men_n412_), .Y(men_men_n413_));
  NA4        u0385(.A(n), .B(f), .C(c), .D(men_men_n120_), .Y(men_men_n414_));
  NOi21      u0386(.An(men_men_n413_), .B(men_men_n414_), .Y(men_men_n415_));
  NOi32      u0387(.An(d), .Bn(a), .C(c), .Y(men_men_n416_));
  NA2        u0388(.A(men_men_n416_), .B(men_men_n190_), .Y(men_men_n417_));
  NAi21      u0389(.An(i), .B(u), .Y(men_men_n418_));
  NAi31      u0390(.An(k), .B(m), .C(j), .Y(men_men_n419_));
  NO3        u0391(.A(men_men_n419_), .B(men_men_n418_), .C(n), .Y(men_men_n420_));
  NOi21      u0392(.An(men_men_n420_), .B(men_men_n417_), .Y(men_men_n421_));
  NO3        u0393(.A(men_men_n421_), .B(men_men_n415_), .C(men_men_n411_), .Y(men_men_n422_));
  NO2        u0394(.A(men_men_n414_), .B(men_men_n311_), .Y(men_men_n423_));
  NOi32      u0395(.An(f), .Bn(d), .C(c), .Y(men_men_n424_));
  AOI220     u0396(.A0(men_men_n424_), .A1(men_men_n322_), .B0(men_men_n423_), .B1(men_men_n226_), .Y(men_men_n425_));
  NA3        u0397(.A(men_men_n425_), .B(men_men_n422_), .C(men_men_n407_), .Y(men_men_n426_));
  NO2        u0398(.A(men_men_n59_), .B(men_men_n120_), .Y(men_men_n427_));
  NA2        u0399(.A(men_men_n263_), .B(men_men_n427_), .Y(men_men_n428_));
  INV        u0400(.A(e), .Y(men_men_n429_));
  NA2        u0401(.A(men_men_n46_), .B(e), .Y(men_men_n430_));
  OAI220     u0402(.A0(men_men_n430_), .A1(men_men_n210_), .B0(men_men_n214_), .B1(men_men_n429_), .Y(men_men_n431_));
  AN2        u0403(.A(u), .B(e), .Y(men_men_n432_));
  NA3        u0404(.A(men_men_n432_), .B(men_men_n213_), .C(i), .Y(men_men_n433_));
  OAI210     u0405(.A0(men_men_n91_), .A1(men_men_n429_), .B0(men_men_n433_), .Y(men_men_n434_));
  NO2        u0406(.A(men_men_n103_), .B(men_men_n429_), .Y(men_men_n435_));
  NO3        u0407(.A(men_men_n435_), .B(men_men_n434_), .C(men_men_n431_), .Y(men_men_n436_));
  NOi32      u0408(.An(h), .Bn(e), .C(u), .Y(men_men_n437_));
  NA3        u0409(.A(men_men_n437_), .B(men_men_n308_), .C(m), .Y(men_men_n438_));
  NOi21      u0410(.An(u), .B(h), .Y(men_men_n439_));
  AN3        u0411(.A(m), .B(l), .C(i), .Y(men_men_n440_));
  NA3        u0412(.A(men_men_n440_), .B(men_men_n439_), .C(e), .Y(men_men_n441_));
  AN3        u0413(.A(h), .B(u), .C(e), .Y(men_men_n442_));
  NA2        u0414(.A(men_men_n442_), .B(men_men_n100_), .Y(men_men_n443_));
  AN3        u0415(.A(men_men_n443_), .B(men_men_n441_), .C(men_men_n438_), .Y(men_men_n444_));
  AOI210     u0416(.A0(men_men_n444_), .A1(men_men_n436_), .B0(men_men_n428_), .Y(men_men_n445_));
  NA3        u0417(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n446_));
  NO2        u0418(.A(men_men_n446_), .B(men_men_n428_), .Y(men_men_n447_));
  NAi31      u0419(.An(b), .B(c), .C(a), .Y(men_men_n448_));
  NO2        u0420(.A(men_men_n448_), .B(n), .Y(men_men_n449_));
  OAI210     u0421(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n450_));
  NO2        u0422(.A(men_men_n450_), .B(men_men_n153_), .Y(men_men_n451_));
  NA2        u0423(.A(men_men_n451_), .B(men_men_n449_), .Y(men_men_n452_));
  INV        u0424(.A(men_men_n452_), .Y(men_men_n453_));
  NO4        u0425(.A(men_men_n453_), .B(men_men_n447_), .C(men_men_n445_), .D(men_men_n426_), .Y(men_men_n454_));
  NA2        u0426(.A(i), .B(u), .Y(men_men_n455_));
  NO3        u0427(.A(men_men_n293_), .B(men_men_n455_), .C(c), .Y(men_men_n456_));
  NOi21      u0428(.An(a), .B(n), .Y(men_men_n457_));
  NOi21      u0429(.An(d), .B(c), .Y(men_men_n458_));
  NA2        u0430(.A(men_men_n458_), .B(men_men_n457_), .Y(men_men_n459_));
  NA3        u0431(.A(i), .B(u), .C(f), .Y(men_men_n460_));
  NA2        u0432(.A(men_men_n456_), .B(men_men_n307_), .Y(men_men_n461_));
  OR2        u0433(.A(n), .B(m), .Y(men_men_n462_));
  NO2        u0434(.A(men_men_n462_), .B(men_men_n158_), .Y(men_men_n463_));
  NO2        u0435(.A(men_men_n191_), .B(men_men_n153_), .Y(men_men_n464_));
  OAI210     u0436(.A0(men_men_n463_), .A1(men_men_n184_), .B0(men_men_n464_), .Y(men_men_n465_));
  INV        u0437(.A(men_men_n392_), .Y(men_men_n466_));
  NA3        u0438(.A(men_men_n466_), .B(men_men_n380_), .C(d), .Y(men_men_n467_));
  NO2        u0439(.A(men_men_n448_), .B(men_men_n49_), .Y(men_men_n468_));
  NO3        u0440(.A(men_men_n66_), .B(men_men_n116_), .C(e), .Y(men_men_n469_));
  NAi21      u0441(.An(k), .B(j), .Y(men_men_n470_));
  NA2        u0442(.A(men_men_n266_), .B(men_men_n470_), .Y(men_men_n471_));
  NA3        u0443(.A(men_men_n471_), .B(men_men_n469_), .C(men_men_n468_), .Y(men_men_n472_));
  NAi21      u0444(.An(e), .B(d), .Y(men_men_n473_));
  NO2        u0445(.A(men_men_n473_), .B(men_men_n56_), .Y(men_men_n474_));
  NO2        u0446(.A(men_men_n267_), .B(men_men_n224_), .Y(men_men_n475_));
  NA3        u0447(.A(men_men_n475_), .B(men_men_n474_), .C(men_men_n238_), .Y(men_men_n476_));
  NA4        u0448(.A(men_men_n476_), .B(men_men_n472_), .C(men_men_n467_), .D(men_men_n465_), .Y(men_men_n477_));
  NO2        u0449(.A(men_men_n352_), .B(men_men_n224_), .Y(men_men_n478_));
  NA2        u0450(.A(men_men_n478_), .B(men_men_n474_), .Y(men_men_n479_));
  NOi31      u0451(.An(n), .B(m), .C(k), .Y(men_men_n480_));
  AOI220     u0452(.A0(men_men_n480_), .A1(men_men_n408_), .B0(men_men_n232_), .B1(men_men_n50_), .Y(men_men_n481_));
  NAi31      u0453(.An(u), .B(f), .C(c), .Y(men_men_n482_));
  OR3        u0454(.A(men_men_n482_), .B(men_men_n481_), .C(e), .Y(men_men_n483_));
  NA3        u0455(.A(men_men_n483_), .B(men_men_n479_), .C(men_men_n323_), .Y(men_men_n484_));
  NOi41      u0456(.An(men_men_n461_), .B(men_men_n484_), .C(men_men_n477_), .D(men_men_n281_), .Y(men_men_n485_));
  NOi32      u0457(.An(c), .Bn(a), .C(b), .Y(men_men_n486_));
  NA2        u0458(.A(men_men_n486_), .B(men_men_n117_), .Y(men_men_n487_));
  NA2        u0459(.A(men_men_n291_), .B(men_men_n158_), .Y(men_men_n488_));
  AN2        u0460(.A(e), .B(d), .Y(men_men_n489_));
  NA2        u0461(.A(men_men_n489_), .B(men_men_n488_), .Y(men_men_n490_));
  INV        u0462(.A(men_men_n153_), .Y(men_men_n491_));
  NO2        u0463(.A(men_men_n136_), .B(men_men_n41_), .Y(men_men_n492_));
  NO2        u0464(.A(men_men_n66_), .B(e), .Y(men_men_n493_));
  NA4        u0465(.A(men_men_n337_), .B(men_men_n172_), .C(men_men_n275_), .D(men_men_n123_), .Y(men_men_n494_));
  NA2        u0466(.A(men_men_n494_), .B(men_men_n493_), .Y(men_men_n495_));
  AOI210     u0467(.A0(men_men_n495_), .A1(men_men_n490_), .B0(men_men_n487_), .Y(men_men_n496_));
  NO2        u0468(.A(men_men_n220_), .B(men_men_n215_), .Y(men_men_n497_));
  NOi21      u0469(.An(a), .B(b), .Y(men_men_n498_));
  NA3        u0470(.A(e), .B(d), .C(c), .Y(men_men_n499_));
  NAi21      u0471(.An(men_men_n499_), .B(men_men_n498_), .Y(men_men_n500_));
  AOI210     u0472(.A0(men_men_n284_), .A1(men_men_n497_), .B0(men_men_n500_), .Y(men_men_n501_));
  NO4        u0473(.A(men_men_n197_), .B(men_men_n106_), .C(men_men_n56_), .D(b), .Y(men_men_n502_));
  NA2        u0474(.A(men_men_n403_), .B(men_men_n159_), .Y(men_men_n503_));
  OR2        u0475(.A(k), .B(j), .Y(men_men_n504_));
  NA2        u0476(.A(l), .B(k), .Y(men_men_n505_));
  NA3        u0477(.A(men_men_n505_), .B(men_men_n504_), .C(men_men_n232_), .Y(men_men_n506_));
  AOI210     u0478(.A0(men_men_n245_), .A1(men_men_n355_), .B0(men_men_n86_), .Y(men_men_n507_));
  NOi21      u0479(.An(men_men_n506_), .B(men_men_n507_), .Y(men_men_n508_));
  OR3        u0480(.A(men_men_n508_), .B(men_men_n149_), .C(men_men_n139_), .Y(men_men_n509_));
  NA2        u0481(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n510_));
  NA2        u0482(.A(men_men_n416_), .B(men_men_n117_), .Y(men_men_n511_));
  NO4        u0483(.A(men_men_n511_), .B(men_men_n97_), .C(men_men_n116_), .D(e), .Y(men_men_n512_));
  NO3        u0484(.A(men_men_n512_), .B(men_men_n510_), .C(men_men_n338_), .Y(men_men_n513_));
  NA3        u0485(.A(men_men_n513_), .B(men_men_n509_), .C(men_men_n503_), .Y(men_men_n514_));
  NO4        u0486(.A(men_men_n514_), .B(men_men_n502_), .C(men_men_n501_), .D(men_men_n496_), .Y(men_men_n515_));
  NA2        u0487(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n516_));
  NOi21      u0488(.An(d), .B(e), .Y(men_men_n517_));
  NO2        u0489(.A(men_men_n197_), .B(men_men_n56_), .Y(men_men_n518_));
  NAi31      u0490(.An(j), .B(l), .C(i), .Y(men_men_n519_));
  OAI210     u0491(.A0(men_men_n519_), .A1(men_men_n137_), .B0(men_men_n106_), .Y(men_men_n520_));
  NA4        u0492(.A(men_men_n520_), .B(men_men_n518_), .C(men_men_n517_), .D(b), .Y(men_men_n521_));
  NO3        u0493(.A(men_men_n417_), .B(men_men_n363_), .C(men_men_n211_), .Y(men_men_n522_));
  NO2        u0494(.A(men_men_n417_), .B(men_men_n392_), .Y(men_men_n523_));
  NO4        u0495(.A(men_men_n523_), .B(men_men_n522_), .C(men_men_n193_), .D(men_men_n320_), .Y(men_men_n524_));
  NA4        u0496(.A(men_men_n524_), .B(men_men_n521_), .C(men_men_n516_), .D(men_men_n255_), .Y(men_men_n525_));
  OAI210     u0497(.A0(men_men_n132_), .A1(men_men_n130_), .B0(n), .Y(men_men_n526_));
  NO2        u0498(.A(men_men_n526_), .B(men_men_n136_), .Y(men_men_n527_));
  AO210      u0499(.A0(men_men_n312_), .A1(men_men_n225_), .B0(men_men_n257_), .Y(men_men_n528_));
  OA210      u0500(.A0(men_men_n528_), .A1(men_men_n527_), .B0(men_men_n202_), .Y(men_men_n529_));
  XO2        u0501(.A(i), .B(h), .Y(men_men_n530_));
  NA3        u0502(.A(men_men_n530_), .B(men_men_n166_), .C(n), .Y(men_men_n531_));
  NAi41      u0503(.An(men_men_n312_), .B(men_men_n531_), .C(men_men_n481_), .D(men_men_n405_), .Y(men_men_n532_));
  NOi32      u0504(.An(men_men_n532_), .Bn(men_men_n493_), .C(men_men_n286_), .Y(men_men_n533_));
  NAi31      u0505(.An(c), .B(f), .C(d), .Y(men_men_n534_));
  AOI210     u0506(.A0(men_men_n296_), .A1(men_men_n205_), .B0(men_men_n534_), .Y(men_men_n535_));
  NOi21      u0507(.An(men_men_n84_), .B(men_men_n535_), .Y(men_men_n536_));
  NA3        u0508(.A(men_men_n401_), .B(men_men_n100_), .C(men_men_n99_), .Y(men_men_n537_));
  NA2        u0509(.A(men_men_n239_), .B(men_men_n112_), .Y(men_men_n538_));
  AOI210     u0510(.A0(men_men_n538_), .A1(men_men_n189_), .B0(men_men_n534_), .Y(men_men_n539_));
  NOi21      u0511(.An(men_men_n537_), .B(men_men_n539_), .Y(men_men_n540_));
  AO220      u0512(.A0(men_men_n304_), .A1(men_men_n278_), .B0(men_men_n173_), .B1(men_men_n67_), .Y(men_men_n541_));
  NA3        u0513(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n542_));
  NO2        u0514(.A(men_men_n542_), .B(men_men_n459_), .Y(men_men_n543_));
  INV        u0515(.A(men_men_n543_), .Y(men_men_n544_));
  NAi41      u0516(.An(men_men_n541_), .B(men_men_n544_), .C(men_men_n540_), .D(men_men_n536_), .Y(men_men_n545_));
  NO4        u0517(.A(men_men_n545_), .B(men_men_n533_), .C(men_men_n529_), .D(men_men_n525_), .Y(men_men_n546_));
  NA4        u0518(.A(men_men_n546_), .B(men_men_n515_), .C(men_men_n485_), .D(men_men_n454_), .Y(men11));
  NO2        u0519(.A(men_men_n73_), .B(f), .Y(men_men_n548_));
  NA2        u0520(.A(j), .B(u), .Y(men_men_n549_));
  NAi31      u0521(.An(i), .B(m), .C(l), .Y(men_men_n550_));
  NA3        u0522(.A(m), .B(k), .C(j), .Y(men_men_n551_));
  OAI220     u0523(.A0(men_men_n551_), .A1(men_men_n136_), .B0(men_men_n550_), .B1(men_men_n549_), .Y(men_men_n552_));
  NOi32      u0524(.An(e), .Bn(b), .C(f), .Y(men_men_n553_));
  NA2        u0525(.A(men_men_n274_), .B(men_men_n117_), .Y(men_men_n554_));
  NA2        u0526(.A(men_men_n46_), .B(j), .Y(men_men_n555_));
  OAI220     u0527(.A0(men_men_n555_), .A1(men_men_n314_), .B0(men_men_n554_), .B1(men_men_n225_), .Y(men_men_n556_));
  NAi31      u0528(.An(d), .B(e), .C(a), .Y(men_men_n557_));
  NO2        u0529(.A(men_men_n557_), .B(n), .Y(men_men_n558_));
  AOI220     u0530(.A0(men_men_n558_), .A1(men_men_n104_), .B0(men_men_n556_), .B1(men_men_n553_), .Y(men_men_n559_));
  NAi41      u0531(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n560_));
  AN2        u0532(.A(men_men_n560_), .B(men_men_n391_), .Y(men_men_n561_));
  AOI210     u0533(.A0(men_men_n561_), .A1(men_men_n417_), .B0(men_men_n287_), .Y(men_men_n562_));
  NA2        u0534(.A(j), .B(i), .Y(men_men_n563_));
  NAi31      u0535(.An(n), .B(m), .C(k), .Y(men_men_n564_));
  NO3        u0536(.A(men_men_n564_), .B(men_men_n563_), .C(men_men_n116_), .Y(men_men_n565_));
  NO4        u0537(.A(n), .B(d), .C(men_men_n120_), .D(a), .Y(men_men_n566_));
  OR2        u0538(.A(n), .B(c), .Y(men_men_n567_));
  NO2        u0539(.A(men_men_n567_), .B(men_men_n155_), .Y(men_men_n568_));
  NO2        u0540(.A(men_men_n568_), .B(men_men_n566_), .Y(men_men_n569_));
  NOi32      u0541(.An(u), .Bn(f), .C(i), .Y(men_men_n570_));
  NA2        u0542(.A(men_men_n552_), .B(f), .Y(men_men_n571_));
  NO2        u0543(.A(men_men_n291_), .B(men_men_n49_), .Y(men_men_n572_));
  NO2        u0544(.A(men_men_n571_), .B(men_men_n569_), .Y(men_men_n573_));
  AOI210     u0545(.A0(men_men_n565_), .A1(men_men_n562_), .B0(men_men_n573_), .Y(men_men_n574_));
  NA2        u0546(.A(men_men_n145_), .B(men_men_n34_), .Y(men_men_n575_));
  OAI220     u0547(.A0(men_men_n575_), .A1(m), .B0(men_men_n555_), .B1(men_men_n245_), .Y(men_men_n576_));
  NOi41      u0548(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n577_));
  NAi32      u0549(.An(e), .Bn(b), .C(c), .Y(men_men_n578_));
  OR2        u0550(.A(men_men_n578_), .B(men_men_n86_), .Y(men_men_n579_));
  AN2        u0551(.A(men_men_n356_), .B(men_men_n334_), .Y(men_men_n580_));
  NA2        u0552(.A(men_men_n580_), .B(men_men_n579_), .Y(men_men_n581_));
  OA210      u0553(.A0(men_men_n581_), .A1(men_men_n577_), .B0(men_men_n576_), .Y(men_men_n582_));
  OAI220     u0554(.A0(men_men_n419_), .A1(men_men_n418_), .B0(men_men_n550_), .B1(men_men_n549_), .Y(men_men_n583_));
  NAi31      u0555(.An(d), .B(c), .C(a), .Y(men_men_n584_));
  NO2        u0556(.A(men_men_n584_), .B(n), .Y(men_men_n585_));
  NA3        u0557(.A(men_men_n585_), .B(men_men_n583_), .C(e), .Y(men_men_n586_));
  NO3        u0558(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n225_), .Y(men_men_n587_));
  NO2        u0559(.A(men_men_n242_), .B(men_men_n114_), .Y(men_men_n588_));
  OAI210     u0560(.A0(men_men_n587_), .A1(men_men_n420_), .B0(men_men_n588_), .Y(men_men_n589_));
  NA2        u0561(.A(men_men_n589_), .B(men_men_n586_), .Y(men_men_n590_));
  NO2        u0562(.A(men_men_n293_), .B(n), .Y(men_men_n591_));
  NO2        u0563(.A(men_men_n449_), .B(men_men_n591_), .Y(men_men_n592_));
  NA2        u0564(.A(men_men_n583_), .B(f), .Y(men_men_n593_));
  NAi32      u0565(.An(d), .Bn(a), .C(b), .Y(men_men_n594_));
  NA2        u0566(.A(h), .B(f), .Y(men_men_n595_));
  NO2        u0567(.A(men_men_n595_), .B(men_men_n97_), .Y(men_men_n596_));
  NO3        u0568(.A(men_men_n185_), .B(men_men_n182_), .C(u), .Y(men_men_n597_));
  NA2        u0569(.A(men_men_n597_), .B(men_men_n58_), .Y(men_men_n598_));
  OAI210     u0570(.A0(men_men_n593_), .A1(men_men_n592_), .B0(men_men_n598_), .Y(men_men_n599_));
  AN3        u0571(.A(j), .B(h), .C(u), .Y(men_men_n600_));
  NO2        u0572(.A(men_men_n152_), .B(c), .Y(men_men_n601_));
  NA3        u0573(.A(men_men_n601_), .B(men_men_n600_), .C(men_men_n480_), .Y(men_men_n602_));
  NA3        u0574(.A(f), .B(d), .C(b), .Y(men_men_n603_));
  NO4        u0575(.A(men_men_n603_), .B(men_men_n185_), .C(men_men_n182_), .D(u), .Y(men_men_n604_));
  NAi21      u0576(.An(men_men_n604_), .B(men_men_n602_), .Y(men_men_n605_));
  NO4        u0577(.A(men_men_n605_), .B(men_men_n599_), .C(men_men_n590_), .D(men_men_n582_), .Y(men_men_n606_));
  AN3        u0578(.A(men_men_n606_), .B(men_men_n574_), .C(men_men_n559_), .Y(men_men_n607_));
  INV        u0579(.A(k), .Y(men_men_n608_));
  NA3        u0580(.A(l), .B(men_men_n608_), .C(i), .Y(men_men_n609_));
  INV        u0581(.A(men_men_n609_), .Y(men_men_n610_));
  NA4        u0582(.A(men_men_n416_), .B(men_men_n439_), .C(men_men_n190_), .D(men_men_n117_), .Y(men_men_n611_));
  NAi32      u0583(.An(h), .Bn(f), .C(u), .Y(men_men_n612_));
  NAi41      u0584(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n613_));
  OAI210     u0585(.A0(men_men_n557_), .A1(n), .B0(men_men_n613_), .Y(men_men_n614_));
  NA2        u0586(.A(men_men_n614_), .B(m), .Y(men_men_n615_));
  NAi31      u0587(.An(h), .B(u), .C(f), .Y(men_men_n616_));
  OR3        u0588(.A(men_men_n616_), .B(men_men_n293_), .C(men_men_n49_), .Y(men_men_n617_));
  NA4        u0589(.A(men_men_n439_), .B(men_men_n125_), .C(men_men_n117_), .D(e), .Y(men_men_n618_));
  AN2        u0590(.A(men_men_n618_), .B(men_men_n617_), .Y(men_men_n619_));
  OA210      u0591(.A0(men_men_n615_), .A1(men_men_n612_), .B0(men_men_n619_), .Y(men_men_n620_));
  NA2        u0592(.A(men_men_n620_), .B(men_men_n611_), .Y(men_men_n621_));
  NAi31      u0593(.An(f), .B(h), .C(u), .Y(men_men_n622_));
  NO4        u0594(.A(men_men_n325_), .B(men_men_n622_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n623_));
  NOi32      u0595(.An(b), .Bn(a), .C(c), .Y(men_men_n624_));
  NOi41      u0596(.An(men_men_n624_), .B(men_men_n371_), .C(men_men_n69_), .D(men_men_n121_), .Y(men_men_n625_));
  OR2        u0597(.A(men_men_n625_), .B(men_men_n623_), .Y(men_men_n626_));
  NOi32      u0598(.An(d), .Bn(a), .C(e), .Y(men_men_n627_));
  NA2        u0599(.A(men_men_n627_), .B(men_men_n117_), .Y(men_men_n628_));
  NO2        u0600(.A(n), .B(c), .Y(men_men_n629_));
  NA3        u0601(.A(men_men_n629_), .B(men_men_n29_), .C(m), .Y(men_men_n630_));
  NAi32      u0602(.An(n), .Bn(f), .C(m), .Y(men_men_n631_));
  NOi32      u0603(.An(e), .Bn(a), .C(d), .Y(men_men_n632_));
  AOI210     u0604(.A0(men_men_n29_), .A1(d), .B0(men_men_n632_), .Y(men_men_n633_));
  AOI210     u0605(.A0(men_men_n633_), .A1(men_men_n224_), .B0(men_men_n575_), .Y(men_men_n634_));
  AOI210     u0606(.A0(men_men_n634_), .A1(men_men_n1620_), .B0(men_men_n626_), .Y(men_men_n635_));
  OAI210     u0607(.A0(men_men_n262_), .A1(men_men_n89_), .B0(men_men_n635_), .Y(men_men_n636_));
  AOI210     u0608(.A0(men_men_n621_), .A1(men_men_n610_), .B0(men_men_n636_), .Y(men_men_n637_));
  NO3        u0609(.A(men_men_n332_), .B(men_men_n61_), .C(n), .Y(men_men_n638_));
  NA3        u0610(.A(men_men_n534_), .B(men_men_n180_), .C(men_men_n179_), .Y(men_men_n639_));
  NA2        u0611(.A(men_men_n482_), .B(men_men_n242_), .Y(men_men_n640_));
  OR2        u0612(.A(men_men_n640_), .B(men_men_n639_), .Y(men_men_n641_));
  NA2        u0613(.A(men_men_n76_), .B(men_men_n117_), .Y(men_men_n642_));
  NO2        u0614(.A(men_men_n642_), .B(men_men_n45_), .Y(men_men_n643_));
  AOI220     u0615(.A0(men_men_n643_), .A1(men_men_n562_), .B0(men_men_n641_), .B1(men_men_n638_), .Y(men_men_n644_));
  NO2        u0616(.A(men_men_n644_), .B(men_men_n89_), .Y(men_men_n645_));
  NA3        u0617(.A(men_men_n577_), .B(men_men_n358_), .C(men_men_n46_), .Y(men_men_n646_));
  NOi32      u0618(.An(e), .Bn(c), .C(f), .Y(men_men_n647_));
  NOi21      u0619(.An(f), .B(u), .Y(men_men_n648_));
  NO2        u0620(.A(men_men_n648_), .B(men_men_n222_), .Y(men_men_n649_));
  AOI220     u0621(.A0(men_men_n649_), .A1(men_men_n413_), .B0(men_men_n647_), .B1(men_men_n184_), .Y(men_men_n650_));
  NA3        u0622(.A(men_men_n650_), .B(men_men_n646_), .C(men_men_n187_), .Y(men_men_n651_));
  AOI210     u0623(.A0(men_men_n561_), .A1(men_men_n417_), .B0(men_men_n313_), .Y(men_men_n652_));
  NA2        u0624(.A(men_men_n652_), .B(men_men_n279_), .Y(men_men_n653_));
  NOi21      u0625(.An(j), .B(l), .Y(men_men_n654_));
  NAi21      u0626(.An(k), .B(h), .Y(men_men_n655_));
  NO2        u0627(.A(men_men_n655_), .B(men_men_n277_), .Y(men_men_n656_));
  NA2        u0628(.A(men_men_n656_), .B(men_men_n654_), .Y(men_men_n657_));
  OR2        u0629(.A(men_men_n657_), .B(men_men_n615_), .Y(men_men_n658_));
  NOi31      u0630(.An(m), .B(n), .C(k), .Y(men_men_n659_));
  NA2        u0631(.A(men_men_n654_), .B(men_men_n659_), .Y(men_men_n660_));
  AOI210     u0632(.A0(men_men_n417_), .A1(men_men_n391_), .B0(men_men_n313_), .Y(men_men_n661_));
  NAi21      u0633(.An(men_men_n660_), .B(men_men_n661_), .Y(men_men_n662_));
  NO2        u0634(.A(men_men_n293_), .B(men_men_n49_), .Y(men_men_n663_));
  NO2        u0635(.A(men_men_n325_), .B(men_men_n622_), .Y(men_men_n664_));
  NO2        u0636(.A(men_men_n557_), .B(men_men_n49_), .Y(men_men_n665_));
  AOI220     u0637(.A0(men_men_n665_), .A1(men_men_n664_), .B0(men_men_n663_), .B1(men_men_n596_), .Y(men_men_n666_));
  NA4        u0638(.A(men_men_n666_), .B(men_men_n662_), .C(men_men_n658_), .D(men_men_n653_), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n112_), .B(men_men_n36_), .Y(men_men_n668_));
  NO2        u0640(.A(k), .B(men_men_n225_), .Y(men_men_n669_));
  NO2        u0641(.A(men_men_n553_), .B(men_men_n380_), .Y(men_men_n670_));
  NO2        u0642(.A(men_men_n670_), .B(n), .Y(men_men_n671_));
  NAi31      u0643(.An(men_men_n668_), .B(men_men_n671_), .C(men_men_n669_), .Y(men_men_n672_));
  NO2        u0644(.A(men_men_n555_), .B(men_men_n185_), .Y(men_men_n673_));
  NA3        u0645(.A(men_men_n578_), .B(men_men_n286_), .C(men_men_n150_), .Y(men_men_n674_));
  NA2        u0646(.A(men_men_n530_), .B(men_men_n166_), .Y(men_men_n675_));
  NO3        u0647(.A(men_men_n414_), .B(men_men_n675_), .C(men_men_n89_), .Y(men_men_n676_));
  AOI210     u0648(.A0(men_men_n674_), .A1(men_men_n673_), .B0(men_men_n676_), .Y(men_men_n677_));
  AN3        u0649(.A(f), .B(d), .C(b), .Y(men_men_n678_));
  OAI210     u0650(.A0(men_men_n678_), .A1(men_men_n135_), .B0(n), .Y(men_men_n679_));
  NA3        u0651(.A(men_men_n530_), .B(men_men_n166_), .C(men_men_n225_), .Y(men_men_n680_));
  AOI210     u0652(.A0(men_men_n679_), .A1(men_men_n244_), .B0(men_men_n680_), .Y(men_men_n681_));
  NAi31      u0653(.An(m), .B(n), .C(k), .Y(men_men_n682_));
  OR2        u0654(.A(men_men_n139_), .B(men_men_n61_), .Y(men_men_n683_));
  OAI210     u0655(.A0(men_men_n683_), .A1(men_men_n682_), .B0(men_men_n264_), .Y(men_men_n684_));
  OAI210     u0656(.A0(men_men_n684_), .A1(men_men_n681_), .B0(j), .Y(men_men_n685_));
  NA3        u0657(.A(men_men_n685_), .B(men_men_n677_), .C(men_men_n672_), .Y(men_men_n686_));
  NO4        u0658(.A(men_men_n686_), .B(men_men_n667_), .C(men_men_n651_), .D(men_men_n645_), .Y(men_men_n687_));
  NA2        u0659(.A(men_men_n401_), .B(men_men_n169_), .Y(men_men_n688_));
  NAi31      u0660(.An(u), .B(h), .C(f), .Y(men_men_n689_));
  OR3        u0661(.A(men_men_n689_), .B(men_men_n293_), .C(n), .Y(men_men_n690_));
  OA210      u0662(.A0(men_men_n557_), .A1(n), .B0(men_men_n613_), .Y(men_men_n691_));
  NA3        u0663(.A(men_men_n437_), .B(men_men_n125_), .C(men_men_n86_), .Y(men_men_n692_));
  OAI210     u0664(.A0(men_men_n691_), .A1(men_men_n93_), .B0(men_men_n692_), .Y(men_men_n693_));
  NOi21      u0665(.An(men_men_n690_), .B(men_men_n693_), .Y(men_men_n694_));
  AOI210     u0666(.A0(men_men_n694_), .A1(men_men_n688_), .B0(men_men_n551_), .Y(men_men_n695_));
  NO3        u0667(.A(u), .B(men_men_n224_), .C(men_men_n56_), .Y(men_men_n696_));
  NAi21      u0668(.An(h), .B(j), .Y(men_men_n697_));
  OAI220     u0669(.A0(men_men_n697_), .A1(men_men_n106_), .B0(men_men_n538_), .B1(men_men_n89_), .Y(men_men_n698_));
  OAI210     u0670(.A0(men_men_n698_), .A1(men_men_n413_), .B0(men_men_n696_), .Y(men_men_n699_));
  OR2        u0671(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n700_));
  NA2        u0672(.A(men_men_n624_), .B(men_men_n360_), .Y(men_men_n701_));
  OA220      u0673(.A0(men_men_n660_), .A1(men_men_n701_), .B0(men_men_n657_), .B1(men_men_n700_), .Y(men_men_n702_));
  NA3        u0674(.A(men_men_n548_), .B(men_men_n102_), .C(men_men_n101_), .Y(men_men_n703_));
  AN2        u0675(.A(h), .B(f), .Y(men_men_n704_));
  NA2        u0676(.A(men_men_n704_), .B(men_men_n37_), .Y(men_men_n705_));
  NA2        u0677(.A(men_men_n102_), .B(men_men_n46_), .Y(men_men_n706_));
  OAI220     u0678(.A0(men_men_n706_), .A1(men_men_n349_), .B0(men_men_n705_), .B1(men_men_n487_), .Y(men_men_n707_));
  AOI210     u0679(.A0(men_men_n594_), .A1(men_men_n448_), .B0(men_men_n49_), .Y(men_men_n708_));
  OAI220     u0680(.A0(men_men_n616_), .A1(men_men_n609_), .B0(men_men_n342_), .B1(men_men_n549_), .Y(men_men_n709_));
  AOI210     u0681(.A0(men_men_n709_), .A1(men_men_n708_), .B0(men_men_n707_), .Y(men_men_n710_));
  NA4        u0682(.A(men_men_n710_), .B(men_men_n703_), .C(men_men_n702_), .D(men_men_n699_), .Y(men_men_n711_));
  NO2        u0683(.A(men_men_n266_), .B(f), .Y(men_men_n712_));
  NO2        u0684(.A(men_men_n648_), .B(men_men_n61_), .Y(men_men_n713_));
  NO3        u0685(.A(men_men_n713_), .B(men_men_n712_), .C(men_men_n34_), .Y(men_men_n714_));
  NA2        u0686(.A(men_men_n345_), .B(men_men_n145_), .Y(men_men_n715_));
  NA2        u0687(.A(men_men_n137_), .B(men_men_n49_), .Y(men_men_n716_));
  AOI220     u0688(.A0(men_men_n716_), .A1(men_men_n553_), .B0(men_men_n380_), .B1(men_men_n117_), .Y(men_men_n717_));
  OA220      u0689(.A0(men_men_n717_), .A1(men_men_n575_), .B0(men_men_n378_), .B1(men_men_n115_), .Y(men_men_n718_));
  OAI210     u0690(.A0(men_men_n715_), .A1(men_men_n714_), .B0(men_men_n718_), .Y(men_men_n719_));
  NO3        u0691(.A(men_men_n424_), .B(men_men_n202_), .C(men_men_n201_), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n720_), .B(men_men_n242_), .Y(men_men_n721_));
  NA3        u0693(.A(men_men_n721_), .B(men_men_n268_), .C(j), .Y(men_men_n722_));
  NA2        u0694(.A(men_men_n486_), .B(men_men_n86_), .Y(men_men_n723_));
  NO4        u0695(.A(men_men_n551_), .B(men_men_n723_), .C(men_men_n136_), .D(men_men_n224_), .Y(men_men_n724_));
  INV        u0696(.A(men_men_n724_), .Y(men_men_n725_));
  NA4        u0697(.A(men_men_n725_), .B(men_men_n722_), .C(men_men_n537_), .D(men_men_n422_), .Y(men_men_n726_));
  NO4        u0698(.A(men_men_n726_), .B(men_men_n719_), .C(men_men_n711_), .D(men_men_n695_), .Y(men_men_n727_));
  NA4        u0699(.A(men_men_n727_), .B(men_men_n687_), .C(men_men_n637_), .D(men_men_n607_), .Y(men08));
  NO2        u0700(.A(k), .B(h), .Y(men_men_n729_));
  AO210      u0701(.A0(men_men_n266_), .A1(men_men_n470_), .B0(men_men_n729_), .Y(men_men_n730_));
  NO2        u0702(.A(men_men_n730_), .B(men_men_n311_), .Y(men_men_n731_));
  NA2        u0703(.A(men_men_n647_), .B(men_men_n86_), .Y(men_men_n732_));
  NA2        u0704(.A(men_men_n732_), .B(men_men_n482_), .Y(men_men_n733_));
  NA2        u0705(.A(men_men_n733_), .B(men_men_n731_), .Y(men_men_n734_));
  NA2        u0706(.A(men_men_n86_), .B(men_men_n114_), .Y(men_men_n735_));
  NO2        u0707(.A(men_men_n735_), .B(men_men_n57_), .Y(men_men_n736_));
  NO4        u0708(.A(men_men_n398_), .B(men_men_n116_), .C(j), .D(men_men_n225_), .Y(men_men_n737_));
  NA2        u0709(.A(men_men_n603_), .B(men_men_n244_), .Y(men_men_n738_));
  AOI220     u0710(.A0(men_men_n738_), .A1(men_men_n366_), .B0(men_men_n737_), .B1(men_men_n736_), .Y(men_men_n739_));
  AOI210     u0711(.A0(men_men_n603_), .A1(men_men_n162_), .B0(men_men_n86_), .Y(men_men_n740_));
  NA4        u0712(.A(men_men_n227_), .B(men_men_n145_), .C(men_men_n45_), .D(h), .Y(men_men_n741_));
  AN2        u0713(.A(l), .B(k), .Y(men_men_n742_));
  NA4        u0714(.A(men_men_n742_), .B(men_men_n112_), .C(men_men_n75_), .D(men_men_n225_), .Y(men_men_n743_));
  OAI210     u0715(.A0(men_men_n741_), .A1(u), .B0(men_men_n743_), .Y(men_men_n744_));
  NA2        u0716(.A(men_men_n744_), .B(men_men_n740_), .Y(men_men_n745_));
  NA4        u0717(.A(men_men_n745_), .B(men_men_n739_), .C(men_men_n734_), .D(men_men_n367_), .Y(men_men_n746_));
  AN2        u0718(.A(men_men_n558_), .B(men_men_n98_), .Y(men_men_n747_));
  NO4        u0719(.A(men_men_n182_), .B(men_men_n412_), .C(men_men_n116_), .D(u), .Y(men_men_n748_));
  AOI210     u0720(.A0(men_men_n748_), .A1(men_men_n738_), .B0(men_men_n543_), .Y(men_men_n749_));
  NO2        u0721(.A(men_men_n38_), .B(men_men_n224_), .Y(men_men_n750_));
  AOI220     u0722(.A0(men_men_n649_), .A1(men_men_n365_), .B0(men_men_n750_), .B1(men_men_n591_), .Y(men_men_n751_));
  NAi31      u0723(.An(men_men_n747_), .B(men_men_n751_), .C(men_men_n749_), .Y(men_men_n752_));
  NO2        u0724(.A(men_men_n561_), .B(men_men_n35_), .Y(men_men_n753_));
  OAI210     u0725(.A0(men_men_n578_), .A1(men_men_n47_), .B0(men_men_n683_), .Y(men_men_n754_));
  NO2        u0726(.A(men_men_n505_), .B(men_men_n137_), .Y(men_men_n755_));
  AOI210     u0727(.A0(men_men_n755_), .A1(men_men_n754_), .B0(men_men_n753_), .Y(men_men_n756_));
  NO3        u0728(.A(men_men_n332_), .B(men_men_n136_), .C(men_men_n41_), .Y(men_men_n757_));
  NAi21      u0729(.An(men_men_n757_), .B(men_men_n743_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n730_), .B(men_men_n140_), .Y(men_men_n759_));
  AOI220     u0731(.A0(men_men_n759_), .A1(men_men_n423_), .B0(men_men_n758_), .B1(men_men_n78_), .Y(men_men_n760_));
  OAI210     u0732(.A0(men_men_n756_), .A1(men_men_n89_), .B0(men_men_n760_), .Y(men_men_n761_));
  NA2        u0733(.A(men_men_n380_), .B(men_men_n43_), .Y(men_men_n762_));
  NA3        u0734(.A(men_men_n721_), .B(men_men_n351_), .C(men_men_n404_), .Y(men_men_n763_));
  NA2        u0735(.A(men_men_n742_), .B(men_men_n232_), .Y(men_men_n764_));
  NO2        u0736(.A(men_men_n764_), .B(men_men_n344_), .Y(men_men_n765_));
  AOI210     u0737(.A0(men_men_n765_), .A1(men_men_n712_), .B0(men_men_n512_), .Y(men_men_n766_));
  NA3        u0738(.A(m), .B(l), .C(k), .Y(men_men_n767_));
  AOI210     u0739(.A0(men_men_n692_), .A1(men_men_n690_), .B0(men_men_n767_), .Y(men_men_n768_));
  NO2        u0740(.A(men_men_n560_), .B(men_men_n287_), .Y(men_men_n769_));
  NOi21      u0741(.An(men_men_n769_), .B(men_men_n554_), .Y(men_men_n770_));
  NA4        u0742(.A(men_men_n117_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n771_));
  NA3        u0743(.A(men_men_n125_), .B(men_men_n432_), .C(i), .Y(men_men_n772_));
  NO2        u0744(.A(men_men_n772_), .B(men_men_n771_), .Y(men_men_n773_));
  NO3        u0745(.A(men_men_n773_), .B(men_men_n770_), .C(men_men_n768_), .Y(men_men_n774_));
  NA4        u0746(.A(men_men_n774_), .B(men_men_n766_), .C(men_men_n763_), .D(men_men_n762_), .Y(men_men_n775_));
  NO4        u0747(.A(men_men_n775_), .B(men_men_n761_), .C(men_men_n752_), .D(men_men_n746_), .Y(men_men_n776_));
  NA2        u0748(.A(men_men_n649_), .B(men_men_n413_), .Y(men_men_n777_));
  NOi31      u0749(.An(u), .B(h), .C(f), .Y(men_men_n778_));
  NA2        u0750(.A(men_men_n665_), .B(men_men_n778_), .Y(men_men_n779_));
  AO210      u0751(.A0(men_men_n779_), .A1(men_men_n617_), .B0(men_men_n563_), .Y(men_men_n780_));
  NO3        u0752(.A(men_men_n417_), .B(men_men_n549_), .C(h), .Y(men_men_n781_));
  AOI210     u0753(.A0(men_men_n781_), .A1(men_men_n117_), .B0(men_men_n523_), .Y(men_men_n782_));
  NA4        u0754(.A(men_men_n782_), .B(men_men_n780_), .C(men_men_n777_), .D(men_men_n265_), .Y(men_men_n783_));
  NA2        u0755(.A(men_men_n742_), .B(men_men_n75_), .Y(men_men_n784_));
  NO4        u0756(.A(men_men_n720_), .B(men_men_n182_), .C(n), .D(i), .Y(men_men_n785_));
  NOi21      u0757(.An(h), .B(j), .Y(men_men_n786_));
  NA2        u0758(.A(men_men_n786_), .B(f), .Y(men_men_n787_));
  NO2        u0759(.A(men_men_n787_), .B(men_men_n259_), .Y(men_men_n788_));
  NO2        u0760(.A(men_men_n788_), .B(men_men_n785_), .Y(men_men_n789_));
  OAI220     u0761(.A0(men_men_n789_), .A1(men_men_n784_), .B0(men_men_n619_), .B1(men_men_n62_), .Y(men_men_n790_));
  AOI210     u0762(.A0(men_men_n783_), .A1(l), .B0(men_men_n790_), .Y(men_men_n791_));
  NO2        u0763(.A(j), .B(i), .Y(men_men_n792_));
  NA3        u0764(.A(men_men_n792_), .B(men_men_n82_), .C(l), .Y(men_men_n793_));
  NA2        u0765(.A(men_men_n792_), .B(men_men_n33_), .Y(men_men_n794_));
  NA2        u0766(.A(men_men_n442_), .B(men_men_n125_), .Y(men_men_n795_));
  OA220      u0767(.A0(men_men_n795_), .A1(men_men_n794_), .B0(men_men_n793_), .B1(men_men_n615_), .Y(men_men_n796_));
  NO3        u0768(.A(men_men_n157_), .B(men_men_n49_), .C(men_men_n114_), .Y(men_men_n797_));
  NO3        u0769(.A(men_men_n567_), .B(men_men_n155_), .C(men_men_n75_), .Y(men_men_n798_));
  NO3        u0770(.A(men_men_n505_), .B(men_men_n460_), .C(j), .Y(men_men_n799_));
  OAI210     u0771(.A0(men_men_n798_), .A1(men_men_n797_), .B0(men_men_n799_), .Y(men_men_n800_));
  OAI210     u0772(.A0(men_men_n779_), .A1(men_men_n62_), .B0(men_men_n800_), .Y(men_men_n801_));
  NA2        u0773(.A(k), .B(j), .Y(men_men_n802_));
  NO3        u0774(.A(men_men_n311_), .B(men_men_n802_), .C(men_men_n40_), .Y(men_men_n803_));
  AOI210     u0775(.A0(men_men_n553_), .A1(n), .B0(men_men_n577_), .Y(men_men_n804_));
  NA2        u0776(.A(men_men_n804_), .B(men_men_n580_), .Y(men_men_n805_));
  AN3        u0777(.A(men_men_n805_), .B(men_men_n803_), .C(men_men_n101_), .Y(men_men_n806_));
  NO3        u0778(.A(men_men_n182_), .B(men_men_n412_), .C(men_men_n116_), .Y(men_men_n807_));
  AOI220     u0779(.A0(men_men_n807_), .A1(men_men_n260_), .B0(men_men_n640_), .B1(men_men_n322_), .Y(men_men_n808_));
  NAi31      u0780(.An(men_men_n633_), .B(men_men_n95_), .C(men_men_n86_), .Y(men_men_n809_));
  NA2        u0781(.A(men_men_n809_), .B(men_men_n808_), .Y(men_men_n810_));
  NO2        u0782(.A(men_men_n311_), .B(men_men_n140_), .Y(men_men_n811_));
  AOI220     u0783(.A0(men_men_n811_), .A1(men_men_n649_), .B0(men_men_n757_), .B1(men_men_n740_), .Y(men_men_n812_));
  NO2        u0784(.A(men_men_n616_), .B(men_men_n121_), .Y(men_men_n813_));
  OAI210     u0785(.A0(men_men_n813_), .A1(men_men_n799_), .B0(men_men_n708_), .Y(men_men_n814_));
  NA2        u0786(.A(men_men_n814_), .B(men_men_n812_), .Y(men_men_n815_));
  OR4        u0787(.A(men_men_n815_), .B(men_men_n810_), .C(men_men_n806_), .D(men_men_n801_), .Y(men_men_n816_));
  NA3        u0788(.A(men_men_n804_), .B(men_men_n580_), .C(men_men_n579_), .Y(men_men_n817_));
  NA4        u0789(.A(men_men_n817_), .B(men_men_n227_), .C(men_men_n470_), .D(men_men_n34_), .Y(men_men_n818_));
  NO4        u0790(.A(men_men_n505_), .B(men_men_n455_), .C(j), .D(f), .Y(men_men_n819_));
  OAI220     u0791(.A0(men_men_n741_), .A1(men_men_n732_), .B0(men_men_n349_), .B1(men_men_n38_), .Y(men_men_n820_));
  AOI210     u0792(.A0(men_men_n819_), .A1(men_men_n272_), .B0(men_men_n820_), .Y(men_men_n821_));
  NA3        u0793(.A(men_men_n570_), .B(men_men_n308_), .C(h), .Y(men_men_n822_));
  NO2        u0794(.A(men_men_n94_), .B(men_men_n47_), .Y(men_men_n823_));
  OAI220     u0795(.A0(men_men_n822_), .A1(men_men_n630_), .B0(men_men_n793_), .B1(men_men_n700_), .Y(men_men_n824_));
  AOI210     u0796(.A0(men_men_n823_), .A1(men_men_n671_), .B0(men_men_n824_), .Y(men_men_n825_));
  NA3        u0797(.A(men_men_n825_), .B(men_men_n821_), .C(men_men_n818_), .Y(men_men_n826_));
  BUFFER     u0798(.A(men_men_n98_), .Y(men_men_n827_));
  AOI220     u0799(.A0(men_men_n827_), .A1(men_men_n250_), .B0(men_men_n799_), .B1(men_men_n663_), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n691_), .B(men_men_n75_), .Y(men_men_n829_));
  AOI210     u0801(.A0(men_men_n819_), .A1(men_men_n829_), .B0(men_men_n353_), .Y(men_men_n830_));
  OAI210     u0802(.A0(men_men_n767_), .A1(men_men_n689_), .B0(men_men_n542_), .Y(men_men_n831_));
  NA3        u0803(.A(men_men_n263_), .B(men_men_n59_), .C(b), .Y(men_men_n832_));
  AOI220     u0804(.A0(men_men_n629_), .A1(men_men_n29_), .B0(men_men_n486_), .B1(men_men_n86_), .Y(men_men_n833_));
  NA2        u0805(.A(men_men_n833_), .B(men_men_n832_), .Y(men_men_n834_));
  NO2        u0806(.A(men_men_n822_), .B(men_men_n511_), .Y(men_men_n835_));
  AOI210     u0807(.A0(men_men_n834_), .A1(men_men_n831_), .B0(men_men_n835_), .Y(men_men_n836_));
  NA3        u0808(.A(men_men_n836_), .B(men_men_n830_), .C(men_men_n828_), .Y(men_men_n837_));
  NOi41      u0809(.An(men_men_n796_), .B(men_men_n837_), .C(men_men_n826_), .D(men_men_n816_), .Y(men_men_n838_));
  OR3        u0810(.A(men_men_n741_), .B(men_men_n244_), .C(u), .Y(men_men_n839_));
  NO3        u0811(.A(men_men_n359_), .B(men_men_n313_), .C(men_men_n116_), .Y(men_men_n840_));
  NA2        u0812(.A(men_men_n840_), .B(men_men_n805_), .Y(men_men_n841_));
  NA2        u0813(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n842_));
  NO3        u0814(.A(men_men_n842_), .B(men_men_n794_), .C(men_men_n293_), .Y(men_men_n843_));
  NO3        u0815(.A(men_men_n549_), .B(men_men_n96_), .C(h), .Y(men_men_n844_));
  AOI210     u0816(.A0(men_men_n844_), .A1(men_men_n736_), .B0(men_men_n843_), .Y(men_men_n845_));
  NA4        u0817(.A(men_men_n845_), .B(men_men_n841_), .C(men_men_n839_), .D(men_men_n425_), .Y(men_men_n846_));
  OR2        u0818(.A(men_men_n689_), .B(men_men_n94_), .Y(men_men_n847_));
  NOi31      u0819(.An(b), .B(d), .C(a), .Y(men_men_n848_));
  NO2        u0820(.A(men_men_n848_), .B(men_men_n627_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n849_), .B(n), .Y(men_men_n850_));
  NOi21      u0822(.An(men_men_n833_), .B(men_men_n850_), .Y(men_men_n851_));
  OAI220     u0823(.A0(men_men_n851_), .A1(men_men_n847_), .B0(men_men_n822_), .B1(men_men_n628_), .Y(men_men_n852_));
  NO2        u0824(.A(men_men_n578_), .B(men_men_n86_), .Y(men_men_n853_));
  NO3        u0825(.A(men_men_n648_), .B(men_men_n344_), .C(men_men_n121_), .Y(men_men_n854_));
  NOi21      u0826(.An(men_men_n854_), .B(men_men_n167_), .Y(men_men_n855_));
  AOI210     u0827(.A0(men_men_n840_), .A1(men_men_n853_), .B0(men_men_n855_), .Y(men_men_n856_));
  OAI210     u0828(.A0(men_men_n741_), .A1(men_men_n414_), .B0(men_men_n856_), .Y(men_men_n857_));
  NO2        u0829(.A(men_men_n720_), .B(n), .Y(men_men_n858_));
  AOI220     u0830(.A0(men_men_n811_), .A1(men_men_n696_), .B0(men_men_n858_), .B1(men_men_n731_), .Y(men_men_n859_));
  NO2        u0831(.A(men_men_n339_), .B(men_men_n249_), .Y(men_men_n860_));
  OAI210     u0832(.A0(men_men_n98_), .A1(men_men_n95_), .B0(men_men_n860_), .Y(men_men_n861_));
  NA2        u0833(.A(men_men_n125_), .B(men_men_n86_), .Y(men_men_n862_));
  AOI210     u0834(.A0(men_men_n446_), .A1(men_men_n438_), .B0(men_men_n862_), .Y(men_men_n863_));
  NAi21      u0835(.An(men_men_n863_), .B(men_men_n861_), .Y(men_men_n864_));
  NA2        u0836(.A(men_men_n765_), .B(men_men_n34_), .Y(men_men_n865_));
  NAi21      u0837(.An(men_men_n771_), .B(men_men_n456_), .Y(men_men_n866_));
  NO2        u0838(.A(men_men_n287_), .B(i), .Y(men_men_n867_));
  NAi41      u0839(.An(men_men_n864_), .B(men_men_n866_), .C(men_men_n865_), .D(men_men_n859_), .Y(men_men_n868_));
  NO4        u0840(.A(men_men_n868_), .B(men_men_n857_), .C(men_men_n852_), .D(men_men_n846_), .Y(men_men_n869_));
  NA4        u0841(.A(men_men_n869_), .B(men_men_n838_), .C(men_men_n791_), .D(men_men_n776_), .Y(men09));
  INV        u0842(.A(men_men_n126_), .Y(men_men_n871_));
  NA2        u0843(.A(f), .B(e), .Y(men_men_n872_));
  NO2        u0844(.A(men_men_n237_), .B(men_men_n116_), .Y(men_men_n873_));
  NA2        u0845(.A(men_men_n873_), .B(u), .Y(men_men_n874_));
  NA4        u0846(.A(men_men_n325_), .B(men_men_n172_), .C(men_men_n275_), .D(men_men_n123_), .Y(men_men_n875_));
  AOI210     u0847(.A0(men_men_n875_), .A1(u), .B0(men_men_n492_), .Y(men_men_n876_));
  AOI210     u0848(.A0(men_men_n876_), .A1(men_men_n874_), .B0(men_men_n872_), .Y(men_men_n877_));
  NA2        u0849(.A(men_men_n463_), .B(e), .Y(men_men_n878_));
  NO2        u0850(.A(men_men_n878_), .B(men_men_n534_), .Y(men_men_n879_));
  AOI210     u0851(.A0(men_men_n877_), .A1(men_men_n871_), .B0(men_men_n879_), .Y(men_men_n880_));
  NO2        u0852(.A(men_men_n214_), .B(men_men_n224_), .Y(men_men_n881_));
  NA3        u0853(.A(m), .B(l), .C(i), .Y(men_men_n882_));
  OAI220     u0854(.A0(men_men_n616_), .A1(men_men_n882_), .B0(men_men_n371_), .B1(men_men_n550_), .Y(men_men_n883_));
  NA4        u0855(.A(men_men_n90_), .B(men_men_n89_), .C(u), .D(f), .Y(men_men_n884_));
  OA210      u0856(.A0(men_men_n883_), .A1(men_men_n881_), .B0(men_men_n591_), .Y(men_men_n885_));
  NA3        u0857(.A(men_men_n847_), .B(men_men_n593_), .C(men_men_n542_), .Y(men_men_n886_));
  OA210      u0858(.A0(men_men_n886_), .A1(men_men_n885_), .B0(men_men_n850_), .Y(men_men_n887_));
  INV        u0859(.A(men_men_n356_), .Y(men_men_n888_));
  NO2        u0860(.A(men_men_n132_), .B(men_men_n130_), .Y(men_men_n889_));
  NOi31      u0861(.An(k), .B(m), .C(l), .Y(men_men_n890_));
  NO2        u0862(.A(men_men_n358_), .B(men_men_n890_), .Y(men_men_n891_));
  AOI210     u0863(.A0(men_men_n891_), .A1(men_men_n889_), .B0(men_men_n622_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n832_), .B(men_men_n349_), .Y(men_men_n893_));
  NA2        u0865(.A(men_men_n360_), .B(men_men_n362_), .Y(men_men_n894_));
  OAI210     u0866(.A0(men_men_n214_), .A1(men_men_n224_), .B0(men_men_n894_), .Y(men_men_n895_));
  AOI220     u0867(.A0(men_men_n895_), .A1(men_men_n893_), .B0(men_men_n892_), .B1(men_men_n888_), .Y(men_men_n896_));
  NA2        u0868(.A(men_men_n176_), .B(men_men_n118_), .Y(men_men_n897_));
  NA3        u0869(.A(men_men_n897_), .B(men_men_n730_), .C(men_men_n140_), .Y(men_men_n898_));
  NA3        u0870(.A(men_men_n898_), .B(men_men_n199_), .C(men_men_n31_), .Y(men_men_n899_));
  NA4        u0871(.A(men_men_n899_), .B(men_men_n896_), .C(men_men_n650_), .D(men_men_n84_), .Y(men_men_n900_));
  NO2        u0872(.A(men_men_n612_), .B(men_men_n519_), .Y(men_men_n901_));
  NOi21      u0873(.An(f), .B(d), .Y(men_men_n902_));
  NA2        u0874(.A(men_men_n902_), .B(m), .Y(men_men_n903_));
  NO2        u0875(.A(men_men_n903_), .B(men_men_n52_), .Y(men_men_n904_));
  NOi32      u0876(.An(u), .Bn(f), .C(d), .Y(men_men_n905_));
  NA4        u0877(.A(men_men_n905_), .B(men_men_n629_), .C(men_men_n29_), .D(m), .Y(men_men_n906_));
  NOi21      u0878(.An(men_men_n326_), .B(men_men_n906_), .Y(men_men_n907_));
  AOI210     u0879(.A0(men_men_n904_), .A1(men_men_n568_), .B0(men_men_n907_), .Y(men_men_n908_));
  NA3        u0880(.A(men_men_n325_), .B(men_men_n275_), .C(men_men_n123_), .Y(men_men_n909_));
  AN2        u0881(.A(f), .B(d), .Y(men_men_n910_));
  NA3        u0882(.A(men_men_n498_), .B(men_men_n910_), .C(men_men_n86_), .Y(men_men_n911_));
  NO3        u0883(.A(men_men_n911_), .B(men_men_n75_), .C(men_men_n225_), .Y(men_men_n912_));
  NO2        u0884(.A(men_men_n301_), .B(men_men_n56_), .Y(men_men_n913_));
  NA2        u0885(.A(men_men_n909_), .B(men_men_n912_), .Y(men_men_n914_));
  NAi31      u0886(.An(men_men_n510_), .B(men_men_n914_), .C(men_men_n908_), .Y(men_men_n915_));
  NO4        u0887(.A(men_men_n648_), .B(men_men_n137_), .C(men_men_n344_), .D(men_men_n158_), .Y(men_men_n916_));
  NO2        u0888(.A(men_men_n682_), .B(men_men_n344_), .Y(men_men_n917_));
  AN2        u0889(.A(men_men_n917_), .B(men_men_n712_), .Y(men_men_n918_));
  NO3        u0890(.A(men_men_n918_), .B(men_men_n916_), .C(men_men_n246_), .Y(men_men_n919_));
  NA2        u0891(.A(men_men_n627_), .B(men_men_n86_), .Y(men_men_n920_));
  NO2        u0892(.A(men_men_n894_), .B(men_men_n920_), .Y(men_men_n921_));
  NA3        u0893(.A(men_men_n166_), .B(men_men_n112_), .C(men_men_n111_), .Y(men_men_n922_));
  OAI220     u0894(.A0(men_men_n911_), .A1(men_men_n450_), .B0(men_men_n356_), .B1(men_men_n922_), .Y(men_men_n923_));
  NOi41      u0895(.An(men_men_n235_), .B(men_men_n923_), .C(men_men_n921_), .D(men_men_n320_), .Y(men_men_n924_));
  NA2        u0896(.A(c), .B(men_men_n120_), .Y(men_men_n925_));
  NO2        u0897(.A(men_men_n925_), .B(men_men_n429_), .Y(men_men_n926_));
  NA3        u0898(.A(men_men_n926_), .B(men_men_n532_), .C(f), .Y(men_men_n927_));
  OR2        u0899(.A(men_men_n689_), .B(men_men_n564_), .Y(men_men_n928_));
  OAI210     u0900(.A0(men_men_n595_), .A1(men_men_n642_), .B0(men_men_n928_), .Y(men_men_n929_));
  NA2        u0901(.A(men_men_n849_), .B(men_men_n115_), .Y(men_men_n930_));
  NA2        u0902(.A(men_men_n930_), .B(men_men_n929_), .Y(men_men_n931_));
  NA4        u0903(.A(men_men_n931_), .B(men_men_n927_), .C(men_men_n924_), .D(men_men_n919_), .Y(men_men_n932_));
  NO4        u0904(.A(men_men_n932_), .B(men_men_n915_), .C(men_men_n900_), .D(men_men_n887_), .Y(men_men_n933_));
  NA2        u0905(.A(men_men_n116_), .B(j), .Y(men_men_n934_));
  AOI210     u0906(.A0(men_men_n832_), .A1(men_men_n349_), .B0(men_men_n884_), .Y(men_men_n935_));
  NO2        u0907(.A(men_men_n242_), .B(men_men_n236_), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n936_), .B(men_men_n239_), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n450_), .B(men_men_n872_), .Y(men_men_n938_));
  NA2        u0910(.A(men_men_n938_), .B(men_men_n585_), .Y(men_men_n939_));
  NA2        u0911(.A(men_men_n939_), .B(men_men_n937_), .Y(men_men_n940_));
  NA2        u0912(.A(e), .B(d), .Y(men_men_n941_));
  OAI220     u0913(.A0(men_men_n941_), .A1(c), .B0(men_men_n339_), .B1(d), .Y(men_men_n942_));
  NA3        u0914(.A(men_men_n942_), .B(men_men_n475_), .C(men_men_n530_), .Y(men_men_n943_));
  AOI210     u0915(.A0(men_men_n538_), .A1(men_men_n189_), .B0(men_men_n242_), .Y(men_men_n944_));
  AOI210     u0916(.A0(men_men_n649_), .A1(men_men_n365_), .B0(men_men_n944_), .Y(men_men_n945_));
  NA2        u0917(.A(men_men_n301_), .B(men_men_n172_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n912_), .B(men_men_n946_), .Y(men_men_n947_));
  NA3        u0919(.A(men_men_n175_), .B(men_men_n87_), .C(men_men_n34_), .Y(men_men_n948_));
  NA4        u0920(.A(men_men_n948_), .B(men_men_n947_), .C(men_men_n945_), .D(men_men_n943_), .Y(men_men_n949_));
  NO3        u0921(.A(men_men_n949_), .B(men_men_n940_), .C(men_men_n935_), .Y(men_men_n950_));
  NA2        u0922(.A(men_men_n888_), .B(men_men_n31_), .Y(men_men_n951_));
  AO210      u0923(.A0(men_men_n951_), .A1(men_men_n732_), .B0(men_men_n228_), .Y(men_men_n952_));
  OAI220     u0924(.A0(men_men_n648_), .A1(men_men_n61_), .B0(men_men_n313_), .B1(j), .Y(men_men_n953_));
  AOI220     u0925(.A0(men_men_n953_), .A1(men_men_n917_), .B0(men_men_n638_), .B1(men_men_n647_), .Y(men_men_n954_));
  OAI210     u0926(.A0(men_men_n878_), .A1(men_men_n179_), .B0(men_men_n954_), .Y(men_men_n955_));
  OAI210     u0927(.A0(men_men_n873_), .A1(men_men_n946_), .B0(men_men_n905_), .Y(men_men_n956_));
  NO2        u0928(.A(men_men_n956_), .B(men_men_n630_), .Y(men_men_n957_));
  AOI210     u0929(.A0(men_men_n122_), .A1(men_men_n121_), .B0(men_men_n274_), .Y(men_men_n958_));
  NO2        u0930(.A(men_men_n958_), .B(men_men_n906_), .Y(men_men_n959_));
  AO210      u0931(.A0(men_men_n893_), .A1(men_men_n883_), .B0(men_men_n959_), .Y(men_men_n960_));
  NOi31      u0932(.An(men_men_n568_), .B(men_men_n903_), .C(men_men_n309_), .Y(men_men_n961_));
  NO4        u0933(.A(men_men_n961_), .B(men_men_n960_), .C(men_men_n957_), .D(men_men_n955_), .Y(men_men_n962_));
  AO220      u0934(.A0(men_men_n475_), .A1(men_men_n786_), .B0(men_men_n184_), .B1(f), .Y(men_men_n963_));
  OAI210     u0935(.A0(men_men_n963_), .A1(men_men_n478_), .B0(men_men_n942_), .Y(men_men_n964_));
  NO2        u0936(.A(men_men_n460_), .B(men_men_n71_), .Y(men_men_n965_));
  OAI210     u0937(.A0(men_men_n886_), .A1(men_men_n965_), .B0(men_men_n736_), .Y(men_men_n966_));
  AN4        u0938(.A(men_men_n966_), .B(men_men_n964_), .C(men_men_n962_), .D(men_men_n952_), .Y(men_men_n967_));
  NA4        u0939(.A(men_men_n967_), .B(men_men_n950_), .C(men_men_n933_), .D(men_men_n880_), .Y(men12));
  NO2        u0940(.A(men_men_n473_), .B(c), .Y(men_men_n969_));
  NO4        u0941(.A(men_men_n462_), .B(men_men_n266_), .C(men_men_n608_), .D(men_men_n225_), .Y(men_men_n970_));
  NA2        u0942(.A(men_men_n970_), .B(men_men_n969_), .Y(men_men_n971_));
  NA2        u0943(.A(men_men_n568_), .B(men_men_n965_), .Y(men_men_n972_));
  NO2        u0944(.A(men_men_n473_), .B(men_men_n120_), .Y(men_men_n973_));
  NO2        u0945(.A(men_men_n889_), .B(men_men_n371_), .Y(men_men_n974_));
  NO2        u0946(.A(men_men_n689_), .B(men_men_n398_), .Y(men_men_n975_));
  AOI220     u0947(.A0(men_men_n975_), .A1(men_men_n566_), .B0(men_men_n974_), .B1(men_men_n973_), .Y(men_men_n976_));
  NA4        u0948(.A(men_men_n976_), .B(men_men_n972_), .C(men_men_n971_), .D(men_men_n461_), .Y(men_men_n977_));
  AOI210     u0949(.A0(men_men_n245_), .A1(men_men_n355_), .B0(men_men_n211_), .Y(men_men_n978_));
  OR2        u0950(.A(men_men_n978_), .B(men_men_n970_), .Y(men_men_n979_));
  AOI210     u0951(.A0(men_men_n352_), .A1(men_men_n410_), .B0(men_men_n225_), .Y(men_men_n980_));
  OAI210     u0952(.A0(men_men_n980_), .A1(men_men_n979_), .B0(men_men_n424_), .Y(men_men_n981_));
  NO2        u0953(.A(men_men_n668_), .B(men_men_n277_), .Y(men_men_n982_));
  NO2        u0954(.A(men_men_n616_), .B(men_men_n882_), .Y(men_men_n983_));
  AOI220     u0955(.A0(men_men_n983_), .A1(men_men_n591_), .B0(men_men_n860_), .B1(men_men_n982_), .Y(men_men_n984_));
  NO2        u0956(.A(men_men_n157_), .B(men_men_n249_), .Y(men_men_n985_));
  NA3        u0957(.A(men_men_n985_), .B(men_men_n252_), .C(i), .Y(men_men_n986_));
  NA3        u0958(.A(men_men_n986_), .B(men_men_n984_), .C(men_men_n981_), .Y(men_men_n987_));
  OR2        u0959(.A(men_men_n340_), .B(men_men_n973_), .Y(men_men_n988_));
  NA2        u0960(.A(men_men_n988_), .B(men_men_n372_), .Y(men_men_n989_));
  NA4        u0961(.A(men_men_n463_), .B(men_men_n458_), .C(men_men_n190_), .D(u), .Y(men_men_n990_));
  NA2        u0962(.A(men_men_n990_), .B(men_men_n989_), .Y(men_men_n991_));
  NO3        u0963(.A(men_men_n694_), .B(men_men_n94_), .C(men_men_n45_), .Y(men_men_n992_));
  NO4        u0964(.A(men_men_n992_), .B(men_men_n991_), .C(men_men_n987_), .D(men_men_n977_), .Y(men_men_n993_));
  NO2        u0965(.A(men_men_n388_), .B(men_men_n387_), .Y(men_men_n994_));
  INV        u0966(.A(men_men_n613_), .Y(men_men_n995_));
  NA2        u0967(.A(men_men_n578_), .B(men_men_n150_), .Y(men_men_n996_));
  NOi21      u0968(.An(men_men_n34_), .B(men_men_n682_), .Y(men_men_n997_));
  AOI220     u0969(.A0(men_men_n997_), .A1(men_men_n996_), .B0(men_men_n995_), .B1(men_men_n994_), .Y(men_men_n998_));
  OAI210     u0970(.A0(men_men_n264_), .A1(men_men_n45_), .B0(men_men_n998_), .Y(men_men_n999_));
  NA2        u0971(.A(men_men_n456_), .B(men_men_n279_), .Y(men_men_n1000_));
  NO3        u0972(.A(men_men_n862_), .B(men_men_n91_), .C(men_men_n429_), .Y(men_men_n1001_));
  NAi31      u0973(.An(men_men_n1001_), .B(men_men_n1000_), .C(men_men_n336_), .Y(men_men_n1002_));
  NO2        u0974(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n1003_));
  NO2        u0975(.A(men_men_n526_), .B(men_men_n313_), .Y(men_men_n1004_));
  NO2        u0976(.A(men_men_n1004_), .B(men_men_n384_), .Y(men_men_n1005_));
  NO2        u0977(.A(men_men_n1005_), .B(men_men_n150_), .Y(men_men_n1006_));
  NA2        u0978(.A(men_men_n659_), .B(men_men_n381_), .Y(men_men_n1007_));
  OAI210     u0979(.A0(men_men_n772_), .A1(men_men_n1007_), .B0(men_men_n385_), .Y(men_men_n1008_));
  NO4        u0980(.A(men_men_n1008_), .B(men_men_n1006_), .C(men_men_n1002_), .D(men_men_n999_), .Y(men_men_n1009_));
  NA2        u0981(.A(men_men_n365_), .B(u), .Y(men_men_n1010_));
  NA2        u0982(.A(men_men_n169_), .B(i), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n46_), .B(i), .Y(men_men_n1012_));
  OAI220     u0984(.A0(men_men_n1012_), .A1(men_men_n210_), .B0(men_men_n1011_), .B1(men_men_n94_), .Y(men_men_n1013_));
  AOI210     u0985(.A0(men_men_n440_), .A1(men_men_n37_), .B0(men_men_n1013_), .Y(men_men_n1014_));
  NA2        u0986(.A(men_men_n578_), .B(men_men_n402_), .Y(men_men_n1015_));
  AOI210     u0987(.A0(men_men_n1015_), .A1(n), .B0(men_men_n577_), .Y(men_men_n1016_));
  OAI220     u0988(.A0(men_men_n1016_), .A1(men_men_n1010_), .B0(men_men_n1014_), .B1(men_men_n349_), .Y(men_men_n1017_));
  NO2        u0989(.A(men_men_n689_), .B(men_men_n519_), .Y(men_men_n1018_));
  NA3        u0990(.A(men_men_n360_), .B(men_men_n654_), .C(i), .Y(men_men_n1019_));
  OAI210     u0991(.A0(men_men_n460_), .A1(men_men_n325_), .B0(men_men_n1019_), .Y(men_men_n1020_));
  OAI220     u0992(.A0(men_men_n1020_), .A1(men_men_n1018_), .B0(men_men_n708_), .B1(men_men_n798_), .Y(men_men_n1021_));
  NA2        u0993(.A(men_men_n632_), .B(men_men_n117_), .Y(men_men_n1022_));
  OR3        u0994(.A(men_men_n325_), .B(men_men_n455_), .C(f), .Y(men_men_n1023_));
  NA3        u0995(.A(men_men_n654_), .B(men_men_n82_), .C(i), .Y(men_men_n1024_));
  OA220      u0996(.A0(men_men_n1024_), .A1(men_men_n1022_), .B0(men_men_n1023_), .B1(men_men_n615_), .Y(men_men_n1025_));
  NA3        u0997(.A(men_men_n341_), .B(men_men_n122_), .C(u), .Y(men_men_n1026_));
  AOI210     u0998(.A0(men_men_n705_), .A1(men_men_n1026_), .B0(m), .Y(men_men_n1027_));
  OAI210     u0999(.A0(men_men_n1027_), .A1(men_men_n974_), .B0(men_men_n340_), .Y(men_men_n1028_));
  NA2        u1000(.A(men_men_n723_), .B(men_men_n920_), .Y(men_men_n1029_));
  INV        u1001(.A(men_men_n884_), .Y(men_men_n1030_));
  NA2        u1002(.A(men_men_n233_), .B(men_men_n79_), .Y(men_men_n1031_));
  NA3        u1003(.A(men_men_n1031_), .B(men_men_n1024_), .C(men_men_n1023_), .Y(men_men_n1032_));
  AOI220     u1004(.A0(men_men_n1032_), .A1(men_men_n272_), .B0(men_men_n1030_), .B1(men_men_n1029_), .Y(men_men_n1033_));
  NA4        u1005(.A(men_men_n1033_), .B(men_men_n1028_), .C(men_men_n1025_), .D(men_men_n1021_), .Y(men_men_n1034_));
  NA2        u1006(.A(men_men_n693_), .B(men_men_n90_), .Y(men_men_n1035_));
  NO2        u1007(.A(men_men_n481_), .B(men_men_n225_), .Y(men_men_n1036_));
  AOI220     u1008(.A0(men_men_n1036_), .A1(men_men_n403_), .B0(men_men_n988_), .B1(men_men_n229_), .Y(men_men_n1037_));
  AOI220     u1009(.A0(men_men_n975_), .A1(men_men_n985_), .B0(men_men_n614_), .B1(men_men_n92_), .Y(men_men_n1038_));
  NA3        u1010(.A(men_men_n1038_), .B(men_men_n1037_), .C(men_men_n1035_), .Y(men_men_n1039_));
  OAI210     u1011(.A0(men_men_n1030_), .A1(men_men_n983_), .B0(men_men_n566_), .Y(men_men_n1040_));
  AOI210     u1012(.A0(men_men_n441_), .A1(men_men_n433_), .B0(men_men_n862_), .Y(men_men_n1041_));
  OAI210     u1013(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n113_), .Y(men_men_n1042_));
  AOI210     u1014(.A0(men_men_n1042_), .A1(men_men_n558_), .B0(men_men_n1041_), .Y(men_men_n1043_));
  NA2        u1015(.A(men_men_n1027_), .B(men_men_n973_), .Y(men_men_n1044_));
  NO3        u1016(.A(men_men_n934_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1045_));
  AOI220     u1017(.A0(men_men_n1045_), .A1(men_men_n652_), .B0(men_men_n673_), .B1(men_men_n553_), .Y(men_men_n1046_));
  NA4        u1018(.A(men_men_n1046_), .B(men_men_n1044_), .C(men_men_n1043_), .D(men_men_n1040_), .Y(men_men_n1047_));
  NO4        u1019(.A(men_men_n1047_), .B(men_men_n1039_), .C(men_men_n1034_), .D(men_men_n1017_), .Y(men_men_n1048_));
  NAi31      u1020(.An(men_men_n146_), .B(men_men_n442_), .C(n), .Y(men_men_n1049_));
  NO3        u1021(.A(men_men_n130_), .B(men_men_n358_), .C(men_men_n890_), .Y(men_men_n1050_));
  NO2        u1022(.A(men_men_n1050_), .B(men_men_n1049_), .Y(men_men_n1051_));
  NO3        u1023(.A(men_men_n287_), .B(men_men_n146_), .C(men_men_n429_), .Y(men_men_n1052_));
  AOI210     u1024(.A0(men_men_n1052_), .A1(men_men_n520_), .B0(men_men_n1051_), .Y(men_men_n1053_));
  INV        u1025(.A(men_men_n1053_), .Y(men_men_n1054_));
  NA2        u1026(.A(men_men_n242_), .B(men_men_n180_), .Y(men_men_n1055_));
  NO3        u1027(.A(men_men_n322_), .B(men_men_n463_), .C(men_men_n184_), .Y(men_men_n1056_));
  NOi31      u1028(.An(men_men_n1055_), .B(men_men_n1056_), .C(men_men_n225_), .Y(men_men_n1057_));
  NAi21      u1029(.An(men_men_n578_), .B(men_men_n1036_), .Y(men_men_n1058_));
  NA2        u1030(.A(men_men_n459_), .B(men_men_n920_), .Y(men_men_n1059_));
  NO3        u1031(.A(men_men_n460_), .B(men_men_n325_), .C(men_men_n75_), .Y(men_men_n1060_));
  AOI220     u1032(.A0(men_men_n1060_), .A1(men_men_n1059_), .B0(men_men_n502_), .B1(u), .Y(men_men_n1061_));
  NA2        u1033(.A(men_men_n1061_), .B(men_men_n1058_), .Y(men_men_n1062_));
  OAI220     u1034(.A0(men_men_n1049_), .A1(men_men_n245_), .B0(men_men_n1019_), .B1(men_men_n628_), .Y(men_men_n1063_));
  NO2        u1035(.A(men_men_n690_), .B(men_men_n398_), .Y(men_men_n1064_));
  NA2        u1036(.A(men_men_n978_), .B(men_men_n969_), .Y(men_men_n1065_));
  NO3        u1037(.A(men_men_n567_), .B(men_men_n155_), .C(men_men_n224_), .Y(men_men_n1066_));
  OAI210     u1038(.A0(men_men_n1066_), .A1(men_men_n548_), .B0(men_men_n399_), .Y(men_men_n1067_));
  OAI220     u1039(.A0(men_men_n975_), .A1(men_men_n983_), .B0(men_men_n568_), .B1(men_men_n449_), .Y(men_men_n1068_));
  NA4        u1040(.A(men_men_n1068_), .B(men_men_n1067_), .C(men_men_n1065_), .D(men_men_n646_), .Y(men_men_n1069_));
  OAI210     u1041(.A0(men_men_n978_), .A1(men_men_n970_), .B0(men_men_n1055_), .Y(men_men_n1070_));
  NA3        u1042(.A(men_men_n1015_), .B(men_men_n507_), .C(men_men_n46_), .Y(men_men_n1071_));
  AOI210     u1043(.A0(men_men_n401_), .A1(men_men_n399_), .B0(men_men_n348_), .Y(men_men_n1072_));
  NA4        u1044(.A(men_men_n1072_), .B(men_men_n1071_), .C(men_men_n1070_), .D(men_men_n288_), .Y(men_men_n1073_));
  OR4        u1045(.A(men_men_n1073_), .B(men_men_n1069_), .C(men_men_n1064_), .D(men_men_n1063_), .Y(men_men_n1074_));
  NO4        u1046(.A(men_men_n1074_), .B(men_men_n1062_), .C(men_men_n1057_), .D(men_men_n1054_), .Y(men_men_n1075_));
  NA4        u1047(.A(men_men_n1075_), .B(men_men_n1048_), .C(men_men_n1009_), .D(men_men_n993_), .Y(men13));
  NA2        u1048(.A(men_men_n46_), .B(men_men_n89_), .Y(men_men_n1077_));
  AN2        u1049(.A(c), .B(b), .Y(men_men_n1078_));
  NA3        u1050(.A(men_men_n263_), .B(men_men_n1078_), .C(m), .Y(men_men_n1079_));
  NA2        u1051(.A(men_men_n517_), .B(f), .Y(men_men_n1080_));
  NO4        u1052(.A(men_men_n1080_), .B(men_men_n1079_), .C(men_men_n1077_), .D(men_men_n609_), .Y(men_men_n1081_));
  NA2        u1053(.A(men_men_n279_), .B(men_men_n1078_), .Y(men_men_n1082_));
  NO4        u1054(.A(men_men_n1082_), .B(men_men_n1080_), .C(men_men_n1011_), .D(a), .Y(men_men_n1083_));
  NAi32      u1055(.An(d), .Bn(c), .C(e), .Y(men_men_n1084_));
  NA2        u1056(.A(men_men_n145_), .B(men_men_n45_), .Y(men_men_n1085_));
  NO4        u1057(.A(men_men_n1085_), .B(men_men_n1084_), .C(men_men_n616_), .D(men_men_n321_), .Y(men_men_n1086_));
  NA2        u1058(.A(men_men_n697_), .B(men_men_n236_), .Y(men_men_n1087_));
  NA2        u1059(.A(men_men_n432_), .B(men_men_n224_), .Y(men_men_n1088_));
  AN2        u1060(.A(d), .B(c), .Y(men_men_n1089_));
  NA2        u1061(.A(men_men_n1089_), .B(men_men_n120_), .Y(men_men_n1090_));
  NO4        u1062(.A(men_men_n1090_), .B(men_men_n1088_), .C(men_men_n185_), .D(men_men_n176_), .Y(men_men_n1091_));
  NA2        u1063(.A(men_men_n517_), .B(c), .Y(men_men_n1092_));
  NO4        u1064(.A(men_men_n1085_), .B(men_men_n612_), .C(men_men_n1092_), .D(men_men_n321_), .Y(men_men_n1093_));
  AO210      u1065(.A0(men_men_n1091_), .A1(men_men_n1087_), .B0(men_men_n1093_), .Y(men_men_n1094_));
  OR4        u1066(.A(men_men_n1094_), .B(men_men_n1086_), .C(men_men_n1083_), .D(men_men_n1081_), .Y(men_men_n1095_));
  NAi32      u1067(.An(f), .Bn(e), .C(c), .Y(men_men_n1096_));
  NO2        u1068(.A(men_men_n1096_), .B(men_men_n152_), .Y(men_men_n1097_));
  NA2        u1069(.A(men_men_n1097_), .B(u), .Y(men_men_n1098_));
  OR3        u1070(.A(men_men_n236_), .B(men_men_n185_), .C(men_men_n176_), .Y(men_men_n1099_));
  NO2        u1071(.A(men_men_n1099_), .B(men_men_n1098_), .Y(men_men_n1100_));
  NO2        u1072(.A(men_men_n1092_), .B(men_men_n321_), .Y(men_men_n1101_));
  NO2        u1073(.A(j), .B(men_men_n45_), .Y(men_men_n1102_));
  NA2        u1074(.A(men_men_n656_), .B(men_men_n1102_), .Y(men_men_n1103_));
  NOi21      u1075(.An(men_men_n1101_), .B(men_men_n1103_), .Y(men_men_n1104_));
  NO2        u1076(.A(men_men_n802_), .B(men_men_n116_), .Y(men_men_n1105_));
  NOi41      u1077(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1106_));
  NA2        u1078(.A(men_men_n1106_), .B(men_men_n1105_), .Y(men_men_n1107_));
  NO2        u1079(.A(men_men_n1107_), .B(men_men_n1098_), .Y(men_men_n1108_));
  OR3        u1080(.A(e), .B(d), .C(c), .Y(men_men_n1109_));
  NA3        u1081(.A(k), .B(j), .C(i), .Y(men_men_n1110_));
  NO3        u1082(.A(men_men_n1110_), .B(men_men_n321_), .C(men_men_n93_), .Y(men_men_n1111_));
  NOi21      u1083(.An(men_men_n1111_), .B(men_men_n1109_), .Y(men_men_n1112_));
  OR4        u1084(.A(men_men_n1112_), .B(men_men_n1108_), .C(men_men_n1104_), .D(men_men_n1100_), .Y(men_men_n1113_));
  NA3        u1085(.A(men_men_n489_), .B(men_men_n351_), .C(men_men_n56_), .Y(men_men_n1114_));
  NO2        u1086(.A(men_men_n1114_), .B(men_men_n1103_), .Y(men_men_n1115_));
  NO4        u1087(.A(men_men_n1114_), .B(men_men_n612_), .C(men_men_n470_), .D(men_men_n45_), .Y(men_men_n1116_));
  NO2        u1088(.A(f), .B(c), .Y(men_men_n1117_));
  NOi21      u1089(.An(men_men_n1117_), .B(men_men_n462_), .Y(men_men_n1118_));
  NA2        u1090(.A(men_men_n1118_), .B(men_men_n59_), .Y(men_men_n1119_));
  OR2        u1091(.A(k), .B(i), .Y(men_men_n1120_));
  NO3        u1092(.A(men_men_n1120_), .B(men_men_n256_), .C(l), .Y(men_men_n1121_));
  NOi31      u1093(.An(men_men_n1121_), .B(men_men_n1119_), .C(j), .Y(men_men_n1122_));
  OR3        u1094(.A(men_men_n1122_), .B(men_men_n1116_), .C(men_men_n1115_), .Y(men_men_n1123_));
  OR3        u1095(.A(men_men_n1123_), .B(men_men_n1113_), .C(men_men_n1095_), .Y(men02));
  OR2        u1096(.A(l), .B(k), .Y(men_men_n1125_));
  OR3        u1097(.A(h), .B(u), .C(f), .Y(men_men_n1126_));
  OR3        u1098(.A(n), .B(m), .C(i), .Y(men_men_n1127_));
  NO4        u1099(.A(men_men_n1127_), .B(men_men_n1126_), .C(men_men_n1125_), .D(men_men_n1109_), .Y(men_men_n1128_));
  NOi31      u1100(.An(e), .B(d), .C(c), .Y(men_men_n1129_));
  AOI210     u1101(.A0(men_men_n1111_), .A1(men_men_n1129_), .B0(men_men_n1086_), .Y(men_men_n1130_));
  AN3        u1102(.A(u), .B(f), .C(c), .Y(men_men_n1131_));
  NA3        u1103(.A(men_men_n1131_), .B(men_men_n489_), .C(h), .Y(men_men_n1132_));
  OR2        u1104(.A(men_men_n1110_), .B(men_men_n321_), .Y(men_men_n1133_));
  OR2        u1105(.A(men_men_n1133_), .B(men_men_n1132_), .Y(men_men_n1134_));
  NO3        u1106(.A(men_men_n1114_), .B(men_men_n1085_), .C(men_men_n612_), .Y(men_men_n1135_));
  NO2        u1107(.A(men_men_n1135_), .B(men_men_n1100_), .Y(men_men_n1136_));
  NA3        u1108(.A(l), .B(k), .C(j), .Y(men_men_n1137_));
  NA2        u1109(.A(i), .B(h), .Y(men_men_n1138_));
  NO3        u1110(.A(men_men_n1138_), .B(men_men_n1137_), .C(men_men_n137_), .Y(men_men_n1139_));
  NO3        u1111(.A(men_men_n147_), .B(men_men_n299_), .C(men_men_n225_), .Y(men_men_n1140_));
  AOI210     u1112(.A0(men_men_n1140_), .A1(men_men_n1139_), .B0(men_men_n1104_), .Y(men_men_n1141_));
  NA3        u1113(.A(c), .B(b), .C(a), .Y(men_men_n1142_));
  NO3        u1114(.A(men_men_n1142_), .B(men_men_n941_), .C(men_men_n224_), .Y(men_men_n1143_));
  NO4        u1115(.A(men_men_n1110_), .B(men_men_n313_), .C(men_men_n49_), .D(men_men_n116_), .Y(men_men_n1144_));
  AOI210     u1116(.A0(men_men_n1144_), .A1(men_men_n1143_), .B0(men_men_n1115_), .Y(men_men_n1145_));
  AN4        u1117(.A(men_men_n1145_), .B(men_men_n1141_), .C(men_men_n1136_), .D(men_men_n1134_), .Y(men_men_n1146_));
  NO2        u1118(.A(men_men_n1090_), .B(men_men_n1088_), .Y(men_men_n1147_));
  NA2        u1119(.A(men_men_n1107_), .B(men_men_n1099_), .Y(men_men_n1148_));
  AOI210     u1120(.A0(men_men_n1148_), .A1(men_men_n1147_), .B0(men_men_n1081_), .Y(men_men_n1149_));
  NAi41      u1121(.An(men_men_n1128_), .B(men_men_n1149_), .C(men_men_n1146_), .D(men_men_n1130_), .Y(men03));
  NO2        u1122(.A(men_men_n550_), .B(men_men_n622_), .Y(men_men_n1151_));
  NA4        u1123(.A(men_men_n90_), .B(men_men_n89_), .C(u), .D(men_men_n224_), .Y(men_men_n1152_));
  NA4        u1124(.A(men_men_n600_), .B(m), .C(men_men_n116_), .D(men_men_n224_), .Y(men_men_n1153_));
  NA3        u1125(.A(men_men_n1153_), .B(men_men_n389_), .C(men_men_n1152_), .Y(men_men_n1154_));
  NO3        u1126(.A(men_men_n1154_), .B(men_men_n1151_), .C(men_men_n1042_), .Y(men_men_n1155_));
  NO3        u1127(.A(men_men_n895_), .B(men_men_n883_), .C(men_men_n750_), .Y(men_men_n1156_));
  OAI220     u1128(.A0(men_men_n1156_), .A1(men_men_n723_), .B0(men_men_n1155_), .B1(men_men_n613_), .Y(men_men_n1157_));
  NOi31      u1129(.An(i), .B(k), .C(j), .Y(men_men_n1158_));
  NA4        u1130(.A(men_men_n1158_), .B(men_men_n1129_), .C(men_men_n360_), .D(men_men_n351_), .Y(men_men_n1159_));
  OAI210     u1131(.A0(men_men_n862_), .A1(men_men_n443_), .B0(men_men_n1159_), .Y(men_men_n1160_));
  NOi31      u1132(.An(m), .B(n), .C(f), .Y(men_men_n1161_));
  NA2        u1133(.A(men_men_n1161_), .B(men_men_n51_), .Y(men_men_n1162_));
  AN2        u1134(.A(e), .B(c), .Y(men_men_n1163_));
  NA2        u1135(.A(men_men_n1163_), .B(a), .Y(men_men_n1164_));
  OAI220     u1136(.A0(men_men_n1164_), .A1(men_men_n1162_), .B0(men_men_n928_), .B1(men_men_n448_), .Y(men_men_n1165_));
  NA2        u1137(.A(men_men_n530_), .B(l), .Y(men_men_n1166_));
  NOi31      u1138(.An(men_men_n905_), .B(men_men_n1079_), .C(men_men_n1166_), .Y(men_men_n1167_));
  NO4        u1139(.A(men_men_n1167_), .B(men_men_n1165_), .C(men_men_n1160_), .D(men_men_n1041_), .Y(men_men_n1168_));
  NO2        u1140(.A(men_men_n299_), .B(a), .Y(men_men_n1169_));
  INV        u1141(.A(men_men_n1086_), .Y(men_men_n1170_));
  NO2        u1142(.A(men_men_n1138_), .B(men_men_n505_), .Y(men_men_n1171_));
  NO2        u1143(.A(men_men_n89_), .B(u), .Y(men_men_n1172_));
  AOI210     u1144(.A0(men_men_n1172_), .A1(men_men_n1171_), .B0(men_men_n1121_), .Y(men_men_n1173_));
  OR2        u1145(.A(men_men_n1173_), .B(men_men_n1119_), .Y(men_men_n1174_));
  NA3        u1146(.A(men_men_n1174_), .B(men_men_n1170_), .C(men_men_n1168_), .Y(men_men_n1175_));
  NO4        u1147(.A(men_men_n1175_), .B(men_men_n1157_), .C(men_men_n864_), .D(men_men_n590_), .Y(men_men_n1176_));
  NA2        u1148(.A(c), .B(b), .Y(men_men_n1177_));
  NO2        u1149(.A(men_men_n735_), .B(men_men_n1177_), .Y(men_men_n1178_));
  OAI210     u1150(.A0(men_men_n903_), .A1(men_men_n876_), .B0(men_men_n436_), .Y(men_men_n1179_));
  OAI210     u1151(.A0(men_men_n1179_), .A1(men_men_n904_), .B0(men_men_n1178_), .Y(men_men_n1180_));
  NAi21      u1152(.An(men_men_n444_), .B(men_men_n1178_), .Y(men_men_n1181_));
  OAI210     u1153(.A0(men_men_n572_), .A1(men_men_n39_), .B0(men_men_n1169_), .Y(men_men_n1182_));
  NA2        u1154(.A(men_men_n1182_), .B(men_men_n1181_), .Y(men_men_n1183_));
  NA2        u1155(.A(men_men_n303_), .B(u), .Y(men_men_n1184_));
  NAi21      u1156(.An(f), .B(d), .Y(men_men_n1185_));
  NO2        u1157(.A(men_men_n1185_), .B(men_men_n1142_), .Y(men_men_n1186_));
  INV        u1158(.A(men_men_n1186_), .Y(men_men_n1187_));
  AOI210     u1159(.A0(men_men_n1184_), .A1(men_men_n309_), .B0(men_men_n1187_), .Y(men_men_n1188_));
  AOI210     u1160(.A0(men_men_n1188_), .A1(men_men_n117_), .B0(men_men_n1183_), .Y(men_men_n1189_));
  NA2        u1161(.A(men_men_n492_), .B(men_men_n491_), .Y(men_men_n1190_));
  NO2        u1162(.A(men_men_n191_), .B(men_men_n249_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n1191_), .B(m), .Y(men_men_n1192_));
  NA3        u1164(.A(men_men_n958_), .B(men_men_n1166_), .C(men_men_n172_), .Y(men_men_n1193_));
  OAI210     u1165(.A0(men_men_n1193_), .A1(men_men_n326_), .B0(men_men_n493_), .Y(men_men_n1194_));
  AOI210     u1166(.A0(men_men_n1194_), .A1(men_men_n1190_), .B0(men_men_n1192_), .Y(men_men_n1195_));
  NA2        u1167(.A(men_men_n585_), .B(men_men_n431_), .Y(men_men_n1196_));
  NA2        u1168(.A(men_men_n165_), .B(men_men_n33_), .Y(men_men_n1197_));
  AOI210     u1169(.A0(men_men_n1007_), .A1(men_men_n1197_), .B0(men_men_n225_), .Y(men_men_n1198_));
  NA2        u1170(.A(men_men_n1198_), .B(men_men_n1186_), .Y(men_men_n1199_));
  NO2        u1171(.A(men_men_n392_), .B(men_men_n391_), .Y(men_men_n1200_));
  AOI210     u1172(.A0(men_men_n1191_), .A1(men_men_n451_), .B0(men_men_n1001_), .Y(men_men_n1201_));
  NAi41      u1173(.An(men_men_n1200_), .B(men_men_n1201_), .C(men_men_n1199_), .D(men_men_n1196_), .Y(men_men_n1202_));
  NO2        u1174(.A(men_men_n1202_), .B(men_men_n1195_), .Y(men_men_n1203_));
  NA4        u1175(.A(men_men_n1203_), .B(men_men_n1189_), .C(men_men_n1180_), .D(men_men_n1176_), .Y(men00));
  AOI210     u1176(.A0(men_men_n312_), .A1(men_men_n225_), .B0(men_men_n292_), .Y(men_men_n1205_));
  NO2        u1177(.A(men_men_n1205_), .B(men_men_n603_), .Y(men_men_n1206_));
  AOI210     u1178(.A0(men_men_n938_), .A1(men_men_n985_), .B0(men_men_n1160_), .Y(men_men_n1207_));
  NO3        u1179(.A(men_men_n1135_), .B(men_men_n1001_), .C(men_men_n747_), .Y(men_men_n1208_));
  NA3        u1180(.A(men_men_n1208_), .B(men_men_n1207_), .C(men_men_n1043_), .Y(men_men_n1209_));
  NA2        u1181(.A(men_men_n532_), .B(f), .Y(men_men_n1210_));
  OAI210     u1182(.A0(men_men_n1050_), .A1(men_men_n40_), .B0(men_men_n675_), .Y(men_men_n1211_));
  NA3        u1183(.A(men_men_n1211_), .B(men_men_n271_), .C(n), .Y(men_men_n1212_));
  AOI210     u1184(.A0(men_men_n1212_), .A1(men_men_n1210_), .B0(men_men_n1090_), .Y(men_men_n1213_));
  NO4        u1185(.A(men_men_n1213_), .B(men_men_n1209_), .C(men_men_n1206_), .D(men_men_n1113_), .Y(men_men_n1214_));
  NA3        u1186(.A(men_men_n175_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1215_));
  NA3        u1187(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1216_));
  NOi31      u1188(.An(n), .B(m), .C(i), .Y(men_men_n1217_));
  NA3        u1189(.A(men_men_n1217_), .B(men_men_n678_), .C(men_men_n51_), .Y(men_men_n1218_));
  OAI210     u1190(.A0(men_men_n1216_), .A1(men_men_n1215_), .B0(men_men_n1218_), .Y(men_men_n1219_));
  INV        u1191(.A(men_men_n602_), .Y(men_men_n1220_));
  NO4        u1192(.A(men_men_n1220_), .B(men_men_n1219_), .C(men_men_n1200_), .D(men_men_n961_), .Y(men_men_n1221_));
  NO4        u1193(.A(men_men_n508_), .B(men_men_n374_), .C(men_men_n1177_), .D(men_men_n59_), .Y(men_men_n1222_));
  NA3        u1194(.A(men_men_n404_), .B(men_men_n232_), .C(u), .Y(men_men_n1223_));
  OA220      u1195(.A0(men_men_n1223_), .A1(men_men_n1216_), .B0(men_men_n405_), .B1(men_men_n139_), .Y(men_men_n1224_));
  NO2        u1196(.A(h), .B(u), .Y(men_men_n1225_));
  NA4        u1197(.A(men_men_n520_), .B(men_men_n489_), .C(men_men_n1225_), .D(men_men_n1078_), .Y(men_men_n1226_));
  OAI220     u1198(.A0(men_men_n550_), .A1(men_men_n622_), .B0(men_men_n94_), .B1(men_men_n93_), .Y(men_men_n1227_));
  NA2        u1199(.A(men_men_n1227_), .B(men_men_n558_), .Y(men_men_n1228_));
  AOI220     u1200(.A0(men_men_n333_), .A1(men_men_n260_), .B0(men_men_n186_), .B1(men_men_n154_), .Y(men_men_n1229_));
  NA4        u1201(.A(men_men_n1229_), .B(men_men_n1228_), .C(men_men_n1226_), .D(men_men_n1224_), .Y(men_men_n1230_));
  NO3        u1202(.A(men_men_n1230_), .B(men_men_n1222_), .C(men_men_n281_), .Y(men_men_n1231_));
  INV        u1203(.A(men_men_n338_), .Y(men_men_n1232_));
  AOI210     u1204(.A0(men_men_n260_), .A1(men_men_n365_), .B0(men_men_n604_), .Y(men_men_n1233_));
  NA3        u1205(.A(men_men_n1233_), .B(men_men_n1232_), .C(men_men_n160_), .Y(men_men_n1234_));
  NA3        u1206(.A(men_men_n188_), .B(men_men_n116_), .C(u), .Y(men_men_n1235_));
  NA3        u1207(.A(men_men_n489_), .B(men_men_n40_), .C(f), .Y(men_men_n1236_));
  NOi31      u1208(.An(men_men_n913_), .B(men_men_n1236_), .C(men_men_n1235_), .Y(men_men_n1237_));
  NAi31      u1209(.An(men_men_n195_), .B(men_men_n901_), .C(men_men_n489_), .Y(men_men_n1238_));
  NAi21      u1210(.An(men_men_n1237_), .B(men_men_n1238_), .Y(men_men_n1239_));
  NO2        u1211(.A(men_men_n291_), .B(men_men_n75_), .Y(men_men_n1240_));
  NO3        u1212(.A(men_men_n448_), .B(men_men_n872_), .C(n), .Y(men_men_n1241_));
  AOI210     u1213(.A0(men_men_n1241_), .A1(men_men_n1240_), .B0(men_men_n1128_), .Y(men_men_n1242_));
  NAi31      u1214(.An(men_men_n1093_), .B(men_men_n1242_), .C(men_men_n74_), .Y(men_men_n1243_));
  NO4        u1215(.A(men_men_n1243_), .B(men_men_n1239_), .C(men_men_n1234_), .D(men_men_n541_), .Y(men_men_n1244_));
  AN3        u1216(.A(men_men_n1244_), .B(men_men_n1231_), .C(men_men_n1221_), .Y(men_men_n1245_));
  NA2        u1217(.A(men_men_n558_), .B(men_men_n104_), .Y(men_men_n1246_));
  NA3        u1218(.A(men_men_n1161_), .B(men_men_n632_), .C(men_men_n488_), .Y(men_men_n1247_));
  NA4        u1219(.A(men_men_n1247_), .B(men_men_n586_), .C(men_men_n1246_), .D(men_men_n254_), .Y(men_men_n1248_));
  NA2        u1220(.A(men_men_n1154_), .B(men_men_n558_), .Y(men_men_n1249_));
  NA4        u1221(.A(men_men_n678_), .B(men_men_n216_), .C(men_men_n232_), .D(men_men_n169_), .Y(men_men_n1250_));
  NA2        u1222(.A(men_men_n1250_), .B(men_men_n1249_), .Y(men_men_n1251_));
  OAI210     u1223(.A0(men_men_n487_), .A1(men_men_n124_), .B0(men_men_n906_), .Y(men_men_n1252_));
  AOI220     u1224(.A0(men_men_n1252_), .A1(men_men_n1193_), .B0(men_men_n585_), .B1(men_men_n431_), .Y(men_men_n1253_));
  OR4        u1225(.A(men_men_n1090_), .B(men_men_n287_), .C(men_men_n234_), .D(e), .Y(men_men_n1254_));
  NA2        u1226(.A(n), .B(e), .Y(men_men_n1255_));
  NO2        u1227(.A(men_men_n1255_), .B(men_men_n152_), .Y(men_men_n1256_));
  NA2        u1228(.A(men_men_n1256_), .B(men_men_n289_), .Y(men_men_n1257_));
  OAI210     u1229(.A0(men_men_n375_), .A1(men_men_n327_), .B0(men_men_n468_), .Y(men_men_n1258_));
  NA4        u1230(.A(men_men_n1258_), .B(men_men_n1257_), .C(men_men_n1254_), .D(men_men_n1253_), .Y(men_men_n1259_));
  AOI210     u1231(.A0(men_men_n1256_), .A1(men_men_n892_), .B0(men_men_n863_), .Y(men_men_n1260_));
  AOI220     u1232(.A0(men_men_n997_), .A1(men_men_n601_), .B0(men_men_n678_), .B1(men_men_n257_), .Y(men_men_n1261_));
  NO2        u1233(.A(men_men_n68_), .B(h), .Y(men_men_n1262_));
  NO3        u1234(.A(men_men_n1090_), .B(men_men_n1088_), .C(men_men_n764_), .Y(men_men_n1263_));
  NO2        u1235(.A(men_men_n1125_), .B(men_men_n137_), .Y(men_men_n1264_));
  AN2        u1236(.A(men_men_n1264_), .B(men_men_n1140_), .Y(men_men_n1265_));
  OAI210     u1237(.A0(men_men_n1265_), .A1(men_men_n1263_), .B0(men_men_n1262_), .Y(men_men_n1266_));
  NA4        u1238(.A(men_men_n1266_), .B(men_men_n1261_), .C(men_men_n1260_), .D(men_men_n908_), .Y(men_men_n1267_));
  NO4        u1239(.A(men_men_n1267_), .B(men_men_n1259_), .C(men_men_n1251_), .D(men_men_n1248_), .Y(men_men_n1268_));
  NA2        u1240(.A(men_men_n877_), .B(men_men_n797_), .Y(men_men_n1269_));
  NA4        u1241(.A(men_men_n1269_), .B(men_men_n1268_), .C(men_men_n1245_), .D(men_men_n1214_), .Y(men01));
  AN2        u1242(.A(men_men_n1067_), .B(men_men_n1065_), .Y(men_men_n1271_));
  NO3        u1243(.A(men_men_n843_), .B(men_men_n835_), .C(men_men_n297_), .Y(men_men_n1272_));
  NO2        u1244(.A(men_men_n618_), .B(men_men_n306_), .Y(men_men_n1273_));
  OAI210     u1245(.A0(men_men_n1273_), .A1(men_men_n415_), .B0(i), .Y(men_men_n1274_));
  NA3        u1246(.A(men_men_n1274_), .B(men_men_n1272_), .C(men_men_n1271_), .Y(men_men_n1275_));
  NA2        u1247(.A(men_men_n614_), .B(men_men_n92_), .Y(men_men_n1276_));
  NA2        u1248(.A(men_men_n578_), .B(men_men_n286_), .Y(men_men_n1277_));
  NA2        u1249(.A(men_men_n1004_), .B(men_men_n1277_), .Y(men_men_n1278_));
  NA4        u1250(.A(men_men_n1278_), .B(men_men_n1276_), .C(men_men_n954_), .D(men_men_n350_), .Y(men_men_n1279_));
  NA2        u1251(.A(men_men_n45_), .B(f), .Y(men_men_n1280_));
  NA2        u1252(.A(men_men_n742_), .B(men_men_n99_), .Y(men_men_n1281_));
  OAI220     u1253(.A0(men_men_n1281_), .A1(men_men_n1280_), .B0(men_men_n371_), .B1(men_men_n301_), .Y(men_men_n1282_));
  OAI210     u1254(.A0(men_men_n822_), .A1(men_men_n628_), .B0(men_men_n1250_), .Y(men_men_n1283_));
  AOI210     u1255(.A0(men_men_n1282_), .A1(men_men_n663_), .B0(men_men_n1283_), .Y(men_men_n1284_));
  NA2        u1256(.A(men_men_n122_), .B(l), .Y(men_men_n1285_));
  OA220      u1257(.A0(men_men_n1285_), .A1(men_men_n611_), .B0(men_men_n691_), .B1(men_men_n389_), .Y(men_men_n1286_));
  NAi41      u1258(.An(men_men_n168_), .B(men_men_n1286_), .C(men_men_n1284_), .D(men_men_n937_), .Y(men_men_n1287_));
  NO2        u1259(.A(men_men_n707_), .B(men_men_n535_), .Y(men_men_n1288_));
  OR2        u1260(.A(men_men_n205_), .B(men_men_n203_), .Y(men_men_n1289_));
  NA3        u1261(.A(men_men_n1289_), .B(men_men_n1288_), .C(men_men_n142_), .Y(men_men_n1290_));
  NO4        u1262(.A(men_men_n1290_), .B(men_men_n1287_), .C(men_men_n1279_), .D(men_men_n1275_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n315_), .B(men_men_n553_), .Y(men_men_n1292_));
  NA2        u1264(.A(men_men_n561_), .B(men_men_n417_), .Y(men_men_n1293_));
  NA2        u1265(.A(men_men_n76_), .B(i), .Y(men_men_n1294_));
  AOI210     u1266(.A0(men_men_n617_), .A1(men_men_n611_), .B0(men_men_n1294_), .Y(men_men_n1295_));
  NOi21      u1267(.An(men_men_n587_), .B(men_men_n608_), .Y(men_men_n1296_));
  AOI210     u1268(.A0(men_men_n1296_), .A1(men_men_n1293_), .B0(men_men_n1295_), .Y(men_men_n1297_));
  AOI210     u1269(.A0(men_men_n214_), .A1(men_men_n91_), .B0(men_men_n224_), .Y(men_men_n1298_));
  OAI210     u1270(.A0(men_men_n850_), .A1(men_men_n449_), .B0(men_men_n1298_), .Y(men_men_n1299_));
  AN3        u1271(.A(m), .B(l), .C(k), .Y(men_men_n1300_));
  OAI210     u1272(.A0(men_men_n377_), .A1(men_men_n34_), .B0(men_men_n1300_), .Y(men_men_n1301_));
  NA2        u1273(.A(men_men_n213_), .B(men_men_n34_), .Y(men_men_n1302_));
  AO210      u1274(.A0(men_men_n1302_), .A1(men_men_n1301_), .B0(men_men_n349_), .Y(men_men_n1303_));
  NA4        u1275(.A(men_men_n1303_), .B(men_men_n1299_), .C(men_men_n1297_), .D(men_men_n1292_), .Y(men_men_n1304_));
  INV        u1276(.A(men_men_n626_), .Y(men_men_n1305_));
  OAI210     u1277(.A0(men_men_n1285_), .A1(men_men_n620_), .B0(men_men_n1305_), .Y(men_men_n1306_));
  NA2        u1278(.A(men_men_n296_), .B(men_men_n205_), .Y(men_men_n1307_));
  OAI210     u1279(.A0(men_men_n1307_), .A1(men_men_n406_), .B0(men_men_n696_), .Y(men_men_n1308_));
  NO3        u1280(.A(men_men_n862_), .B(men_men_n214_), .C(men_men_n429_), .Y(men_men_n1309_));
  NO2        u1281(.A(men_men_n1309_), .B(men_men_n1001_), .Y(men_men_n1310_));
  OAI210     u1282(.A0(men_men_n1282_), .A1(men_men_n343_), .B0(men_men_n708_), .Y(men_men_n1311_));
  NA4        u1283(.A(men_men_n1311_), .B(men_men_n1310_), .C(men_men_n1308_), .D(men_men_n825_), .Y(men_men_n1312_));
  NO3        u1284(.A(men_men_n1312_), .B(men_men_n1306_), .C(men_men_n1304_), .Y(men_men_n1313_));
  NA3        u1285(.A(men_men_n629_), .B(men_men_n29_), .C(f), .Y(men_men_n1314_));
  NO2        u1286(.A(men_men_n1314_), .B(men_men_n214_), .Y(men_men_n1315_));
  AOI210     u1287(.A0(men_men_n527_), .A1(men_men_n58_), .B0(men_men_n1315_), .Y(men_men_n1316_));
  OR3        u1288(.A(men_men_n1281_), .B(men_men_n630_), .C(men_men_n1280_), .Y(men_men_n1317_));
  NA3        u1289(.A(men_men_n778_), .B(men_men_n76_), .C(i), .Y(men_men_n1318_));
  NO2        u1290(.A(men_men_n1318_), .B(men_men_n1022_), .Y(men_men_n1319_));
  NO2        u1291(.A(men_men_n217_), .B(men_men_n115_), .Y(men_men_n1320_));
  NO3        u1292(.A(men_men_n1320_), .B(men_men_n1319_), .C(men_men_n1219_), .Y(men_men_n1321_));
  NA4        u1293(.A(men_men_n1321_), .B(men_men_n1317_), .C(men_men_n1316_), .D(men_men_n796_), .Y(men_men_n1322_));
  NO2        u1294(.A(men_men_n1011_), .B(men_men_n244_), .Y(men_men_n1323_));
  NO2        u1295(.A(men_men_n1012_), .B(men_men_n580_), .Y(men_men_n1324_));
  OAI210     u1296(.A0(men_men_n1324_), .A1(men_men_n1323_), .B0(men_men_n358_), .Y(men_men_n1325_));
  NO3        u1297(.A(men_men_n81_), .B(men_men_n313_), .C(men_men_n45_), .Y(men_men_n1326_));
  NA2        u1298(.A(men_men_n1326_), .B(men_men_n577_), .Y(men_men_n1327_));
  NA2        u1299(.A(men_men_n1327_), .B(men_men_n702_), .Y(men_men_n1328_));
  OR2        u1300(.A(men_men_n1223_), .B(men_men_n1216_), .Y(men_men_n1329_));
  NO2        u1301(.A(men_men_n389_), .B(men_men_n73_), .Y(men_men_n1330_));
  AOI210     u1302(.A0(men_men_n769_), .A1(men_men_n643_), .B0(men_men_n1330_), .Y(men_men_n1331_));
  NA2        u1303(.A(men_men_n1326_), .B(men_men_n853_), .Y(men_men_n1332_));
  NA4        u1304(.A(men_men_n1332_), .B(men_men_n1331_), .C(men_men_n1329_), .D(men_men_n407_), .Y(men_men_n1333_));
  NOi41      u1305(.An(men_men_n1325_), .B(men_men_n1333_), .C(men_men_n1328_), .D(men_men_n1322_), .Y(men_men_n1334_));
  NO2        u1306(.A(men_men_n136_), .B(men_men_n45_), .Y(men_men_n1335_));
  NO2        u1307(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1336_));
  AO220      u1308(.A0(men_men_n1336_), .A1(men_men_n649_), .B0(men_men_n1335_), .B1(men_men_n740_), .Y(men_men_n1337_));
  NA2        u1309(.A(men_men_n1337_), .B(men_men_n358_), .Y(men_men_n1338_));
  INV        u1310(.A(men_men_n139_), .Y(men_men_n1339_));
  NO3        u1311(.A(men_men_n1138_), .B(men_men_n185_), .C(men_men_n89_), .Y(men_men_n1340_));
  NA2        u1312(.A(men_men_n1340_), .B(men_men_n1339_), .Y(men_men_n1341_));
  NA2        u1313(.A(men_men_n1341_), .B(men_men_n1338_), .Y(men_men_n1342_));
  NO2        u1314(.A(men_men_n640_), .B(men_men_n639_), .Y(men_men_n1343_));
  NO4        u1315(.A(men_men_n1138_), .B(men_men_n1343_), .C(men_men_n183_), .D(men_men_n89_), .Y(men_men_n1344_));
  NO3        u1316(.A(men_men_n1344_), .B(men_men_n1342_), .C(men_men_n667_), .Y(men_men_n1345_));
  NA4        u1317(.A(men_men_n1345_), .B(men_men_n1334_), .C(men_men_n1313_), .D(men_men_n1291_), .Y(men06));
  NO2        u1318(.A(men_men_n430_), .B(men_men_n584_), .Y(men_men_n1347_));
  NO2        u1319(.A(men_men_n771_), .B(i), .Y(men_men_n1348_));
  OAI210     u1320(.A0(men_men_n1348_), .A1(men_men_n282_), .B0(men_men_n1347_), .Y(men_men_n1349_));
  NO2        u1321(.A(men_men_n236_), .B(men_men_n106_), .Y(men_men_n1350_));
  OAI210     u1322(.A0(men_men_n1350_), .A1(men_men_n1340_), .B0(men_men_n403_), .Y(men_men_n1351_));
  NO3        u1323(.A(men_men_n624_), .B(men_men_n848_), .C(men_men_n627_), .Y(men_men_n1352_));
  OR2        u1324(.A(men_men_n1352_), .B(men_men_n928_), .Y(men_men_n1353_));
  NA4        u1325(.A(men_men_n1353_), .B(men_men_n1351_), .C(men_men_n1349_), .D(men_men_n1325_), .Y(men_men_n1354_));
  NO3        u1326(.A(men_men_n1354_), .B(men_men_n1328_), .C(men_men_n270_), .Y(men_men_n1355_));
  NO2        u1327(.A(men_men_n313_), .B(men_men_n45_), .Y(men_men_n1356_));
  AOI210     u1328(.A0(men_men_n1356_), .A1(men_men_n577_), .B0(men_men_n1323_), .Y(men_men_n1357_));
  AOI210     u1329(.A0(men_men_n1356_), .A1(men_men_n581_), .B0(men_men_n1337_), .Y(men_men_n1358_));
  AOI210     u1330(.A0(men_men_n1358_), .A1(men_men_n1357_), .B0(men_men_n355_), .Y(men_men_n1359_));
  OAI210     u1331(.A0(men_men_n91_), .A1(men_men_n40_), .B0(men_men_n706_), .Y(men_men_n1360_));
  NA2        u1332(.A(men_men_n1360_), .B(men_men_n671_), .Y(men_men_n1361_));
  NO2        u1333(.A(men_men_n538_), .B(men_men_n180_), .Y(men_men_n1362_));
  NOi21      u1334(.An(men_men_n141_), .B(men_men_n45_), .Y(men_men_n1363_));
  NO2        u1335(.A(men_men_n633_), .B(men_men_n1162_), .Y(men_men_n1364_));
  OAI210     u1336(.A0(men_men_n482_), .A1(men_men_n261_), .B0(men_men_n948_), .Y(men_men_n1365_));
  NO4        u1337(.A(men_men_n1365_), .B(men_men_n1364_), .C(men_men_n1363_), .D(men_men_n1362_), .Y(men_men_n1366_));
  OR2        u1338(.A(men_men_n625_), .B(men_men_n623_), .Y(men_men_n1367_));
  INV        u1339(.A(men_men_n1367_), .Y(men_men_n1368_));
  NA3        u1340(.A(men_men_n1368_), .B(men_men_n1366_), .C(men_men_n1361_), .Y(men_men_n1369_));
  NO2        u1341(.A(men_men_n787_), .B(men_men_n387_), .Y(men_men_n1370_));
  NO3        u1342(.A(men_men_n708_), .B(men_men_n798_), .C(men_men_n663_), .Y(men_men_n1371_));
  NOi21      u1343(.An(men_men_n1370_), .B(men_men_n1371_), .Y(men_men_n1372_));
  AN2        u1344(.A(men_men_n997_), .B(men_men_n674_), .Y(men_men_n1373_));
  NO4        u1345(.A(men_men_n1373_), .B(men_men_n1372_), .C(men_men_n1369_), .D(men_men_n1359_), .Y(men_men_n1374_));
  NO2        u1346(.A(men_men_n842_), .B(men_men_n293_), .Y(men_men_n1375_));
  OAI220     u1347(.A0(men_men_n771_), .A1(men_men_n47_), .B0(men_men_n236_), .B1(men_men_n642_), .Y(men_men_n1376_));
  OAI210     u1348(.A0(men_men_n293_), .A1(c), .B0(men_men_n670_), .Y(men_men_n1377_));
  AOI220     u1349(.A0(men_men_n1377_), .A1(men_men_n1376_), .B0(men_men_n1375_), .B1(men_men_n282_), .Y(men_men_n1378_));
  NO3        u1350(.A(men_men_n256_), .B(men_men_n106_), .C(men_men_n299_), .Y(men_men_n1379_));
  OAI220     u1351(.A0(men_men_n732_), .A1(men_men_n261_), .B0(men_men_n534_), .B1(men_men_n538_), .Y(men_men_n1380_));
  OAI210     u1352(.A0(l), .A1(i), .B0(k), .Y(men_men_n1381_));
  NO3        u1353(.A(men_men_n1381_), .B(men_men_n622_), .C(j), .Y(men_men_n1382_));
  NOi21      u1354(.An(men_men_n1382_), .B(men_men_n700_), .Y(men_men_n1383_));
  NO4        u1355(.A(men_men_n1383_), .B(men_men_n1380_), .C(men_men_n1379_), .D(men_men_n1165_), .Y(men_men_n1384_));
  NA3        u1356(.A(men_men_n1384_), .B(men_men_n1378_), .C(men_men_n1261_), .Y(men_men_n1385_));
  NOi31      u1357(.An(men_men_n1352_), .B(men_men_n486_), .C(men_men_n416_), .Y(men_men_n1386_));
  OR3        u1358(.A(men_men_n1386_), .B(men_men_n822_), .C(men_men_n564_), .Y(men_men_n1387_));
  OR3        u1359(.A(men_men_n391_), .B(men_men_n236_), .C(men_men_n642_), .Y(men_men_n1388_));
  AOI210     u1360(.A0(men_men_n596_), .A1(men_men_n468_), .B0(men_men_n393_), .Y(men_men_n1389_));
  NA2        u1361(.A(men_men_n1382_), .B(men_men_n829_), .Y(men_men_n1390_));
  NA4        u1362(.A(men_men_n1390_), .B(men_men_n1389_), .C(men_men_n1388_), .D(men_men_n1387_), .Y(men_men_n1391_));
  NA2        u1363(.A(men_men_n1370_), .B(men_men_n797_), .Y(men_men_n1392_));
  AN2        u1364(.A(men_men_n970_), .B(men_men_n969_), .Y(men_men_n1393_));
  NO4        u1365(.A(men_men_n1393_), .B(men_men_n918_), .C(men_men_n523_), .D(men_men_n502_), .Y(men_men_n1394_));
  NA3        u1366(.A(men_men_n1394_), .B(men_men_n1392_), .C(men_men_n1332_), .Y(men_men_n1395_));
  NAi21      u1367(.An(j), .B(i), .Y(men_men_n1396_));
  NO4        u1368(.A(men_men_n1343_), .B(men_men_n1396_), .C(men_men_n462_), .D(men_men_n247_), .Y(men_men_n1397_));
  NO4        u1369(.A(men_men_n1397_), .B(men_men_n1395_), .C(men_men_n1391_), .D(men_men_n1385_), .Y(men_men_n1398_));
  NA4        u1370(.A(men_men_n1398_), .B(men_men_n1374_), .C(men_men_n1355_), .D(men_men_n1345_), .Y(men07));
  NOi21      u1371(.An(j), .B(k), .Y(men_men_n1400_));
  NA4        u1372(.A(men_men_n188_), .B(men_men_n112_), .C(men_men_n1400_), .D(f), .Y(men_men_n1401_));
  NAi32      u1373(.An(m), .Bn(b), .C(n), .Y(men_men_n1402_));
  NO3        u1374(.A(men_men_n1402_), .B(u), .C(f), .Y(men_men_n1403_));
  OAI210     u1375(.A0(men_men_n337_), .A1(men_men_n504_), .B0(men_men_n1403_), .Y(men_men_n1404_));
  NAi21      u1376(.An(f), .B(c), .Y(men_men_n1405_));
  OR2        u1377(.A(e), .B(d), .Y(men_men_n1406_));
  OAI220     u1378(.A0(men_men_n1406_), .A1(men_men_n1405_), .B0(men_men_n655_), .B1(men_men_n339_), .Y(men_men_n1407_));
  NA3        u1379(.A(men_men_n1407_), .B(men_men_n1102_), .C(men_men_n188_), .Y(men_men_n1408_));
  NOi31      u1380(.An(n), .B(m), .C(b), .Y(men_men_n1409_));
  NO3        u1381(.A(men_men_n137_), .B(men_men_n470_), .C(h), .Y(men_men_n1410_));
  NA3        u1382(.A(men_men_n1408_), .B(men_men_n1404_), .C(men_men_n1401_), .Y(men_men_n1411_));
  NOi41      u1383(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1412_));
  NA3        u1384(.A(men_men_n1412_), .B(men_men_n910_), .C(men_men_n432_), .Y(men_men_n1413_));
  NO2        u1385(.A(men_men_n1413_), .B(men_men_n56_), .Y(men_men_n1414_));
  NA2        u1386(.A(men_men_n1140_), .B(men_men_n232_), .Y(men_men_n1415_));
  NO2        u1387(.A(men_men_n1415_), .B(men_men_n61_), .Y(men_men_n1416_));
  NO2        u1388(.A(k), .B(i), .Y(men_men_n1417_));
  NA3        u1389(.A(men_men_n1417_), .B(men_men_n936_), .C(men_men_n188_), .Y(men_men_n1418_));
  NA2        u1390(.A(men_men_n89_), .B(men_men_n45_), .Y(men_men_n1419_));
  NO2        u1391(.A(men_men_n1096_), .B(men_men_n462_), .Y(men_men_n1420_));
  NA3        u1392(.A(men_men_n1420_), .B(men_men_n1419_), .C(men_men_n225_), .Y(men_men_n1421_));
  NO2        u1393(.A(men_men_n1110_), .B(men_men_n321_), .Y(men_men_n1422_));
  NA2        u1394(.A(men_men_n565_), .B(men_men_n82_), .Y(men_men_n1423_));
  NA2        u1395(.A(men_men_n1262_), .B(men_men_n307_), .Y(men_men_n1424_));
  NA4        u1396(.A(men_men_n1424_), .B(men_men_n1423_), .C(men_men_n1421_), .D(men_men_n1418_), .Y(men_men_n1425_));
  NO4        u1397(.A(men_men_n1425_), .B(men_men_n1416_), .C(men_men_n1414_), .D(men_men_n1411_), .Y(men_men_n1426_));
  NO3        u1398(.A(e), .B(d), .C(c), .Y(men_men_n1427_));
  AOI210     u1399(.A0(men_men_n1117_), .A1(men_men_n225_), .B0(men_men_n1427_), .Y(men_men_n1428_));
  OAI210     u1400(.A0(men_men_n137_), .A1(men_men_n225_), .B0(men_men_n631_), .Y(men_men_n1429_));
  NA2        u1401(.A(men_men_n1429_), .B(men_men_n1427_), .Y(men_men_n1430_));
  NO2        u1402(.A(men_men_n1430_), .B(men_men_n1428_), .Y(men_men_n1431_));
  OR2        u1403(.A(h), .B(f), .Y(men_men_n1432_));
  NO3        u1404(.A(n), .B(m), .C(i), .Y(men_men_n1433_));
  OAI210     u1405(.A0(men_men_n1163_), .A1(men_men_n163_), .B0(men_men_n1433_), .Y(men_men_n1434_));
  NO2        u1406(.A(i), .B(u), .Y(men_men_n1435_));
  OR3        u1407(.A(men_men_n1435_), .B(men_men_n1402_), .C(men_men_n72_), .Y(men_men_n1436_));
  OAI220     u1408(.A0(men_men_n1436_), .A1(men_men_n504_), .B0(men_men_n1434_), .B1(men_men_n1432_), .Y(men_men_n1437_));
  NA3        u1409(.A(men_men_n729_), .B(men_men_n716_), .C(men_men_n116_), .Y(men_men_n1438_));
  NA3        u1410(.A(men_men_n1409_), .B(men_men_n1105_), .C(men_men_n704_), .Y(men_men_n1439_));
  AOI210     u1411(.A0(men_men_n1439_), .A1(men_men_n1438_), .B0(men_men_n45_), .Y(men_men_n1440_));
  NO2        u1412(.A(l), .B(k), .Y(men_men_n1441_));
  NOi41      u1413(.An(men_men_n570_), .B(men_men_n1441_), .C(men_men_n499_), .D(men_men_n462_), .Y(men_men_n1442_));
  NO3        u1414(.A(men_men_n462_), .B(d), .C(c), .Y(men_men_n1443_));
  NO4        u1415(.A(men_men_n1442_), .B(men_men_n1440_), .C(men_men_n1437_), .D(men_men_n1431_), .Y(men_men_n1444_));
  NO2        u1416(.A(men_men_n153_), .B(h), .Y(men_men_n1445_));
  NO2        u1417(.A(men_men_n1120_), .B(l), .Y(men_men_n1446_));
  NO2        u1418(.A(u), .B(c), .Y(men_men_n1447_));
  NA3        u1419(.A(men_men_n1447_), .B(men_men_n147_), .C(men_men_n196_), .Y(men_men_n1448_));
  NO2        u1420(.A(men_men_n1448_), .B(men_men_n1446_), .Y(men_men_n1449_));
  NA2        u1421(.A(men_men_n1449_), .B(men_men_n188_), .Y(men_men_n1450_));
  NO2        u1422(.A(men_men_n473_), .B(a), .Y(men_men_n1451_));
  NA3        u1423(.A(men_men_n1451_), .B(k), .C(men_men_n117_), .Y(men_men_n1452_));
  NO2        u1424(.A(i), .B(h), .Y(men_men_n1453_));
  NA2        u1425(.A(men_men_n1453_), .B(men_men_n232_), .Y(men_men_n1454_));
  AOI210     u1426(.A0(men_men_n1185_), .A1(h), .B0(men_men_n437_), .Y(men_men_n1455_));
  NA2        u1427(.A(men_men_n143_), .B(men_men_n232_), .Y(men_men_n1456_));
  AOI210     u1428(.A0(men_men_n271_), .A1(men_men_n120_), .B0(men_men_n553_), .Y(men_men_n1457_));
  OAI220     u1429(.A0(men_men_n1457_), .A1(men_men_n1454_), .B0(men_men_n1456_), .B1(men_men_n1455_), .Y(men_men_n1458_));
  NO2        u1430(.A(men_men_n794_), .B(men_men_n197_), .Y(men_men_n1459_));
  NOi31      u1431(.An(m), .B(n), .C(b), .Y(men_men_n1460_));
  NOi31      u1432(.An(f), .B(d), .C(c), .Y(men_men_n1461_));
  NA2        u1433(.A(men_men_n1461_), .B(men_men_n1460_), .Y(men_men_n1462_));
  INV        u1434(.A(men_men_n1462_), .Y(men_men_n1463_));
  NO3        u1435(.A(men_men_n1463_), .B(men_men_n1459_), .C(men_men_n1458_), .Y(men_men_n1464_));
  NA2        u1436(.A(men_men_n1131_), .B(men_men_n489_), .Y(men_men_n1465_));
  NO4        u1437(.A(men_men_n1465_), .B(men_men_n1105_), .C(men_men_n462_), .D(men_men_n45_), .Y(men_men_n1466_));
  OAI210     u1438(.A0(men_men_n191_), .A1(men_men_n549_), .B0(men_men_n1106_), .Y(men_men_n1467_));
  NO3        u1439(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1468_));
  INV        u1440(.A(men_men_n1467_), .Y(men_men_n1469_));
  NO2        u1441(.A(men_men_n1469_), .B(men_men_n1466_), .Y(men_men_n1470_));
  AN4        u1442(.A(men_men_n1470_), .B(men_men_n1464_), .C(men_men_n1452_), .D(men_men_n1450_), .Y(men_men_n1471_));
  NA2        u1443(.A(men_men_n1409_), .B(men_men_n400_), .Y(men_men_n1472_));
  NO2        u1444(.A(men_men_n1472_), .B(men_men_n1087_), .Y(men_men_n1473_));
  NA2        u1445(.A(men_men_n1443_), .B(men_men_n226_), .Y(men_men_n1474_));
  NO2        u1446(.A(men_men_n197_), .B(b), .Y(men_men_n1475_));
  AOI220     u1447(.A0(men_men_n1217_), .A1(men_men_n1475_), .B0(men_men_n1139_), .B1(men_men_n1465_), .Y(men_men_n1476_));
  NO2        u1448(.A(i), .B(men_men_n224_), .Y(men_men_n1477_));
  NA4        u1449(.A(men_men_n1191_), .B(men_men_n1477_), .C(men_men_n107_), .D(m), .Y(men_men_n1478_));
  NAi41      u1450(.An(men_men_n1473_), .B(men_men_n1478_), .C(men_men_n1476_), .D(men_men_n1474_), .Y(men_men_n1479_));
  NO4        u1451(.A(men_men_n137_), .B(u), .C(f), .D(e), .Y(men_men_n1480_));
  NA3        u1452(.A(men_men_n1417_), .B(men_men_n308_), .C(h), .Y(men_men_n1481_));
  NA2        u1453(.A(men_men_n204_), .B(men_men_n101_), .Y(men_men_n1482_));
  OR2        u1454(.A(e), .B(a), .Y(men_men_n1483_));
  NO2        u1455(.A(men_men_n1406_), .B(men_men_n1405_), .Y(men_men_n1484_));
  AOI210     u1456(.A0(men_men_n30_), .A1(h), .B0(men_men_n1484_), .Y(men_men_n1485_));
  NO2        u1457(.A(men_men_n1485_), .B(men_men_n1127_), .Y(men_men_n1486_));
  NA2        u1458(.A(men_men_n1412_), .B(men_men_n1441_), .Y(men_men_n1487_));
  INV        u1459(.A(men_men_n1487_), .Y(men_men_n1488_));
  OR3        u1460(.A(men_men_n564_), .B(men_men_n563_), .C(men_men_n116_), .Y(men_men_n1489_));
  NA2        u1461(.A(men_men_n1161_), .B(men_men_n429_), .Y(men_men_n1490_));
  OAI220     u1462(.A0(men_men_n1490_), .A1(men_men_n458_), .B0(men_men_n1489_), .B1(men_men_n313_), .Y(men_men_n1491_));
  AO210      u1463(.A0(men_men_n1491_), .A1(men_men_n120_), .B0(men_men_n1488_), .Y(men_men_n1492_));
  NO3        u1464(.A(men_men_n1492_), .B(men_men_n1486_), .C(men_men_n1479_), .Y(men_men_n1493_));
  NA4        u1465(.A(men_men_n1493_), .B(men_men_n1471_), .C(men_men_n1444_), .D(men_men_n1426_), .Y(men_men_n1494_));
  NO2        u1466(.A(men_men_n1177_), .B(men_men_n114_), .Y(men_men_n1495_));
  NA2        u1467(.A(men_men_n400_), .B(men_men_n56_), .Y(men_men_n1496_));
  NA2        u1468(.A(men_men_n226_), .B(men_men_n188_), .Y(men_men_n1497_));
  AOI210     u1469(.A0(men_men_n1497_), .A1(men_men_n1235_), .B0(men_men_n1496_), .Y(men_men_n1498_));
  NO2        u1470(.A(men_men_n412_), .B(j), .Y(men_men_n1499_));
  NA3        u1471(.A(men_men_n1468_), .B(men_men_n1406_), .C(men_men_n1161_), .Y(men_men_n1500_));
  NAi41      u1472(.An(men_men_n1453_), .B(men_men_n1118_), .C(men_men_n176_), .D(men_men_n156_), .Y(men_men_n1501_));
  NA2        u1473(.A(men_men_n1501_), .B(men_men_n1500_), .Y(men_men_n1502_));
  NA3        u1474(.A(u), .B(men_men_n1499_), .C(men_men_n165_), .Y(men_men_n1503_));
  INV        u1475(.A(men_men_n1503_), .Y(men_men_n1504_));
  NO3        u1476(.A(men_men_n787_), .B(men_men_n183_), .C(men_men_n432_), .Y(men_men_n1505_));
  NO3        u1477(.A(men_men_n1505_), .B(men_men_n1504_), .C(men_men_n1502_), .Y(men_men_n1506_));
  NO3        u1478(.A(men_men_n1127_), .B(men_men_n608_), .C(u), .Y(men_men_n1507_));
  NOi21      u1479(.An(men_men_n1497_), .B(men_men_n1507_), .Y(men_men_n1508_));
  AOI210     u1480(.A0(men_men_n1508_), .A1(men_men_n1482_), .B0(men_men_n1096_), .Y(men_men_n1509_));
  OR2        u1481(.A(n), .B(i), .Y(men_men_n1510_));
  OAI210     u1482(.A0(men_men_n1510_), .A1(men_men_n1117_), .B0(men_men_n49_), .Y(men_men_n1511_));
  AOI220     u1483(.A0(men_men_n1511_), .A1(men_men_n1225_), .B0(men_men_n867_), .B1(men_men_n204_), .Y(men_men_n1512_));
  INV        u1484(.A(men_men_n1512_), .Y(men_men_n1513_));
  NO2        u1485(.A(men_men_n236_), .B(k), .Y(men_men_n1514_));
  NO2        u1486(.A(men_men_n1513_), .B(men_men_n1509_), .Y(men_men_n1515_));
  NO2        u1487(.A(men_men_n49_), .B(men_men_n608_), .Y(men_men_n1516_));
  NO3        u1488(.A(men_men_n1142_), .B(men_men_n1406_), .C(men_men_n49_), .Y(men_men_n1517_));
  NA2        u1489(.A(men_men_n1143_), .B(men_men_n1516_), .Y(men_men_n1518_));
  NO2        u1490(.A(men_men_n1127_), .B(h), .Y(men_men_n1519_));
  NA3        u1491(.A(men_men_n1519_), .B(d), .C(men_men_n1088_), .Y(men_men_n1520_));
  OAI220     u1492(.A0(men_men_n1520_), .A1(c), .B0(men_men_n1518_), .B1(j), .Y(men_men_n1521_));
  NA3        u1493(.A(men_men_n1495_), .B(men_men_n489_), .C(f), .Y(men_men_n1522_));
  NA2        u1494(.A(men_men_n188_), .B(men_men_n116_), .Y(men_men_n1523_));
  NO2        u1495(.A(men_men_n1400_), .B(men_men_n42_), .Y(men_men_n1524_));
  AOI210     u1496(.A0(men_men_n117_), .A1(men_men_n40_), .B0(men_men_n1524_), .Y(men_men_n1525_));
  NO2        u1497(.A(men_men_n1525_), .B(men_men_n1522_), .Y(men_men_n1526_));
  AOI210     u1498(.A0(men_men_n549_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1527_));
  NA2        u1499(.A(men_men_n1527_), .B(men_men_n1451_), .Y(men_men_n1528_));
  NO2        u1500(.A(men_men_n1396_), .B(men_men_n183_), .Y(men_men_n1529_));
  NOi21      u1501(.An(d), .B(f), .Y(men_men_n1530_));
  NO3        u1502(.A(men_men_n1461_), .B(men_men_n1530_), .C(men_men_n40_), .Y(men_men_n1531_));
  NA2        u1503(.A(men_men_n1531_), .B(men_men_n1529_), .Y(men_men_n1532_));
  NO2        u1504(.A(men_men_n1406_), .B(f), .Y(men_men_n1533_));
  NA2        u1505(.A(men_men_n1451_), .B(men_men_n1524_), .Y(men_men_n1534_));
  NO2        u1506(.A(men_men_n313_), .B(c), .Y(men_men_n1535_));
  NA2        u1507(.A(men_men_n1535_), .B(men_men_n565_), .Y(men_men_n1536_));
  NA4        u1508(.A(men_men_n1536_), .B(men_men_n1534_), .C(men_men_n1532_), .D(men_men_n1528_), .Y(men_men_n1537_));
  NO3        u1509(.A(men_men_n1537_), .B(men_men_n1526_), .C(men_men_n1521_), .Y(men_men_n1538_));
  NA4        u1510(.A(men_men_n1538_), .B(men_men_n1515_), .C(men_men_n1506_), .D(men_men_n1621_), .Y(men_men_n1539_));
  NO3        u1511(.A(men_men_n1131_), .B(men_men_n1117_), .C(men_men_n40_), .Y(men_men_n1540_));
  OAI220     u1512(.A0(men_men_n489_), .A1(men_men_n313_), .B0(men_men_n136_), .B1(men_men_n59_), .Y(men_men_n1541_));
  OAI210     u1513(.A0(men_men_n1541_), .A1(men_men_n1540_), .B0(men_men_n1422_), .Y(men_men_n1542_));
  OAI210     u1514(.A0(men_men_n1480_), .A1(men_men_n1409_), .B0(men_men_n925_), .Y(men_men_n1543_));
  OAI220     u1515(.A0(men_men_n1084_), .A1(men_men_n137_), .B0(men_men_n697_), .B1(men_men_n183_), .Y(men_men_n1544_));
  NA2        u1516(.A(men_men_n1544_), .B(men_men_n648_), .Y(men_men_n1545_));
  NA3        u1517(.A(men_men_n1545_), .B(men_men_n1543_), .C(men_men_n1542_), .Y(men_men_n1546_));
  NA2        u1518(.A(men_men_n1447_), .B(men_men_n1530_), .Y(men_men_n1547_));
  NO2        u1519(.A(men_men_n1547_), .B(m), .Y(men_men_n1548_));
  NA3        u1520(.A(men_men_n1140_), .B(men_men_n112_), .C(men_men_n232_), .Y(men_men_n1549_));
  OAI220     u1521(.A0(men_men_n157_), .A1(men_men_n190_), .B0(men_men_n470_), .B1(u), .Y(men_men_n1550_));
  OAI210     u1522(.A0(men_men_n1550_), .A1(men_men_n114_), .B0(men_men_n1460_), .Y(men_men_n1551_));
  NA2        u1523(.A(men_men_n1551_), .B(men_men_n1549_), .Y(men_men_n1552_));
  NO3        u1524(.A(men_men_n1552_), .B(men_men_n1548_), .C(men_men_n1546_), .Y(men_men_n1553_));
  NO2        u1525(.A(men_men_n1405_), .B(e), .Y(men_men_n1554_));
  NA2        u1526(.A(men_men_n1554_), .B(men_men_n427_), .Y(men_men_n1555_));
  OAI210     u1527(.A0(men_men_n1533_), .A1(men_men_n1172_), .B0(men_men_n659_), .Y(men_men_n1556_));
  OR3        u1528(.A(men_men_n1514_), .B(men_men_n1262_), .C(men_men_n137_), .Y(men_men_n1557_));
  OAI220     u1529(.A0(men_men_n1557_), .A1(men_men_n1555_), .B0(men_men_n1556_), .B1(men_men_n464_), .Y(men_men_n1558_));
  NO3        u1530(.A(men_men_n1489_), .B(men_men_n371_), .C(a), .Y(men_men_n1559_));
  NO2        u1531(.A(men_men_n1559_), .B(men_men_n1558_), .Y(men_men_n1560_));
  NO2        u1532(.A(men_men_n190_), .B(c), .Y(men_men_n1561_));
  OAI210     u1533(.A0(men_men_n1561_), .A1(men_men_n1554_), .B0(men_men_n188_), .Y(men_men_n1562_));
  AOI220     u1534(.A0(men_men_n1562_), .A1(men_men_n1119_), .B0(men_men_n555_), .B1(men_men_n387_), .Y(men_men_n1563_));
  NA2        u1535(.A(men_men_n563_), .B(u), .Y(men_men_n1564_));
  AOI210     u1536(.A0(men_men_n1564_), .A1(men_men_n1443_), .B0(men_men_n1517_), .Y(men_men_n1565_));
  NO2        u1537(.A(men_men_n1483_), .B(f), .Y(men_men_n1566_));
  NO2        u1538(.A(men_men_n1565_), .B(men_men_n224_), .Y(men_men_n1567_));
  AOI210     u1539(.A0(men_men_n941_), .A1(men_men_n439_), .B0(men_men_n108_), .Y(men_men_n1568_));
  OR2        u1540(.A(men_men_n1568_), .B(men_men_n563_), .Y(men_men_n1569_));
  NA2        u1541(.A(men_men_n1566_), .B(men_men_n1419_), .Y(men_men_n1570_));
  OAI220     u1542(.A0(men_men_n1570_), .A1(men_men_n49_), .B0(men_men_n1569_), .B1(men_men_n183_), .Y(men_men_n1571_));
  NA4        u1543(.A(men_men_n1140_), .B(men_men_n1137_), .C(men_men_n232_), .D(men_men_n68_), .Y(men_men_n1572_));
  NA2        u1544(.A(men_men_n1410_), .B(men_men_n191_), .Y(men_men_n1573_));
  NO2        u1545(.A(men_men_n49_), .B(l), .Y(men_men_n1574_));
  OAI210     u1546(.A0(men_men_n1483_), .A1(men_men_n902_), .B0(men_men_n504_), .Y(men_men_n1575_));
  OAI210     u1547(.A0(men_men_n1575_), .A1(men_men_n1143_), .B0(men_men_n1574_), .Y(men_men_n1576_));
  NO2        u1548(.A(men_men_n266_), .B(u), .Y(men_men_n1577_));
  NO2        u1549(.A(m), .B(i), .Y(men_men_n1578_));
  BUFFER     u1550(.A(men_men_n1578_), .Y(men_men_n1579_));
  AOI220     u1551(.A0(men_men_n1579_), .A1(men_men_n1445_), .B0(men_men_n1118_), .B1(men_men_n1577_), .Y(men_men_n1580_));
  NA4        u1552(.A(men_men_n1580_), .B(men_men_n1576_), .C(men_men_n1573_), .D(men_men_n1572_), .Y(men_men_n1581_));
  NO4        u1553(.A(men_men_n1581_), .B(men_men_n1571_), .C(men_men_n1567_), .D(men_men_n1563_), .Y(men_men_n1582_));
  NA3        u1554(.A(men_men_n1582_), .B(men_men_n1560_), .C(men_men_n1553_), .Y(men_men_n1583_));
  NA3        u1555(.A(men_men_n1003_), .B(men_men_n143_), .C(men_men_n46_), .Y(men_men_n1584_));
  AOI210     u1556(.A0(men_men_n154_), .A1(c), .B0(men_men_n1584_), .Y(men_men_n1585_));
  INV        u1557(.A(men_men_n194_), .Y(men_men_n1586_));
  NA2        u1558(.A(men_men_n1586_), .B(men_men_n1519_), .Y(men_men_n1587_));
  AO210      u1559(.A0(men_men_n138_), .A1(l), .B0(men_men_n1472_), .Y(men_men_n1588_));
  NO2        u1560(.A(men_men_n72_), .B(c), .Y(men_men_n1589_));
  NO4        u1561(.A(men_men_n1432_), .B(men_men_n195_), .C(men_men_n470_), .D(men_men_n45_), .Y(men_men_n1590_));
  AOI210     u1562(.A0(men_men_n1529_), .A1(men_men_n1589_), .B0(men_men_n1590_), .Y(men_men_n1591_));
  NA3        u1563(.A(men_men_n1591_), .B(men_men_n1588_), .C(men_men_n1587_), .Y(men_men_n1592_));
  NO2        u1564(.A(men_men_n1592_), .B(men_men_n1585_), .Y(men_men_n1593_));
  NO4        u1565(.A(men_men_n236_), .B(men_men_n195_), .C(men_men_n271_), .D(k), .Y(men_men_n1594_));
  AOI210     u1566(.A0(men_men_n163_), .A1(men_men_n56_), .B0(men_men_n1554_), .Y(men_men_n1595_));
  NO2        u1567(.A(men_men_n1595_), .B(men_men_n1523_), .Y(men_men_n1596_));
  NO2        u1568(.A(men_men_n1584_), .B(men_men_n114_), .Y(men_men_n1597_));
  NOi21      u1569(.An(men_men_n1410_), .B(e), .Y(men_men_n1598_));
  NO4        u1570(.A(men_men_n1598_), .B(men_men_n1597_), .C(men_men_n1596_), .D(men_men_n1594_), .Y(men_men_n1599_));
  AOI220     u1571(.A0(men_men_n1578_), .A1(men_men_n669_), .B0(men_men_n1102_), .B1(men_men_n166_), .Y(men_men_n1600_));
  NOi31      u1572(.An(men_men_n30_), .B(men_men_n1600_), .C(n), .Y(men_men_n1601_));
  INV        u1573(.A(men_men_n1601_), .Y(men_men_n1602_));
  NA2        u1574(.A(men_men_n59_), .B(a), .Y(men_men_n1603_));
  NO2        u1575(.A(men_men_n1417_), .B(men_men_n122_), .Y(men_men_n1604_));
  OAI220     u1576(.A0(men_men_n1604_), .A1(men_men_n1472_), .B0(men_men_n1490_), .B1(men_men_n1603_), .Y(men_men_n1605_));
  NA4        u1577(.A(men_men_n1619_), .B(men_men_n1602_), .C(men_men_n1599_), .D(men_men_n1593_), .Y(men_men_n1606_));
  OR4        u1578(.A(men_men_n1606_), .B(men_men_n1583_), .C(men_men_n1539_), .D(men_men_n1494_), .Y(men04));
  NOi31      u1579(.An(men_men_n1480_), .B(men_men_n1481_), .C(men_men_n1090_), .Y(men_men_n1608_));
  NA2        u1580(.A(men_men_n1533_), .B(men_men_n867_), .Y(men_men_n1609_));
  NO4        u1581(.A(men_men_n1609_), .B(men_men_n1079_), .C(men_men_n505_), .D(j), .Y(men_men_n1610_));
  OR3        u1582(.A(men_men_n1610_), .B(men_men_n1608_), .C(men_men_n1108_), .Y(men_men_n1611_));
  NO3        u1583(.A(men_men_n1419_), .B(men_men_n93_), .C(k), .Y(men_men_n1612_));
  AOI210     u1584(.A0(men_men_n1612_), .A1(men_men_n1101_), .B0(men_men_n1237_), .Y(men_men_n1613_));
  NA2        u1585(.A(men_men_n1613_), .B(men_men_n1266_), .Y(men_men_n1614_));
  NO4        u1586(.A(men_men_n1614_), .B(men_men_n1611_), .C(men_men_n1116_), .D(men_men_n1095_), .Y(men_men_n1615_));
  NA4        u1587(.A(men_men_n1615_), .B(men_men_n1174_), .C(men_men_n1159_), .D(men_men_n1146_), .Y(men05));
  INV        u1588(.A(men_men_n1605_), .Y(men_men_n1619_));
  INV        u1589(.A(men_men_n631_), .Y(men_men_n1620_));
  INV        u1590(.A(men_men_n1498_), .Y(men_men_n1621_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule