library verilog;
use verilog.vl_types.all;
entity contador5_vlg_vec_tst is
end contador5_vlg_vec_tst;
