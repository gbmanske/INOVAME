//Benchmark atmr_misex3_1774_0.125

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1450_, men_men_n1451_, men_men_n1452_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  INV        o0001(.A(d), .Y(ori_ori_n30_));
  NA3        o0002(.A(e), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n31_));
  NOi32      o0003(.An(m), .Bn(l), .C(n), .Y(ori_ori_n32_));
  NOi32      o0004(.An(i), .Bn(g), .C(h), .Y(ori_ori_n33_));
  NA2        o0005(.A(ori_ori_n33_), .B(ori_ori_n32_), .Y(ori_ori_n34_));
  NOi32      o0006(.An(j), .Bn(g), .C(k), .Y(ori_ori_n35_));
  INV        o0007(.A(h), .Y(ori_ori_n36_));
  NAi21      o0008(.An(j), .B(l), .Y(ori_ori_n37_));
  NAi31      o0009(.An(n), .B(m), .C(l), .Y(ori_ori_n38_));
  INV        o0010(.A(i), .Y(ori_ori_n39_));
  AN2        o0011(.A(h), .B(g), .Y(ori_ori_n40_));
  INV        o0012(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o0013(.A(ori_ori_n41_), .B(ori_ori_n38_), .Y(ori_ori_n42_));
  NAi21      o0014(.An(n), .B(m), .Y(ori_ori_n43_));
  NOi32      o0015(.An(k), .Bn(h), .C(l), .Y(ori_ori_n44_));
  NOi32      o0016(.An(k), .Bn(h), .C(g), .Y(ori_ori_n45_));
  INV        o0017(.A(ori_ori_n45_), .Y(ori_ori_n46_));
  NO2        o0018(.A(ori_ori_n46_), .B(ori_ori_n43_), .Y(ori_ori_n47_));
  NO2        o0019(.A(ori_ori_n47_), .B(ori_ori_n42_), .Y(ori_ori_n48_));
  AOI210     o0020(.A0(ori_ori_n48_), .A1(ori_ori_n34_), .B0(ori_ori_n31_), .Y(ori_ori_n49_));
  INV        o0021(.A(c), .Y(ori_ori_n50_));
  NA2        o0022(.A(e), .B(b), .Y(ori_ori_n51_));
  INV        o0023(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  INV        o0024(.A(d), .Y(ori_ori_n53_));
  NAi21      o0025(.An(i), .B(h), .Y(ori_ori_n54_));
  NA2        o0026(.A(g), .B(f), .Y(ori_ori_n55_));
  NAi31      o0027(.An(l), .B(m), .C(k), .Y(ori_ori_n56_));
  NAi21      o0028(.An(e), .B(h), .Y(ori_ori_n57_));
  NAi41      o0029(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n58_));
  INV        o0030(.A(m), .Y(ori_ori_n59_));
  NOi21      o0031(.An(k), .B(l), .Y(ori_ori_n60_));
  NA2        o0032(.A(ori_ori_n60_), .B(ori_ori_n59_), .Y(ori_ori_n61_));
  AN4        o0033(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n62_));
  NOi21      o0034(.An(h), .B(f), .Y(ori_ori_n63_));
  NA2        o0035(.A(ori_ori_n63_), .B(ori_ori_n62_), .Y(ori_ori_n64_));
  NAi32      o0036(.An(m), .Bn(k), .C(j), .Y(ori_ori_n65_));
  NOi32      o0037(.An(h), .Bn(g), .C(f), .Y(ori_ori_n66_));
  OR2        o0038(.A(ori_ori_n64_), .B(ori_ori_n61_), .Y(ori_ori_n67_));
  INV        o0039(.A(ori_ori_n67_), .Y(ori_ori_n68_));
  INV        o0040(.A(n), .Y(ori_ori_n69_));
  NA2        o0041(.A(b), .B(ori_ori_n69_), .Y(ori_ori_n70_));
  INV        o0042(.A(j), .Y(ori_ori_n71_));
  AN3        o0043(.A(m), .B(k), .C(i), .Y(ori_ori_n72_));
  NA2        o0044(.A(ori_ori_n72_), .B(g), .Y(ori_ori_n73_));
  NO2        o0045(.A(ori_ori_n73_), .B(f), .Y(ori_ori_n74_));
  NAi32      o0046(.An(g), .Bn(f), .C(h), .Y(ori_ori_n75_));
  NAi31      o0047(.An(j), .B(m), .C(l), .Y(ori_ori_n76_));
  NO2        o0048(.A(ori_ori_n76_), .B(ori_ori_n75_), .Y(ori_ori_n77_));
  NA2        o0049(.A(m), .B(l), .Y(ori_ori_n78_));
  NAi31      o0050(.An(k), .B(j), .C(g), .Y(ori_ori_n79_));
  NO3        o0051(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(f), .Y(ori_ori_n80_));
  AN2        o0052(.A(j), .B(g), .Y(ori_ori_n81_));
  NA2        o0053(.A(m), .B(ori_ori_n81_), .Y(ori_ori_n82_));
  NO2        o0054(.A(ori_ori_n82_), .B(f), .Y(ori_ori_n83_));
  NAi41      o0055(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n84_));
  AN2        o0056(.A(e), .B(b), .Y(ori_ori_n85_));
  NOi21      o0057(.An(g), .B(f), .Y(ori_ori_n86_));
  NOi21      o0058(.An(i), .B(h), .Y(ori_ori_n87_));
  NA3        o0059(.A(ori_ori_n87_), .B(ori_ori_n86_), .C(m), .Y(ori_ori_n88_));
  INV        o0060(.A(a), .Y(ori_ori_n89_));
  NA2        o0061(.A(ori_ori_n85_), .B(ori_ori_n89_), .Y(ori_ori_n90_));
  INV        o0062(.A(l), .Y(ori_ori_n91_));
  NOi21      o0063(.An(m), .B(n), .Y(ori_ori_n92_));
  INV        o0064(.A(b), .Y(ori_ori_n93_));
  AN2        o0065(.A(k), .B(i), .Y(ori_ori_n94_));
  NOi32      o0066(.An(c), .Bn(a), .C(d), .Y(ori_ori_n95_));
  NA2        o0067(.A(ori_ori_n95_), .B(ori_ori_n92_), .Y(ori_ori_n96_));
  NO2        o0068(.A(ori_ori_n1031_), .B(ori_ori_n70_), .Y(ori_ori_n97_));
  NOi31      o0069(.An(k), .B(m), .C(j), .Y(ori_ori_n98_));
  NA3        o0070(.A(ori_ori_n98_), .B(ori_ori_n63_), .C(ori_ori_n62_), .Y(ori_ori_n99_));
  NOi31      o0071(.An(k), .B(m), .C(i), .Y(ori_ori_n100_));
  INV        o0072(.A(ori_ori_n99_), .Y(ori_ori_n101_));
  NOi32      o0073(.An(f), .Bn(b), .C(e), .Y(ori_ori_n102_));
  NAi21      o0074(.An(g), .B(h), .Y(ori_ori_n103_));
  NAi21      o0075(.An(m), .B(n), .Y(ori_ori_n104_));
  NAi31      o0076(.An(e), .B(f), .C(b), .Y(ori_ori_n105_));
  NAi31      o0077(.An(j), .B(k), .C(h), .Y(ori_ori_n106_));
  NO2        o0078(.A(k), .B(j), .Y(ori_ori_n107_));
  NO2        o0079(.A(ori_ori_n107_), .B(ori_ori_n104_), .Y(ori_ori_n108_));
  AN2        o0080(.A(k), .B(j), .Y(ori_ori_n109_));
  NAi21      o0081(.An(c), .B(b), .Y(ori_ori_n110_));
  NA2        o0082(.A(f), .B(d), .Y(ori_ori_n111_));
  NO3        o0083(.A(ori_ori_n111_), .B(ori_ori_n110_), .C(ori_ori_n103_), .Y(ori_ori_n112_));
  NA2        o0084(.A(h), .B(c), .Y(ori_ori_n113_));
  NAi31      o0085(.An(f), .B(e), .C(b), .Y(ori_ori_n114_));
  NA2        o0086(.A(ori_ori_n112_), .B(ori_ori_n108_), .Y(ori_ori_n115_));
  NA2        o0087(.A(d), .B(b), .Y(ori_ori_n116_));
  NAi21      o0088(.An(e), .B(f), .Y(ori_ori_n117_));
  NO2        o0089(.A(ori_ori_n117_), .B(ori_ori_n116_), .Y(ori_ori_n118_));
  NA2        o0090(.A(b), .B(a), .Y(ori_ori_n119_));
  NAi21      o0091(.An(c), .B(d), .Y(ori_ori_n120_));
  NAi31      o0092(.An(l), .B(k), .C(h), .Y(ori_ori_n121_));
  NO2        o0093(.A(ori_ori_n104_), .B(ori_ori_n121_), .Y(ori_ori_n122_));
  NA2        o0094(.A(ori_ori_n122_), .B(ori_ori_n118_), .Y(ori_ori_n123_));
  NAi31      o0095(.An(ori_ori_n101_), .B(ori_ori_n123_), .C(ori_ori_n115_), .Y(ori_ori_n124_));
  NAi31      o0096(.An(e), .B(f), .C(b), .Y(ori_ori_n125_));
  INV        o0097(.A(ori_ori_n125_), .Y(ori_ori_n126_));
  NOi21      o0098(.An(h), .B(i), .Y(ori_ori_n127_));
  NOi21      o0099(.An(k), .B(m), .Y(ori_ori_n128_));
  NA3        o0100(.A(ori_ori_n128_), .B(ori_ori_n127_), .C(n), .Y(ori_ori_n129_));
  NOi21      o0101(.An(ori_ori_n126_), .B(ori_ori_n129_), .Y(ori_ori_n130_));
  NOi21      o0102(.An(h), .B(g), .Y(ori_ori_n131_));
  NAi31      o0103(.An(d), .B(f), .C(c), .Y(ori_ori_n132_));
  NAi31      o0104(.An(e), .B(f), .C(c), .Y(ori_ori_n133_));
  NA2        o0105(.A(ori_ori_n133_), .B(ori_ori_n132_), .Y(ori_ori_n134_));
  NA2        o0106(.A(j), .B(h), .Y(ori_ori_n135_));
  OR3        o0107(.A(n), .B(m), .C(k), .Y(ori_ori_n136_));
  NO2        o0108(.A(ori_ori_n136_), .B(ori_ori_n135_), .Y(ori_ori_n137_));
  NAi32      o0109(.An(m), .Bn(k), .C(n), .Y(ori_ori_n138_));
  NO2        o0110(.A(ori_ori_n138_), .B(ori_ori_n135_), .Y(ori_ori_n139_));
  AOI220     o0111(.A0(ori_ori_n139_), .A1(ori_ori_n126_), .B0(ori_ori_n137_), .B1(ori_ori_n134_), .Y(ori_ori_n140_));
  NO2        o0112(.A(n), .B(m), .Y(ori_ori_n141_));
  NA2        o0113(.A(ori_ori_n141_), .B(ori_ori_n44_), .Y(ori_ori_n142_));
  NAi21      o0114(.An(f), .B(e), .Y(ori_ori_n143_));
  NA2        o0115(.A(d), .B(c), .Y(ori_ori_n144_));
  NO2        o0116(.A(ori_ori_n144_), .B(ori_ori_n143_), .Y(ori_ori_n145_));
  NOi21      o0117(.An(ori_ori_n145_), .B(ori_ori_n142_), .Y(ori_ori_n146_));
  NAi31      o0118(.An(m), .B(n), .C(b), .Y(ori_ori_n147_));
  NA2        o0119(.A(k), .B(i), .Y(ori_ori_n148_));
  NAi21      o0120(.An(h), .B(f), .Y(ori_ori_n149_));
  NO2        o0121(.A(ori_ori_n149_), .B(ori_ori_n148_), .Y(ori_ori_n150_));
  NO2        o0122(.A(ori_ori_n147_), .B(ori_ori_n120_), .Y(ori_ori_n151_));
  NA2        o0123(.A(ori_ori_n151_), .B(ori_ori_n150_), .Y(ori_ori_n152_));
  NOi32      o0124(.An(f), .Bn(c), .C(d), .Y(ori_ori_n153_));
  NOi32      o0125(.An(f), .Bn(c), .C(e), .Y(ori_ori_n154_));
  NO2        o0126(.A(ori_ori_n154_), .B(ori_ori_n153_), .Y(ori_ori_n155_));
  OR2        o0127(.A(ori_ori_n142_), .B(ori_ori_n155_), .Y(ori_ori_n156_));
  NAi41      o0128(.An(ori_ori_n146_), .B(ori_ori_n156_), .C(ori_ori_n152_), .D(ori_ori_n140_), .Y(ori_ori_n157_));
  OR3        o0129(.A(ori_ori_n157_), .B(ori_ori_n130_), .C(ori_ori_n124_), .Y(ori_ori_n158_));
  NO4        o0130(.A(ori_ori_n158_), .B(ori_ori_n97_), .C(ori_ori_n68_), .D(ori_ori_n49_), .Y(ori_ori_n159_));
  NAi31      o0131(.An(n), .B(h), .C(g), .Y(ori_ori_n160_));
  NO2        o0132(.A(ori_ori_n160_), .B(ori_ori_n1032_), .Y(ori_ori_n161_));
  NOi32      o0133(.An(m), .Bn(k), .C(l), .Y(ori_ori_n162_));
  NA2        o0134(.A(ori_ori_n162_), .B(g), .Y(ori_ori_n163_));
  NO2        o0135(.A(ori_ori_n163_), .B(n), .Y(ori_ori_n164_));
  NA4        o0136(.A(k), .B(ori_ori_n92_), .C(i), .D(g), .Y(ori_ori_n165_));
  NO2        o0137(.A(ori_ori_n164_), .B(ori_ori_n161_), .Y(ori_ori_n166_));
  NAi41      o0138(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n167_));
  INV        o0139(.A(ori_ori_n167_), .Y(ori_ori_n168_));
  INV        o0140(.A(f), .Y(ori_ori_n169_));
  INV        o0141(.A(g), .Y(ori_ori_n170_));
  NOi31      o0142(.An(i), .B(j), .C(h), .Y(ori_ori_n171_));
  NOi21      o0143(.An(l), .B(m), .Y(ori_ori_n172_));
  NA2        o0144(.A(ori_ori_n172_), .B(ori_ori_n171_), .Y(ori_ori_n173_));
  NO3        o0145(.A(ori_ori_n173_), .B(ori_ori_n170_), .C(ori_ori_n169_), .Y(ori_ori_n174_));
  NA2        o0146(.A(ori_ori_n174_), .B(ori_ori_n168_), .Y(ori_ori_n175_));
  OAI210     o0147(.A0(ori_ori_n166_), .A1(ori_ori_n31_), .B0(ori_ori_n175_), .Y(ori_ori_n176_));
  NOi21      o0148(.An(n), .B(m), .Y(ori_ori_n177_));
  OR2        o0149(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n178_));
  NAi21      o0150(.An(j), .B(h), .Y(ori_ori_n179_));
  XN2        o0151(.A(i), .B(h), .Y(ori_ori_n180_));
  NOi31      o0152(.An(k), .B(n), .C(m), .Y(ori_ori_n181_));
  NAi31      o0153(.An(f), .B(e), .C(c), .Y(ori_ori_n182_));
  NA3        o0154(.A(e), .B(c), .C(b), .Y(ori_ori_n183_));
  NAi32      o0155(.An(m), .Bn(i), .C(k), .Y(ori_ori_n184_));
  INV        o0156(.A(k), .Y(ori_ori_n185_));
  NAi21      o0157(.An(n), .B(a), .Y(ori_ori_n186_));
  NO2        o0158(.A(ori_ori_n186_), .B(ori_ori_n116_), .Y(ori_ori_n187_));
  NAi41      o0159(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n188_));
  NO2        o0160(.A(ori_ori_n188_), .B(e), .Y(ori_ori_n189_));
  NO2        o0161(.A(g), .B(ori_ori_n84_), .Y(ori_ori_n190_));
  NA2        o0162(.A(ori_ori_n190_), .B(ori_ori_n102_), .Y(ori_ori_n191_));
  NAi41      o0163(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n192_));
  NO2        o0164(.A(ori_ori_n192_), .B(ori_ori_n169_), .Y(ori_ori_n193_));
  NA2        o0165(.A(ori_ori_n128_), .B(ori_ori_n87_), .Y(ori_ori_n194_));
  NAi21      o0166(.An(ori_ori_n194_), .B(ori_ori_n193_), .Y(ori_ori_n195_));
  NO2        o0167(.A(n), .B(a), .Y(ori_ori_n196_));
  NAi21      o0168(.An(h), .B(i), .Y(ori_ori_n197_));
  NA2        o0169(.A(ori_ori_n141_), .B(k), .Y(ori_ori_n198_));
  NO2        o0170(.A(ori_ori_n198_), .B(ori_ori_n197_), .Y(ori_ori_n199_));
  NA2        o0171(.A(ori_ori_n199_), .B(ori_ori_n153_), .Y(ori_ori_n200_));
  NA3        o0172(.A(ori_ori_n200_), .B(ori_ori_n195_), .C(ori_ori_n191_), .Y(ori_ori_n201_));
  NOi21      o0173(.An(g), .B(e), .Y(ori_ori_n202_));
  NO2        o0174(.A(ori_ori_n58_), .B(ori_ori_n59_), .Y(ori_ori_n203_));
  NAi21      o0175(.An(f), .B(g), .Y(ori_ori_n204_));
  NOi31      o0176(.An(ori_ori_n178_), .B(ori_ori_n201_), .C(ori_ori_n176_), .Y(ori_ori_n205_));
  NA3        o0177(.A(ori_ori_n53_), .B(c), .C(b), .Y(ori_ori_n206_));
  NAi21      o0178(.An(h), .B(g), .Y(ori_ori_n207_));
  NO2        o0179(.A(ori_ori_n194_), .B(ori_ori_n204_), .Y(ori_ori_n208_));
  NA3        o0180(.A(ori_ori_n128_), .B(ori_ori_n127_), .C(ori_ori_n69_), .Y(ori_ori_n209_));
  NO2        o0181(.A(ori_ori_n209_), .B(ori_ori_n155_), .Y(ori_ori_n210_));
  INV        o0182(.A(ori_ori_n210_), .Y(ori_ori_n211_));
  NA3        o0183(.A(e), .B(c), .C(b), .Y(ori_ori_n212_));
  NOi21      o0184(.An(l), .B(j), .Y(ori_ori_n213_));
  NA2        o0185(.A(ori_ori_n131_), .B(ori_ori_n213_), .Y(ori_ori_n214_));
  OR3        o0186(.A(ori_ori_n58_), .B(ori_ori_n59_), .C(e), .Y(ori_ori_n215_));
  AOI210     o0187(.A0(ori_ori_n1033_), .A1(ori_ori_n214_), .B0(ori_ori_n215_), .Y(ori_ori_n216_));
  INV        o0188(.A(ori_ori_n216_), .Y(ori_ori_n217_));
  NAi32      o0189(.An(j), .Bn(h), .C(i), .Y(ori_ori_n218_));
  NAi21      o0190(.An(m), .B(l), .Y(ori_ori_n219_));
  NA2        o0191(.A(h), .B(g), .Y(ori_ori_n220_));
  NA2        o0192(.A(ori_ori_n217_), .B(ori_ori_n211_), .Y(ori_ori_n221_));
  NO2        o0193(.A(ori_ori_n114_), .B(d), .Y(ori_ori_n222_));
  NAi32      o0194(.An(n), .Bn(m), .C(l), .Y(ori_ori_n223_));
  NO2        o0195(.A(ori_ori_n223_), .B(ori_ori_n218_), .Y(ori_ori_n224_));
  NA2        o0196(.A(ori_ori_n224_), .B(ori_ori_n145_), .Y(ori_ori_n225_));
  NO2        o0197(.A(ori_ori_n1030_), .B(ori_ori_n221_), .Y(ori_ori_n226_));
  NAi21      o0198(.An(m), .B(k), .Y(ori_ori_n227_));
  NO2        o0199(.A(ori_ori_n180_), .B(ori_ori_n227_), .Y(ori_ori_n228_));
  NAi41      o0200(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n229_));
  NA2        o0201(.A(e), .B(c), .Y(ori_ori_n230_));
  NO3        o0202(.A(ori_ori_n230_), .B(n), .C(d), .Y(ori_ori_n231_));
  NAi31      o0203(.An(d), .B(e), .C(b), .Y(ori_ori_n232_));
  NO4        o0204(.A(ori_ori_n229_), .B(ori_ori_n65_), .C(ori_ori_n57_), .D(ori_ori_n170_), .Y(ori_ori_n233_));
  NA2        o0205(.A(ori_ori_n196_), .B(ori_ori_n85_), .Y(ori_ori_n234_));
  OR2        o0206(.A(ori_ori_n234_), .B(ori_ori_n163_), .Y(ori_ori_n235_));
  NOi31      o0207(.An(l), .B(n), .C(m), .Y(ori_ori_n236_));
  NA2        o0208(.A(ori_ori_n236_), .B(ori_ori_n171_), .Y(ori_ori_n237_));
  NO2        o0209(.A(ori_ori_n237_), .B(ori_ori_n155_), .Y(ori_ori_n238_));
  NAi32      o0210(.An(ori_ori_n238_), .Bn(ori_ori_n233_), .C(ori_ori_n235_), .Y(ori_ori_n239_));
  NAi32      o0211(.An(m), .Bn(j), .C(k), .Y(ori_ori_n240_));
  NAi41      o0212(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n241_));
  NA2        o0213(.A(ori_ori_n167_), .B(ori_ori_n241_), .Y(ori_ori_n242_));
  NOi31      o0214(.An(j), .B(m), .C(k), .Y(ori_ori_n243_));
  NO2        o0215(.A(ori_ori_n98_), .B(ori_ori_n243_), .Y(ori_ori_n244_));
  AN3        o0216(.A(h), .B(g), .C(f), .Y(ori_ori_n245_));
  NAi31      o0217(.An(ori_ori_n244_), .B(ori_ori_n245_), .C(ori_ori_n242_), .Y(ori_ori_n246_));
  NO2        o0218(.A(ori_ori_n219_), .B(ori_ori_n218_), .Y(ori_ori_n247_));
  NO2        o0219(.A(ori_ori_n173_), .B(g), .Y(ori_ori_n248_));
  NO2        o0220(.A(ori_ori_n125_), .B(ori_ori_n69_), .Y(ori_ori_n249_));
  AOI220     o0221(.A0(ori_ori_n249_), .A1(ori_ori_n248_), .B0(ori_ori_n193_), .B1(ori_ori_n247_), .Y(ori_ori_n250_));
  NA2        o0222(.A(ori_ori_n250_), .B(ori_ori_n246_), .Y(ori_ori_n251_));
  NA3        o0223(.A(h), .B(g), .C(f), .Y(ori_ori_n252_));
  NO2        o0224(.A(ori_ori_n252_), .B(ori_ori_n61_), .Y(ori_ori_n253_));
  NA2        o0225(.A(ori_ori_n241_), .B(ori_ori_n167_), .Y(ori_ori_n254_));
  NA2        o0226(.A(ori_ori_n131_), .B(e), .Y(ori_ori_n255_));
  NA2        o0227(.A(ori_ori_n254_), .B(ori_ori_n253_), .Y(ori_ori_n256_));
  NOi32      o0228(.An(j), .Bn(g), .C(i), .Y(ori_ori_n257_));
  NA2        o0229(.A(ori_ori_n257_), .B(ori_ori_n92_), .Y(ori_ori_n258_));
  AO210      o0230(.A0(ori_ori_n90_), .A1(ori_ori_n31_), .B0(ori_ori_n258_), .Y(ori_ori_n259_));
  INV        o0231(.A(ori_ori_n227_), .Y(ori_ori_n260_));
  NO3        o0232(.A(ori_ori_n229_), .B(ori_ori_n57_), .C(ori_ori_n170_), .Y(ori_ori_n261_));
  NA2        o0233(.A(ori_ori_n261_), .B(ori_ori_n260_), .Y(ori_ori_n262_));
  NA2        o0234(.A(g), .B(k), .Y(ori_ori_n263_));
  NA3        o0235(.A(m), .B(ori_ori_n91_), .C(ori_ori_n169_), .Y(ori_ori_n264_));
  NA3        o0236(.A(ori_ori_n162_), .B(g), .C(ori_ori_n169_), .Y(ori_ori_n265_));
  NAi41      o0237(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n266_));
  NA2        o0238(.A(ori_ori_n45_), .B(ori_ori_n92_), .Y(ori_ori_n267_));
  NO2        o0239(.A(ori_ori_n267_), .B(ori_ori_n266_), .Y(ori_ori_n268_));
  NA3        o0240(.A(ori_ori_n262_), .B(ori_ori_n259_), .C(ori_ori_n256_), .Y(ori_ori_n269_));
  NO3        o0241(.A(ori_ori_n269_), .B(ori_ori_n251_), .C(ori_ori_n239_), .Y(ori_ori_n270_));
  NA4        o0242(.A(ori_ori_n270_), .B(ori_ori_n226_), .C(ori_ori_n205_), .D(ori_ori_n159_), .Y(ori10));
  NA3        o0243(.A(m), .B(k), .C(i), .Y(ori_ori_n272_));
  NOi21      o0244(.An(e), .B(f), .Y(ori_ori_n273_));
  NO3        o0245(.A(ori_ori_n120_), .B(n), .C(ori_ori_n89_), .Y(ori_ori_n274_));
  NAi31      o0246(.An(b), .B(f), .C(c), .Y(ori_ori_n275_));
  INV        o0247(.A(ori_ori_n275_), .Y(ori_ori_n276_));
  NOi32      o0248(.An(k), .Bn(h), .C(j), .Y(ori_ori_n277_));
  NA2        o0249(.A(ori_ori_n277_), .B(ori_ori_n177_), .Y(ori_ori_n278_));
  NA2        o0250(.A(ori_ori_n129_), .B(ori_ori_n278_), .Y(ori_ori_n279_));
  NA2        o0251(.A(ori_ori_n279_), .B(ori_ori_n276_), .Y(ori_ori_n280_));
  AN2        o0252(.A(j), .B(h), .Y(ori_ori_n281_));
  NO3        o0253(.A(n), .B(m), .C(k), .Y(ori_ori_n282_));
  NA2        o0254(.A(ori_ori_n282_), .B(ori_ori_n281_), .Y(ori_ori_n283_));
  NO3        o0255(.A(ori_ori_n283_), .B(ori_ori_n120_), .C(ori_ori_n169_), .Y(ori_ori_n284_));
  OR2        o0256(.A(m), .B(k), .Y(ori_ori_n285_));
  NO2        o0257(.A(ori_ori_n135_), .B(ori_ori_n285_), .Y(ori_ori_n286_));
  NA4        o0258(.A(n), .B(f), .C(c), .D(ori_ori_n93_), .Y(ori_ori_n287_));
  NOi21      o0259(.An(ori_ori_n286_), .B(ori_ori_n287_), .Y(ori_ori_n288_));
  NOi32      o0260(.An(d), .Bn(a), .C(c), .Y(ori_ori_n289_));
  NA2        o0261(.A(ori_ori_n289_), .B(ori_ori_n143_), .Y(ori_ori_n290_));
  NAi21      o0262(.An(i), .B(g), .Y(ori_ori_n291_));
  NAi31      o0263(.An(k), .B(m), .C(j), .Y(ori_ori_n292_));
  NO3        o0264(.A(ori_ori_n292_), .B(ori_ori_n291_), .C(n), .Y(ori_ori_n293_));
  NOi21      o0265(.An(ori_ori_n293_), .B(ori_ori_n290_), .Y(ori_ori_n294_));
  NO3        o0266(.A(ori_ori_n294_), .B(ori_ori_n288_), .C(ori_ori_n284_), .Y(ori_ori_n295_));
  NO2        o0267(.A(ori_ori_n287_), .B(ori_ori_n219_), .Y(ori_ori_n296_));
  NOi32      o0268(.An(f), .Bn(d), .C(c), .Y(ori_ori_n297_));
  NA2        o0269(.A(ori_ori_n295_), .B(ori_ori_n280_), .Y(ori_ori_n298_));
  NO2        o0270(.A(ori_ori_n53_), .B(ori_ori_n93_), .Y(ori_ori_n299_));
  NA2        o0271(.A(ori_ori_n196_), .B(ori_ori_n299_), .Y(ori_ori_n300_));
  INV        o0272(.A(e), .Y(ori_ori_n301_));
  NA2        o0273(.A(ori_ori_n40_), .B(e), .Y(ori_ori_n302_));
  OAI220     o0274(.A0(ori_ori_n302_), .A1(ori_ori_n1032_), .B0(ori_ori_n163_), .B1(ori_ori_n301_), .Y(ori_ori_n303_));
  NO2        o0275(.A(ori_ori_n73_), .B(ori_ori_n301_), .Y(ori_ori_n304_));
  NO2        o0276(.A(ori_ori_n82_), .B(ori_ori_n301_), .Y(ori_ori_n305_));
  NO3        o0277(.A(ori_ori_n305_), .B(ori_ori_n304_), .C(ori_ori_n303_), .Y(ori_ori_n306_));
  NOi32      o0278(.An(h), .Bn(e), .C(g), .Y(ori_ori_n307_));
  AN3        o0279(.A(m), .B(l), .C(i), .Y(ori_ori_n308_));
  AN3        o0280(.A(h), .B(g), .C(e), .Y(ori_ori_n309_));
  NO2        o0281(.A(ori_ori_n306_), .B(ori_ori_n300_), .Y(ori_ori_n310_));
  NA3        o0282(.A(ori_ori_n289_), .B(ori_ori_n143_), .C(ori_ori_n69_), .Y(ori_ori_n311_));
  NAi31      o0283(.An(b), .B(c), .C(a), .Y(ori_ori_n312_));
  NO2        o0284(.A(ori_ori_n312_), .B(n), .Y(ori_ori_n313_));
  NA2        o0285(.A(ori_ori_n45_), .B(m), .Y(ori_ori_n314_));
  NO2        o0286(.A(ori_ori_n310_), .B(ori_ori_n298_), .Y(ori_ori_n315_));
  NA2        o0287(.A(i), .B(g), .Y(ori_ori_n316_));
  NOi21      o0288(.An(a), .B(n), .Y(ori_ori_n317_));
  NOi21      o0289(.An(d), .B(c), .Y(ori_ori_n318_));
  NA2        o0290(.A(ori_ori_n318_), .B(ori_ori_n317_), .Y(ori_ori_n319_));
  NA3        o0291(.A(i), .B(g), .C(f), .Y(ori_ori_n320_));
  OR2        o0292(.A(ori_ori_n320_), .B(ori_ori_n56_), .Y(ori_ori_n321_));
  NA3        o0293(.A(ori_ori_n308_), .B(g), .C(ori_ori_n143_), .Y(ori_ori_n322_));
  AOI210     o0294(.A0(ori_ori_n322_), .A1(ori_ori_n321_), .B0(ori_ori_n319_), .Y(ori_ori_n323_));
  INV        o0295(.A(ori_ori_n323_), .Y(ori_ori_n324_));
  OR2        o0296(.A(n), .B(m), .Y(ori_ori_n325_));
  NO2        o0297(.A(ori_ori_n325_), .B(ori_ori_n121_), .Y(ori_ori_n326_));
  NO2        o0298(.A(ori_ori_n144_), .B(ori_ori_n117_), .Y(ori_ori_n327_));
  OAI210     o0299(.A0(ori_ori_n326_), .A1(ori_ori_n137_), .B0(ori_ori_n327_), .Y(ori_ori_n328_));
  INV        o0300(.A(ori_ori_n267_), .Y(ori_ori_n329_));
  NO2        o0301(.A(ori_ori_n312_), .B(ori_ori_n43_), .Y(ori_ori_n330_));
  NO2        o0302(.A(ori_ori_n55_), .B(ori_ori_n91_), .Y(ori_ori_n331_));
  NAi21      o0303(.An(k), .B(j), .Y(ori_ori_n332_));
  NA2        o0304(.A(ori_ori_n197_), .B(ori_ori_n332_), .Y(ori_ori_n333_));
  NA3        o0305(.A(ori_ori_n333_), .B(ori_ori_n331_), .C(ori_ori_n330_), .Y(ori_ori_n334_));
  NAi21      o0306(.An(e), .B(d), .Y(ori_ori_n335_));
  INV        o0307(.A(ori_ori_n335_), .Y(ori_ori_n336_));
  NO2        o0308(.A(ori_ori_n198_), .B(ori_ori_n169_), .Y(ori_ori_n337_));
  NA2        o0309(.A(ori_ori_n334_), .B(ori_ori_n328_), .Y(ori_ori_n338_));
  NO2        o0310(.A(ori_ori_n237_), .B(ori_ori_n169_), .Y(ori_ori_n339_));
  NA2        o0311(.A(ori_ori_n339_), .B(ori_ori_n336_), .Y(ori_ori_n340_));
  NOi31      o0312(.An(n), .B(m), .C(k), .Y(ori_ori_n341_));
  AOI220     o0313(.A0(ori_ori_n341_), .A1(ori_ori_n281_), .B0(ori_ori_n177_), .B1(ori_ori_n44_), .Y(ori_ori_n342_));
  NAi31      o0314(.An(g), .B(f), .C(c), .Y(ori_ori_n343_));
  NA2        o0315(.A(ori_ori_n340_), .B(ori_ori_n225_), .Y(ori_ori_n344_));
  NOi31      o0316(.An(ori_ori_n324_), .B(ori_ori_n344_), .C(ori_ori_n338_), .Y(ori_ori_n345_));
  NOi32      o0317(.An(c), .Bn(a), .C(b), .Y(ori_ori_n346_));
  NA2        o0318(.A(ori_ori_n346_), .B(ori_ori_n92_), .Y(ori_ori_n347_));
  AN2        o0319(.A(e), .B(d), .Y(ori_ori_n348_));
  NO2        o0320(.A(ori_ori_n103_), .B(ori_ori_n37_), .Y(ori_ori_n349_));
  NA2        o0321(.A(ori_ori_n349_), .B(f), .Y(ori_ori_n350_));
  NO2        o0322(.A(ori_ori_n350_), .B(ori_ori_n347_), .Y(ori_ori_n351_));
  NOi21      o0323(.An(a), .B(b), .Y(ori_ori_n352_));
  NA3        o0324(.A(e), .B(d), .C(c), .Y(ori_ori_n353_));
  NAi21      o0325(.An(ori_ori_n353_), .B(ori_ori_n352_), .Y(ori_ori_n354_));
  NO2        o0326(.A(ori_ori_n311_), .B(ori_ori_n163_), .Y(ori_ori_n355_));
  NA2        o0327(.A(ori_ori_n276_), .B(ori_ori_n122_), .Y(ori_ori_n356_));
  OR2        o0328(.A(k), .B(j), .Y(ori_ori_n357_));
  NA2        o0329(.A(l), .B(k), .Y(ori_ori_n358_));
  NA2        o0330(.A(ori_ori_n357_), .B(ori_ori_n177_), .Y(ori_ori_n359_));
  AOI210     o0331(.A0(ori_ori_n184_), .A1(ori_ori_n240_), .B0(ori_ori_n69_), .Y(ori_ori_n360_));
  BUFFER     o0332(.A(ori_ori_n359_), .Y(ori_ori_n361_));
  OR3        o0333(.A(ori_ori_n361_), .B(ori_ori_n113_), .C(ori_ori_n105_), .Y(ori_ori_n362_));
  INV        o0334(.A(ori_ori_n99_), .Y(ori_ori_n363_));
  NO3        o0335(.A(ori_ori_n311_), .B(ori_ori_n76_), .C(ori_ori_n103_), .Y(ori_ori_n364_));
  NO2        o0336(.A(ori_ori_n364_), .B(ori_ori_n363_), .Y(ori_ori_n365_));
  NA3        o0337(.A(ori_ori_n365_), .B(ori_ori_n362_), .C(ori_ori_n356_), .Y(ori_ori_n366_));
  NO3        o0338(.A(ori_ori_n366_), .B(ori_ori_n355_), .C(ori_ori_n351_), .Y(ori_ori_n367_));
  NO2        o0339(.A(ori_ori_n149_), .B(ori_ori_n50_), .Y(ori_ori_n368_));
  NAi31      o0340(.An(j), .B(l), .C(i), .Y(ori_ori_n369_));
  OAI210     o0341(.A0(ori_ori_n369_), .A1(ori_ori_n104_), .B0(ori_ori_n84_), .Y(ori_ori_n370_));
  NA2        o0342(.A(ori_ori_n370_), .B(ori_ori_n368_), .Y(ori_ori_n371_));
  NO2        o0343(.A(ori_ori_n290_), .B(ori_ori_n267_), .Y(ori_ori_n372_));
  NO2        o0344(.A(ori_ori_n372_), .B(ori_ori_n146_), .Y(ori_ori_n373_));
  NA3        o0345(.A(ori_ori_n373_), .B(ori_ori_n371_), .C(ori_ori_n178_), .Y(ori_ori_n374_));
  OAI210     o0346(.A0(ori_ori_n100_), .A1(ori_ori_n98_), .B0(n), .Y(ori_ori_n375_));
  NO2        o0347(.A(ori_ori_n375_), .B(ori_ori_n103_), .Y(ori_ori_n376_));
  XO2        o0348(.A(i), .B(h), .Y(ori_ori_n377_));
  NA2        o0349(.A(ori_ori_n342_), .B(ori_ori_n278_), .Y(ori_ori_n378_));
  NAi31      o0350(.An(c), .B(f), .C(d), .Y(ori_ori_n379_));
  NO2        o0351(.A(ori_ori_n209_), .B(ori_ori_n379_), .Y(ori_ori_n380_));
  BUFFER     o0352(.A(ori_ori_n67_), .Y(ori_ori_n381_));
  NA2        o0353(.A(ori_ori_n181_), .B(ori_ori_n87_), .Y(ori_ori_n382_));
  AOI210     o0354(.A0(ori_ori_n382_), .A1(ori_ori_n142_), .B0(ori_ori_n379_), .Y(ori_ori_n383_));
  AOI210     o0355(.A0(ori_ori_n258_), .A1(ori_ori_n34_), .B0(ori_ori_n354_), .Y(ori_ori_n384_));
  NO2        o0356(.A(ori_ori_n384_), .B(ori_ori_n383_), .Y(ori_ori_n385_));
  NA3        o0357(.A(ori_ori_n35_), .B(m), .C(f), .Y(ori_ori_n386_));
  INV        o0358(.A(ori_ori_n216_), .Y(ori_ori_n387_));
  NA3        o0359(.A(ori_ori_n387_), .B(ori_ori_n385_), .C(ori_ori_n381_), .Y(ori_ori_n388_));
  NO2        o0360(.A(ori_ori_n388_), .B(ori_ori_n374_), .Y(ori_ori_n389_));
  NA4        o0361(.A(ori_ori_n389_), .B(ori_ori_n367_), .C(ori_ori_n345_), .D(ori_ori_n315_), .Y(ori11));
  NO2        o0362(.A(ori_ori_n58_), .B(f), .Y(ori_ori_n391_));
  NA2        o0363(.A(j), .B(g), .Y(ori_ori_n392_));
  NAi31      o0364(.An(i), .B(m), .C(l), .Y(ori_ori_n393_));
  NA3        o0365(.A(m), .B(k), .C(j), .Y(ori_ori_n394_));
  OAI220     o0366(.A0(ori_ori_n394_), .A1(ori_ori_n103_), .B0(ori_ori_n393_), .B1(ori_ori_n392_), .Y(ori_ori_n395_));
  NA2        o0367(.A(ori_ori_n395_), .B(ori_ori_n391_), .Y(ori_ori_n396_));
  NOi32      o0368(.An(e), .Bn(b), .C(f), .Y(ori_ori_n397_));
  NA2        o0369(.A(ori_ori_n40_), .B(j), .Y(ori_ori_n398_));
  NAi31      o0370(.An(d), .B(e), .C(a), .Y(ori_ori_n399_));
  NO2        o0371(.A(ori_ori_n399_), .B(n), .Y(ori_ori_n400_));
  NA2        o0372(.A(ori_ori_n400_), .B(ori_ori_n83_), .Y(ori_ori_n401_));
  NAi31      o0373(.An(f), .B(e), .C(a), .Y(ori_ori_n402_));
  AN2        o0374(.A(ori_ori_n402_), .B(ori_ori_n266_), .Y(ori_ori_n403_));
  AOI210     o0375(.A0(ori_ori_n403_), .A1(ori_ori_n290_), .B0(ori_ori_n207_), .Y(ori_ori_n404_));
  NA2        o0376(.A(j), .B(i), .Y(ori_ori_n405_));
  NAi31      o0377(.An(n), .B(m), .C(k), .Y(ori_ori_n406_));
  NO3        o0378(.A(ori_ori_n406_), .B(ori_ori_n405_), .C(ori_ori_n91_), .Y(ori_ori_n407_));
  NO4        o0379(.A(n), .B(d), .C(ori_ori_n93_), .D(a), .Y(ori_ori_n408_));
  OR2        o0380(.A(n), .B(c), .Y(ori_ori_n409_));
  NO2        o0381(.A(ori_ori_n409_), .B(ori_ori_n119_), .Y(ori_ori_n410_));
  NO2        o0382(.A(ori_ori_n410_), .B(ori_ori_n408_), .Y(ori_ori_n411_));
  NA2        o0383(.A(ori_ori_n395_), .B(f), .Y(ori_ori_n412_));
  NO2        o0384(.A(ori_ori_n412_), .B(ori_ori_n411_), .Y(ori_ori_n413_));
  AOI210     o0385(.A0(ori_ori_n407_), .A1(ori_ori_n404_), .B0(ori_ori_n413_), .Y(ori_ori_n414_));
  NA2        o0386(.A(ori_ori_n109_), .B(ori_ori_n33_), .Y(ori_ori_n415_));
  OAI220     o0387(.A0(ori_ori_n415_), .A1(m), .B0(ori_ori_n398_), .B1(ori_ori_n184_), .Y(ori_ori_n416_));
  NOi41      o0388(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n417_));
  NAi32      o0389(.An(e), .Bn(b), .C(c), .Y(ori_ori_n418_));
  OR2        o0390(.A(ori_ori_n418_), .B(ori_ori_n69_), .Y(ori_ori_n419_));
  AN2        o0391(.A(ori_ori_n241_), .B(ori_ori_n229_), .Y(ori_ori_n420_));
  NA2        o0392(.A(ori_ori_n420_), .B(ori_ori_n419_), .Y(ori_ori_n421_));
  OA210      o0393(.A0(ori_ori_n421_), .A1(ori_ori_n417_), .B0(ori_ori_n416_), .Y(ori_ori_n422_));
  OAI220     o0394(.A0(ori_ori_n292_), .A1(ori_ori_n291_), .B0(ori_ori_n393_), .B1(ori_ori_n392_), .Y(ori_ori_n423_));
  NAi31      o0395(.An(d), .B(c), .C(a), .Y(ori_ori_n424_));
  NO2        o0396(.A(ori_ori_n424_), .B(n), .Y(ori_ori_n425_));
  NO2        o0397(.A(ori_ori_n182_), .B(ori_ori_n89_), .Y(ori_ori_n426_));
  NA2        o0398(.A(ori_ori_n293_), .B(ori_ori_n426_), .Y(ori_ori_n427_));
  INV        o0399(.A(ori_ori_n427_), .Y(ori_ori_n428_));
  NAi32      o0400(.An(d), .Bn(a), .C(b), .Y(ori_ori_n429_));
  NO2        o0401(.A(ori_ori_n429_), .B(ori_ori_n43_), .Y(ori_ori_n430_));
  NA2        o0402(.A(h), .B(f), .Y(ori_ori_n431_));
  NO2        o0403(.A(ori_ori_n431_), .B(ori_ori_n79_), .Y(ori_ori_n432_));
  NO3        o0404(.A(ori_ori_n138_), .B(ori_ori_n135_), .C(g), .Y(ori_ori_n433_));
  AOI220     o0405(.A0(ori_ori_n433_), .A1(ori_ori_n52_), .B0(ori_ori_n432_), .B1(ori_ori_n430_), .Y(ori_ori_n434_));
  INV        o0406(.A(ori_ori_n434_), .Y(ori_ori_n435_));
  AN3        o0407(.A(j), .B(h), .C(g), .Y(ori_ori_n436_));
  NO2        o0408(.A(ori_ori_n116_), .B(c), .Y(ori_ori_n437_));
  NA3        o0409(.A(ori_ori_n437_), .B(ori_ori_n436_), .C(ori_ori_n341_), .Y(ori_ori_n438_));
  NA3        o0410(.A(f), .B(d), .C(b), .Y(ori_ori_n439_));
  NO4        o0411(.A(ori_ori_n439_), .B(ori_ori_n138_), .C(ori_ori_n135_), .D(g), .Y(ori_ori_n440_));
  INV        o0412(.A(ori_ori_n438_), .Y(ori_ori_n441_));
  NO4        o0413(.A(ori_ori_n441_), .B(ori_ori_n435_), .C(ori_ori_n428_), .D(ori_ori_n422_), .Y(ori_ori_n442_));
  AN4        o0414(.A(ori_ori_n442_), .B(ori_ori_n414_), .C(ori_ori_n401_), .D(ori_ori_n396_), .Y(ori_ori_n443_));
  INV        o0415(.A(k), .Y(ori_ori_n444_));
  NA4        o0416(.A(ori_ori_n289_), .B(g), .C(ori_ori_n143_), .D(ori_ori_n92_), .Y(ori_ori_n445_));
  NAi32      o0417(.An(h), .Bn(f), .C(g), .Y(ori_ori_n446_));
  NAi41      o0418(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n447_));
  OAI210     o0419(.A0(ori_ori_n399_), .A1(n), .B0(ori_ori_n447_), .Y(ori_ori_n448_));
  NA2        o0420(.A(ori_ori_n448_), .B(m), .Y(ori_ori_n449_));
  OR2        o0421(.A(ori_ori_n449_), .B(ori_ori_n446_), .Y(ori_ori_n450_));
  NO3        o0422(.A(ori_ori_n446_), .B(ori_ori_n58_), .C(ori_ori_n59_), .Y(ori_ori_n451_));
  NAi31      o0423(.An(ori_ori_n451_), .B(ori_ori_n450_), .C(ori_ori_n445_), .Y(ori_ori_n452_));
  NAi31      o0424(.An(f), .B(h), .C(g), .Y(ori_ori_n453_));
  NO2        o0425(.A(n), .B(c), .Y(ori_ori_n454_));
  NA3        o0426(.A(ori_ori_n454_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n455_));
  NOi32      o0427(.An(e), .Bn(a), .C(d), .Y(ori_ori_n456_));
  AOI210     o0428(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n456_), .Y(ori_ori_n457_));
  NO2        o0429(.A(ori_ori_n195_), .B(ori_ori_n71_), .Y(ori_ori_n458_));
  AOI210     o0430(.A0(ori_ori_n452_), .A1(l), .B0(ori_ori_n458_), .Y(ori_ori_n459_));
  NO3        o0431(.A(ori_ori_n227_), .B(ori_ori_n54_), .C(n), .Y(ori_ori_n460_));
  NA3        o0432(.A(ori_ori_n379_), .B(ori_ori_n133_), .C(ori_ori_n132_), .Y(ori_ori_n461_));
  NA2        o0433(.A(ori_ori_n343_), .B(ori_ori_n182_), .Y(ori_ori_n462_));
  NA2        o0434(.A(ori_ori_n60_), .B(ori_ori_n92_), .Y(ori_ori_n463_));
  INV        o0435(.A(ori_ori_n463_), .Y(ori_ori_n464_));
  AOI220     o0436(.A0(ori_ori_n464_), .A1(ori_ori_n404_), .B0(ori_ori_n461_), .B1(ori_ori_n460_), .Y(ori_ori_n465_));
  NO2        o0437(.A(ori_ori_n465_), .B(ori_ori_n71_), .Y(ori_ori_n466_));
  NA3        o0438(.A(ori_ori_n417_), .B(ori_ori_n243_), .C(ori_ori_n40_), .Y(ori_ori_n467_));
  NOi32      o0439(.An(e), .Bn(c), .C(f), .Y(ori_ori_n468_));
  INV        o0440(.A(ori_ori_n167_), .Y(ori_ori_n469_));
  AOI220     o0441(.A0(ori_ori_n469_), .A1(ori_ori_n286_), .B0(ori_ori_n468_), .B1(ori_ori_n137_), .Y(ori_ori_n470_));
  NA3        o0442(.A(ori_ori_n470_), .B(ori_ori_n467_), .C(ori_ori_n140_), .Y(ori_ori_n471_));
  AOI210     o0443(.A0(ori_ori_n403_), .A1(ori_ori_n290_), .B0(ori_ori_n220_), .Y(ori_ori_n472_));
  NAi21      o0444(.An(k), .B(h), .Y(ori_ori_n473_));
  NO2        o0445(.A(ori_ori_n473_), .B(ori_ori_n204_), .Y(ori_ori_n474_));
  NA2        o0446(.A(ori_ori_n474_), .B(j), .Y(ori_ori_n475_));
  OR2        o0447(.A(ori_ori_n475_), .B(ori_ori_n449_), .Y(ori_ori_n476_));
  NOi31      o0448(.An(m), .B(n), .C(k), .Y(ori_ori_n477_));
  NA2        o0449(.A(j), .B(ori_ori_n477_), .Y(ori_ori_n478_));
  AOI210     o0450(.A0(ori_ori_n290_), .A1(ori_ori_n266_), .B0(ori_ori_n220_), .Y(ori_ori_n479_));
  NAi21      o0451(.An(ori_ori_n478_), .B(ori_ori_n479_), .Y(ori_ori_n480_));
  NA2        o0452(.A(ori_ori_n480_), .B(ori_ori_n476_), .Y(ori_ori_n481_));
  NA2        o0453(.A(ori_ori_n87_), .B(m), .Y(ori_ori_n482_));
  NO2        o0454(.A(ori_ori_n398_), .B(ori_ori_n138_), .Y(ori_ori_n483_));
  NA3        o0455(.A(ori_ori_n418_), .B(ori_ori_n206_), .C(ori_ori_n114_), .Y(ori_ori_n484_));
  NA2        o0456(.A(ori_ori_n377_), .B(ori_ori_n128_), .Y(ori_ori_n485_));
  NO3        o0457(.A(ori_ori_n287_), .B(ori_ori_n485_), .C(ori_ori_n71_), .Y(ori_ori_n486_));
  AOI210     o0458(.A0(ori_ori_n484_), .A1(ori_ori_n483_), .B0(ori_ori_n486_), .Y(ori_ori_n487_));
  AN3        o0459(.A(f), .B(d), .C(b), .Y(ori_ori_n488_));
  OAI210     o0460(.A0(ori_ori_n488_), .A1(ori_ori_n102_), .B0(n), .Y(ori_ori_n489_));
  NA3        o0461(.A(ori_ori_n377_), .B(ori_ori_n128_), .C(ori_ori_n170_), .Y(ori_ori_n490_));
  AOI210     o0462(.A0(ori_ori_n489_), .A1(ori_ori_n183_), .B0(ori_ori_n490_), .Y(ori_ori_n491_));
  NAi31      o0463(.An(m), .B(n), .C(k), .Y(ori_ori_n492_));
  NA2        o0464(.A(ori_ori_n491_), .B(j), .Y(ori_ori_n493_));
  NA2        o0465(.A(ori_ori_n493_), .B(ori_ori_n487_), .Y(ori_ori_n494_));
  NO4        o0466(.A(ori_ori_n494_), .B(ori_ori_n481_), .C(ori_ori_n471_), .D(ori_ori_n466_), .Y(ori_ori_n495_));
  NA2        o0467(.A(ori_ori_n274_), .B(ori_ori_n131_), .Y(ori_ori_n496_));
  NAi31      o0468(.An(g), .B(h), .C(f), .Y(ori_ori_n497_));
  OA210      o0469(.A0(ori_ori_n399_), .A1(n), .B0(ori_ori_n447_), .Y(ori_ori_n498_));
  NA3        o0470(.A(ori_ori_n307_), .B(ori_ori_n95_), .C(ori_ori_n69_), .Y(ori_ori_n499_));
  OAI210     o0471(.A0(ori_ori_n498_), .A1(ori_ori_n75_), .B0(ori_ori_n499_), .Y(ori_ori_n500_));
  INV        o0472(.A(ori_ori_n500_), .Y(ori_ori_n501_));
  AOI210     o0473(.A0(ori_ori_n501_), .A1(ori_ori_n496_), .B0(ori_ori_n394_), .Y(ori_ori_n502_));
  OR2        o0474(.A(ori_ori_n58_), .B(ori_ori_n59_), .Y(ori_ori_n503_));
  AN2        o0475(.A(h), .B(f), .Y(ori_ori_n504_));
  NA2        o0476(.A(ori_ori_n504_), .B(ori_ori_n35_), .Y(ori_ori_n505_));
  NO2        o0477(.A(ori_ori_n505_), .B(ori_ori_n347_), .Y(ori_ori_n506_));
  AOI210     o0478(.A0(ori_ori_n429_), .A1(ori_ori_n312_), .B0(ori_ori_n43_), .Y(ori_ori_n507_));
  NO2        o0479(.A(ori_ori_n197_), .B(f), .Y(ori_ori_n508_));
  INV        o0480(.A(ori_ori_n104_), .Y(ori_ori_n509_));
  AOI220     o0481(.A0(ori_ori_n509_), .A1(ori_ori_n397_), .B0(e), .B1(ori_ori_n92_), .Y(ori_ori_n510_));
  OA220      o0482(.A0(ori_ori_n510_), .A1(ori_ori_n415_), .B0(ori_ori_n258_), .B1(ori_ori_n90_), .Y(ori_ori_n511_));
  INV        o0483(.A(ori_ori_n511_), .Y(ori_ori_n512_));
  NO3        o0484(.A(ori_ori_n297_), .B(ori_ori_n154_), .C(ori_ori_n153_), .Y(ori_ori_n513_));
  NA2        o0485(.A(ori_ori_n513_), .B(ori_ori_n182_), .Y(ori_ori_n514_));
  NA3        o0486(.A(ori_ori_n514_), .B(ori_ori_n199_), .C(j), .Y(ori_ori_n515_));
  NO3        o0487(.A(ori_ori_n343_), .B(ori_ori_n135_), .C(i), .Y(ori_ori_n516_));
  NA2        o0488(.A(ori_ori_n346_), .B(ori_ori_n69_), .Y(ori_ori_n517_));
  NA2        o0489(.A(ori_ori_n515_), .B(ori_ori_n295_), .Y(ori_ori_n518_));
  NO4        o0490(.A(ori_ori_n518_), .B(ori_ori_n512_), .C(ori_ori_n506_), .D(ori_ori_n502_), .Y(ori_ori_n519_));
  NA4        o0491(.A(ori_ori_n519_), .B(ori_ori_n495_), .C(ori_ori_n459_), .D(ori_ori_n443_), .Y(ori08));
  NO2        o0492(.A(k), .B(h), .Y(ori_ori_n521_));
  AO210      o0493(.A0(ori_ori_n197_), .A1(ori_ori_n332_), .B0(ori_ori_n521_), .Y(ori_ori_n522_));
  NO2        o0494(.A(ori_ori_n522_), .B(ori_ori_n219_), .Y(ori_ori_n523_));
  NA2        o0495(.A(ori_ori_n468_), .B(ori_ori_n69_), .Y(ori_ori_n524_));
  INV        o0496(.A(ori_ori_n364_), .Y(ori_ori_n525_));
  NA2        o0497(.A(ori_ori_n69_), .B(ori_ori_n89_), .Y(ori_ori_n526_));
  NO2        o0498(.A(ori_ori_n526_), .B(ori_ori_n51_), .Y(ori_ori_n527_));
  NO3        o0499(.A(ori_ori_n272_), .B(ori_ori_n91_), .C(ori_ori_n170_), .Y(ori_ori_n528_));
  NA2        o0500(.A(ori_ori_n439_), .B(ori_ori_n183_), .Y(ori_ori_n529_));
  NA2        o0501(.A(ori_ori_n528_), .B(ori_ori_n527_), .Y(ori_ori_n530_));
  AOI210     o0502(.A0(ori_ori_n439_), .A1(ori_ori_n125_), .B0(ori_ori_n69_), .Y(ori_ori_n531_));
  NA4        o0503(.A(ori_ori_n172_), .B(ori_ori_n109_), .C(ori_ori_n39_), .D(h), .Y(ori_ori_n532_));
  AN2        o0504(.A(l), .B(k), .Y(ori_ori_n533_));
  NA3        o0505(.A(ori_ori_n533_), .B(ori_ori_n87_), .C(ori_ori_n59_), .Y(ori_ori_n534_));
  NA2        o0506(.A(ori_ori_n532_), .B(ori_ori_n534_), .Y(ori_ori_n535_));
  NA2        o0507(.A(ori_ori_n535_), .B(ori_ori_n531_), .Y(ori_ori_n536_));
  NA4        o0508(.A(ori_ori_n536_), .B(ori_ori_n530_), .C(ori_ori_n525_), .D(ori_ori_n250_), .Y(ori_ori_n537_));
  NO4        o0509(.A(ori_ori_n135_), .B(ori_ori_n285_), .C(ori_ori_n91_), .D(g), .Y(ori_ori_n538_));
  NA2        o0510(.A(ori_ori_n538_), .B(ori_ori_n529_), .Y(ori_ori_n539_));
  NA2        o0511(.A(ori_ori_n469_), .B(ori_ori_n247_), .Y(ori_ori_n540_));
  NA2        o0512(.A(ori_ori_n540_), .B(ori_ori_n539_), .Y(ori_ori_n541_));
  NO3        o0513(.A(ori_ori_n227_), .B(ori_ori_n103_), .C(ori_ori_n37_), .Y(ori_ori_n542_));
  NAi21      o0514(.An(ori_ori_n542_), .B(ori_ori_n534_), .Y(ori_ori_n543_));
  NA2        o0515(.A(ori_ori_n522_), .B(ori_ori_n106_), .Y(ori_ori_n544_));
  AOI220     o0516(.A0(ori_ori_n544_), .A1(ori_ori_n296_), .B0(ori_ori_n543_), .B1(ori_ori_n62_), .Y(ori_ori_n545_));
  INV        o0517(.A(ori_ori_n545_), .Y(ori_ori_n546_));
  NA3        o0518(.A(ori_ori_n514_), .B(ori_ori_n236_), .C(ori_ori_n277_), .Y(ori_ori_n547_));
  NA3        o0519(.A(m), .B(l), .C(k), .Y(ori_ori_n548_));
  NO2        o0520(.A(ori_ori_n499_), .B(ori_ori_n548_), .Y(ori_ori_n549_));
  INV        o0521(.A(ori_ori_n549_), .Y(ori_ori_n550_));
  NA2        o0522(.A(ori_ori_n550_), .B(ori_ori_n547_), .Y(ori_ori_n551_));
  NO4        o0523(.A(ori_ori_n551_), .B(ori_ori_n546_), .C(ori_ori_n541_), .D(ori_ori_n537_), .Y(ori_ori_n552_));
  NO2        o0524(.A(ori_ori_n290_), .B(ori_ori_n392_), .Y(ori_ori_n553_));
  AOI210     o0525(.A0(ori_ori_n553_), .A1(ori_ori_n92_), .B0(ori_ori_n372_), .Y(ori_ori_n554_));
  INV        o0526(.A(ori_ori_n554_), .Y(ori_ori_n555_));
  NA2        o0527(.A(ori_ori_n533_), .B(ori_ori_n59_), .Y(ori_ori_n556_));
  NO4        o0528(.A(ori_ori_n513_), .B(ori_ori_n135_), .C(n), .D(i), .Y(ori_ori_n557_));
  NA2        o0529(.A(h), .B(f), .Y(ori_ori_n558_));
  NO2        o0530(.A(ori_ori_n558_), .B(ori_ori_n192_), .Y(ori_ori_n559_));
  NO3        o0531(.A(ori_ori_n559_), .B(ori_ori_n557_), .C(ori_ori_n516_), .Y(ori_ori_n560_));
  NO2        o0532(.A(ori_ori_n560_), .B(ori_ori_n556_), .Y(ori_ori_n561_));
  AOI210     o0533(.A0(ori_ori_n555_), .A1(l), .B0(ori_ori_n561_), .Y(ori_ori_n562_));
  NA2        o0534(.A(ori_ori_n66_), .B(l), .Y(ori_ori_n563_));
  OR2        o0535(.A(ori_ori_n563_), .B(ori_ori_n449_), .Y(ori_ori_n564_));
  NO3        o0536(.A(ori_ori_n120_), .B(ori_ori_n43_), .C(ori_ori_n89_), .Y(ori_ori_n565_));
  AOI210     o0537(.A0(ori_ori_n397_), .A1(n), .B0(ori_ori_n417_), .Y(ori_ori_n566_));
  NA2        o0538(.A(ori_ori_n566_), .B(ori_ori_n420_), .Y(ori_ori_n567_));
  NO3        o0539(.A(ori_ori_n135_), .B(ori_ori_n285_), .C(ori_ori_n91_), .Y(ori_ori_n568_));
  AOI220     o0540(.A0(ori_ori_n568_), .A1(ori_ori_n193_), .B0(ori_ori_n462_), .B1(ori_ori_n224_), .Y(ori_ori_n569_));
  NAi31      o0541(.An(ori_ori_n457_), .B(ori_ori_n77_), .C(ori_ori_n69_), .Y(ori_ori_n570_));
  NA2        o0542(.A(ori_ori_n570_), .B(ori_ori_n569_), .Y(ori_ori_n571_));
  NA2        o0543(.A(ori_ori_n542_), .B(ori_ori_n531_), .Y(ori_ori_n572_));
  NO2        o0544(.A(ori_ori_n548_), .B(ori_ori_n75_), .Y(ori_ori_n573_));
  INV        o0545(.A(ori_ori_n572_), .Y(ori_ori_n574_));
  OR2        o0546(.A(ori_ori_n574_), .B(ori_ori_n571_), .Y(ori_ori_n575_));
  NA3        o0547(.A(ori_ori_n566_), .B(ori_ori_n420_), .C(ori_ori_n419_), .Y(ori_ori_n576_));
  NA4        o0548(.A(ori_ori_n576_), .B(ori_ori_n172_), .C(ori_ori_n332_), .D(ori_ori_n33_), .Y(ori_ori_n577_));
  NO3        o0549(.A(ori_ori_n358_), .B(ori_ori_n316_), .C(f), .Y(ori_ori_n578_));
  NA2        o0550(.A(ori_ori_n578_), .B(ori_ori_n203_), .Y(ori_ori_n579_));
  NA3        o0551(.A(f), .B(ori_ori_n213_), .C(h), .Y(ori_ori_n580_));
  NOi21      o0552(.An(ori_ori_n507_), .B(ori_ori_n580_), .Y(ori_ori_n581_));
  NO2        o0553(.A(ori_ori_n563_), .B(ori_ori_n503_), .Y(ori_ori_n582_));
  INV        o0554(.A(ori_ori_n582_), .Y(ori_ori_n583_));
  NAi41      o0555(.An(ori_ori_n581_), .B(ori_ori_n583_), .C(ori_ori_n579_), .D(ori_ori_n577_), .Y(ori_ori_n584_));
  BUFFER     o0556(.A(ori_ori_n573_), .Y(ori_ori_n585_));
  NA2        o0557(.A(ori_ori_n585_), .B(ori_ori_n187_), .Y(ori_ori_n586_));
  NO2        o0558(.A(ori_ori_n498_), .B(ori_ori_n59_), .Y(ori_ori_n587_));
  AOI210     o0559(.A0(ori_ori_n578_), .A1(ori_ori_n587_), .B0(ori_ori_n238_), .Y(ori_ori_n588_));
  OAI210     o0560(.A0(ori_ori_n548_), .A1(ori_ori_n497_), .B0(ori_ori_n386_), .Y(ori_ori_n589_));
  NA3        o0561(.A(ori_ori_n196_), .B(ori_ori_n53_), .C(b), .Y(ori_ori_n590_));
  AOI220     o0562(.A0(ori_ori_n454_), .A1(ori_ori_n29_), .B0(ori_ori_n346_), .B1(ori_ori_n69_), .Y(ori_ori_n591_));
  NA2        o0563(.A(ori_ori_n591_), .B(ori_ori_n590_), .Y(ori_ori_n592_));
  NA2        o0564(.A(ori_ori_n592_), .B(ori_ori_n589_), .Y(ori_ori_n593_));
  NA3        o0565(.A(ori_ori_n593_), .B(ori_ori_n588_), .C(ori_ori_n586_), .Y(ori_ori_n594_));
  NOi41      o0566(.An(ori_ori_n564_), .B(ori_ori_n594_), .C(ori_ori_n584_), .D(ori_ori_n575_), .Y(ori_ori_n595_));
  NO3        o0567(.A(ori_ori_n244_), .B(ori_ori_n220_), .C(ori_ori_n91_), .Y(ori_ori_n596_));
  NA2        o0568(.A(ori_ori_n596_), .B(ori_ori_n567_), .Y(ori_ori_n597_));
  NO3        o0569(.A(ori_ori_n392_), .B(ori_ori_n78_), .C(h), .Y(ori_ori_n598_));
  NA2        o0570(.A(ori_ori_n598_), .B(ori_ori_n527_), .Y(ori_ori_n599_));
  NA2        o0571(.A(ori_ori_n599_), .B(ori_ori_n597_), .Y(ori_ori_n600_));
  OR2        o0572(.A(ori_ori_n497_), .B(ori_ori_n76_), .Y(ori_ori_n601_));
  NOi31      o0573(.An(b), .B(d), .C(a), .Y(ori_ori_n602_));
  NO2        o0574(.A(ori_ori_n418_), .B(ori_ori_n69_), .Y(ori_ori_n603_));
  NA2        o0575(.A(ori_ori_n596_), .B(ori_ori_n603_), .Y(ori_ori_n604_));
  OAI210     o0576(.A0(ori_ori_n532_), .A1(ori_ori_n287_), .B0(ori_ori_n604_), .Y(ori_ori_n605_));
  NO2        o0577(.A(ori_ori_n513_), .B(n), .Y(ori_ori_n606_));
  NA2        o0578(.A(ori_ori_n606_), .B(ori_ori_n523_), .Y(ori_ori_n607_));
  NO2        o0579(.A(ori_ori_n230_), .B(ori_ori_n186_), .Y(ori_ori_n608_));
  OAI210     o0580(.A0(ori_ori_n80_), .A1(ori_ori_n77_), .B0(ori_ori_n608_), .Y(ori_ori_n609_));
  INV        o0581(.A(ori_ori_n609_), .Y(ori_ori_n610_));
  NA2        o0582(.A(ori_ori_n538_), .B(ori_ori_n249_), .Y(ori_ori_n611_));
  NA2        o0583(.A(ori_ori_n451_), .B(j), .Y(ori_ori_n612_));
  AN2        o0584(.A(ori_ori_n612_), .B(ori_ori_n611_), .Y(ori_ori_n613_));
  NAi31      o0585(.An(ori_ori_n610_), .B(ori_ori_n613_), .C(ori_ori_n607_), .Y(ori_ori_n614_));
  NO3        o0586(.A(ori_ori_n614_), .B(ori_ori_n605_), .C(ori_ori_n600_), .Y(ori_ori_n615_));
  NA4        o0587(.A(ori_ori_n615_), .B(ori_ori_n595_), .C(ori_ori_n562_), .D(ori_ori_n552_), .Y(ori09));
  INV        o0588(.A(ori_ori_n96_), .Y(ori_ori_n617_));
  NA2        o0589(.A(f), .B(e), .Y(ori_ori_n618_));
  NA2        o0590(.A(l), .B(g), .Y(ori_ori_n619_));
  NO2        o0591(.A(ori_ori_n619_), .B(ori_ori_n618_), .Y(ori_ori_n620_));
  NA2        o0592(.A(ori_ori_n326_), .B(e), .Y(ori_ori_n621_));
  NO2        o0593(.A(ori_ori_n621_), .B(ori_ori_n379_), .Y(ori_ori_n622_));
  AOI210     o0594(.A0(ori_ori_n620_), .A1(ori_ori_n617_), .B0(ori_ori_n622_), .Y(ori_ori_n623_));
  NA2        o0595(.A(ori_ori_n72_), .B(g), .Y(ori_ori_n624_));
  INV        o0596(.A(ori_ori_n241_), .Y(ori_ori_n625_));
  NO2        o0597(.A(ori_ori_n100_), .B(ori_ori_n98_), .Y(ori_ori_n626_));
  NOi31      o0598(.An(k), .B(m), .C(l), .Y(ori_ori_n627_));
  NO2        o0599(.A(ori_ori_n243_), .B(ori_ori_n627_), .Y(ori_ori_n628_));
  AOI210     o0600(.A0(ori_ori_n628_), .A1(ori_ori_n626_), .B0(ori_ori_n453_), .Y(ori_ori_n629_));
  NA2        o0601(.A(ori_ori_n590_), .B(ori_ori_n234_), .Y(ori_ori_n630_));
  NA2        o0602(.A(ori_ori_n245_), .B(m), .Y(ori_ori_n631_));
  OAI210     o0603(.A0(ori_ori_n163_), .A1(ori_ori_n169_), .B0(ori_ori_n631_), .Y(ori_ori_n632_));
  AOI220     o0604(.A0(ori_ori_n632_), .A1(ori_ori_n630_), .B0(ori_ori_n629_), .B1(ori_ori_n625_), .Y(ori_ori_n633_));
  NA2        o0605(.A(ori_ori_n522_), .B(ori_ori_n106_), .Y(ori_ori_n634_));
  NA3        o0606(.A(ori_ori_n634_), .B(ori_ori_n151_), .C(e), .Y(ori_ori_n635_));
  NA4        o0607(.A(ori_ori_n635_), .B(ori_ori_n633_), .C(ori_ori_n470_), .D(ori_ori_n67_), .Y(ori_ori_n636_));
  NO2        o0608(.A(ori_ori_n446_), .B(ori_ori_n369_), .Y(ori_ori_n637_));
  NA2        o0609(.A(ori_ori_n637_), .B(ori_ori_n151_), .Y(ori_ori_n638_));
  NA2        o0610(.A(f), .B(m), .Y(ori_ori_n639_));
  NO2        o0611(.A(ori_ori_n639_), .B(ori_ori_n46_), .Y(ori_ori_n640_));
  NOi32      o0612(.An(g), .Bn(f), .C(d), .Y(ori_ori_n641_));
  NA4        o0613(.A(ori_ori_n641_), .B(ori_ori_n454_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n642_));
  INV        o0614(.A(ori_ori_n642_), .Y(ori_ori_n643_));
  AOI210     o0615(.A0(ori_ori_n640_), .A1(ori_ori_n410_), .B0(ori_ori_n643_), .Y(ori_ori_n644_));
  AN2        o0616(.A(f), .B(d), .Y(ori_ori_n645_));
  NA3        o0617(.A(ori_ori_n352_), .B(ori_ori_n645_), .C(ori_ori_n69_), .Y(ori_ori_n646_));
  NAi31      o0618(.An(ori_ori_n363_), .B(ori_ori_n644_), .C(ori_ori_n638_), .Y(ori_ori_n647_));
  NO3        o0619(.A(ori_ori_n104_), .B(ori_ori_n232_), .C(ori_ori_n121_), .Y(ori_ori_n648_));
  NO2        o0620(.A(ori_ori_n492_), .B(ori_ori_n232_), .Y(ori_ori_n649_));
  AN2        o0621(.A(ori_ori_n649_), .B(ori_ori_n508_), .Y(ori_ori_n650_));
  NO2        o0622(.A(ori_ori_n650_), .B(ori_ori_n648_), .Y(ori_ori_n651_));
  NO2        o0623(.A(ori_ori_n646_), .B(ori_ori_n314_), .Y(ori_ori_n652_));
  NOi21      o0624(.An(ori_ori_n178_), .B(ori_ori_n652_), .Y(ori_ori_n653_));
  NA2        o0625(.A(c), .B(ori_ori_n93_), .Y(ori_ori_n654_));
  NO2        o0626(.A(ori_ori_n654_), .B(ori_ori_n301_), .Y(ori_ori_n655_));
  NA3        o0627(.A(ori_ori_n655_), .B(ori_ori_n378_), .C(f), .Y(ori_ori_n656_));
  NA3        o0628(.A(ori_ori_n656_), .B(ori_ori_n653_), .C(ori_ori_n651_), .Y(ori_ori_n657_));
  NO3        o0629(.A(ori_ori_n657_), .B(ori_ori_n647_), .C(ori_ori_n636_), .Y(ori_ori_n658_));
  OR2        o0630(.A(ori_ori_n646_), .B(ori_ori_n59_), .Y(ori_ori_n659_));
  NA2        o0631(.A(l), .B(g), .Y(ori_ori_n660_));
  AOI210     o0632(.A0(ori_ori_n660_), .A1(ori_ori_n214_), .B0(ori_ori_n659_), .Y(ori_ori_n661_));
  NO2        o0633(.A(ori_ori_n234_), .B(ori_ori_n624_), .Y(ori_ori_n662_));
  NO2        o0634(.A(ori_ori_n106_), .B(ori_ori_n104_), .Y(ori_ori_n663_));
  NO2        o0635(.A(ori_ori_n182_), .B(ori_ori_n179_), .Y(ori_ori_n664_));
  AOI220     o0636(.A0(ori_ori_n664_), .A1(ori_ori_n181_), .B0(ori_ori_n222_), .B1(ori_ori_n663_), .Y(ori_ori_n665_));
  NO2        o0637(.A(ori_ori_n314_), .B(ori_ori_n618_), .Y(ori_ori_n666_));
  NA2        o0638(.A(ori_ori_n666_), .B(ori_ori_n425_), .Y(ori_ori_n667_));
  NA2        o0639(.A(ori_ori_n667_), .B(ori_ori_n665_), .Y(ori_ori_n668_));
  NA2        o0640(.A(e), .B(d), .Y(ori_ori_n669_));
  OAI220     o0641(.A0(ori_ori_n669_), .A1(c), .B0(ori_ori_n230_), .B1(d), .Y(ori_ori_n670_));
  NA3        o0642(.A(ori_ori_n670_), .B(ori_ori_n337_), .C(ori_ori_n377_), .Y(ori_ori_n671_));
  AOI210     o0643(.A0(ori_ori_n382_), .A1(ori_ori_n142_), .B0(ori_ori_n182_), .Y(ori_ori_n672_));
  AOI210     o0644(.A0(ori_ori_n469_), .A1(ori_ori_n247_), .B0(ori_ori_n672_), .Y(ori_ori_n673_));
  NA2        o0645(.A(ori_ori_n673_), .B(ori_ori_n671_), .Y(ori_ori_n674_));
  NO4        o0646(.A(ori_ori_n674_), .B(ori_ori_n668_), .C(ori_ori_n662_), .D(ori_ori_n661_), .Y(ori_ori_n675_));
  OR2        o0647(.A(ori_ori_n524_), .B(ori_ori_n173_), .Y(ori_ori_n676_));
  NO2        o0648(.A(ori_ori_n621_), .B(ori_ori_n132_), .Y(ori_ori_n677_));
  INV        o0649(.A(ori_ori_n677_), .Y(ori_ori_n678_));
  AN2        o0650(.A(ori_ori_n137_), .B(f), .Y(ori_ori_n679_));
  OAI210     o0651(.A0(ori_ori_n679_), .A1(ori_ori_n339_), .B0(ori_ori_n670_), .Y(ori_ori_n680_));
  NO2        o0652(.A(ori_ori_n320_), .B(ori_ori_n56_), .Y(ori_ori_n681_));
  NA2        o0653(.A(ori_ori_n681_), .B(ori_ori_n527_), .Y(ori_ori_n682_));
  AN4        o0654(.A(ori_ori_n682_), .B(ori_ori_n680_), .C(ori_ori_n678_), .D(ori_ori_n676_), .Y(ori_ori_n683_));
  NA4        o0655(.A(ori_ori_n683_), .B(ori_ori_n675_), .C(ori_ori_n658_), .D(ori_ori_n623_), .Y(ori12));
  NO2        o0656(.A(ori_ori_n335_), .B(c), .Y(ori_ori_n685_));
  NO4        o0657(.A(ori_ori_n325_), .B(ori_ori_n197_), .C(ori_ori_n444_), .D(ori_ori_n170_), .Y(ori_ori_n686_));
  NA2        o0658(.A(ori_ori_n686_), .B(ori_ori_n685_), .Y(ori_ori_n687_));
  NA2        o0659(.A(ori_ori_n410_), .B(ori_ori_n681_), .Y(ori_ori_n688_));
  NO2        o0660(.A(ori_ori_n335_), .B(ori_ori_n93_), .Y(ori_ori_n689_));
  NO2        o0661(.A(ori_ori_n626_), .B(ori_ori_n252_), .Y(ori_ori_n690_));
  NO2        o0662(.A(ori_ori_n497_), .B(ori_ori_n272_), .Y(ori_ori_n691_));
  AOI220     o0663(.A0(ori_ori_n691_), .A1(ori_ori_n408_), .B0(ori_ori_n690_), .B1(ori_ori_n689_), .Y(ori_ori_n692_));
  NA4        o0664(.A(ori_ori_n692_), .B(ori_ori_n688_), .C(ori_ori_n687_), .D(ori_ori_n324_), .Y(ori_ori_n693_));
  AOI210     o0665(.A0(ori_ori_n184_), .A1(ori_ori_n240_), .B0(ori_ori_n160_), .Y(ori_ori_n694_));
  BUFFER     o0666(.A(ori_ori_n686_), .Y(ori_ori_n695_));
  AOI210     o0667(.A0(ori_ori_n237_), .A1(ori_ori_n283_), .B0(ori_ori_n170_), .Y(ori_ori_n696_));
  OAI210     o0668(.A0(ori_ori_n696_), .A1(ori_ori_n695_), .B0(ori_ori_n297_), .Y(ori_ori_n697_));
  NO2        o0669(.A(ori_ori_n482_), .B(ori_ori_n204_), .Y(ori_ori_n698_));
  NA2        o0670(.A(ori_ori_n608_), .B(ori_ori_n698_), .Y(ori_ori_n699_));
  NO2        o0671(.A(ori_ori_n120_), .B(ori_ori_n186_), .Y(ori_ori_n700_));
  NA3        o0672(.A(ori_ori_n700_), .B(ori_ori_n189_), .C(i), .Y(ori_ori_n701_));
  NA3        o0673(.A(ori_ori_n701_), .B(ori_ori_n699_), .C(ori_ori_n697_), .Y(ori_ori_n702_));
  NO3        o0674(.A(ori_ori_n104_), .B(ori_ori_n121_), .C(ori_ori_n170_), .Y(ori_ori_n703_));
  NA2        o0675(.A(ori_ori_n703_), .B(ori_ori_n397_), .Y(ori_ori_n704_));
  NA4        o0676(.A(ori_ori_n326_), .B(ori_ori_n318_), .C(ori_ori_n143_), .D(g), .Y(ori_ori_n705_));
  NA2        o0677(.A(ori_ori_n705_), .B(ori_ori_n704_), .Y(ori_ori_n706_));
  NO3        o0678(.A(ori_ori_n501_), .B(ori_ori_n76_), .C(ori_ori_n39_), .Y(ori_ori_n707_));
  NO4        o0679(.A(ori_ori_n707_), .B(ori_ori_n706_), .C(ori_ori_n702_), .D(ori_ori_n693_), .Y(ori_ori_n708_));
  NO2        o0680(.A(ori_ori_n264_), .B(ori_ori_n263_), .Y(ori_ori_n709_));
  NA2        o0681(.A(ori_ori_n447_), .B(ori_ori_n58_), .Y(ori_ori_n710_));
  NA2        o0682(.A(ori_ori_n418_), .B(ori_ori_n114_), .Y(ori_ori_n711_));
  NOi21      o0683(.An(ori_ori_n33_), .B(ori_ori_n492_), .Y(ori_ori_n712_));
  AOI220     o0684(.A0(ori_ori_n712_), .A1(ori_ori_n711_), .B0(ori_ori_n710_), .B1(ori_ori_n709_), .Y(ori_ori_n713_));
  INV        o0685(.A(ori_ori_n713_), .Y(ori_ori_n714_));
  INV        o0686(.A(ori_ori_n43_), .Y(ori_ori_n715_));
  NO2        o0687(.A(ori_ori_n375_), .B(ori_ori_n220_), .Y(ori_ori_n716_));
  INV        o0688(.A(ori_ori_n716_), .Y(ori_ori_n717_));
  NO2        o0689(.A(ori_ori_n717_), .B(ori_ori_n114_), .Y(ori_ori_n718_));
  INV        o0690(.A(ori_ori_n262_), .Y(ori_ori_n719_));
  NO3        o0691(.A(ori_ori_n719_), .B(ori_ori_n718_), .C(ori_ori_n714_), .Y(ori_ori_n720_));
  NA2        o0692(.A(ori_ori_n247_), .B(g), .Y(ori_ori_n721_));
  NA2        o0693(.A(ori_ori_n131_), .B(i), .Y(ori_ori_n722_));
  NA2        o0694(.A(ori_ori_n40_), .B(i), .Y(ori_ori_n723_));
  NO2        o0695(.A(ori_ori_n723_), .B(ori_ori_n1032_), .Y(ori_ori_n724_));
  INV        o0696(.A(ori_ori_n724_), .Y(ori_ori_n725_));
  NO2        o0697(.A(ori_ori_n114_), .B(ori_ori_n69_), .Y(ori_ori_n726_));
  OR2        o0698(.A(ori_ori_n726_), .B(ori_ori_n417_), .Y(ori_ori_n727_));
  NA2        o0699(.A(ori_ori_n418_), .B(ori_ori_n275_), .Y(ori_ori_n728_));
  AOI210     o0700(.A0(ori_ori_n728_), .A1(n), .B0(ori_ori_n727_), .Y(ori_ori_n729_));
  OAI220     o0701(.A0(ori_ori_n729_), .A1(ori_ori_n721_), .B0(ori_ori_n725_), .B1(ori_ori_n234_), .Y(ori_ori_n730_));
  NA2        o0702(.A(ori_ori_n456_), .B(ori_ori_n92_), .Y(ori_ori_n731_));
  NA3        o0703(.A(f), .B(ori_ori_n94_), .C(g), .Y(ori_ori_n732_));
  AOI210     o0704(.A0(ori_ori_n505_), .A1(ori_ori_n732_), .B0(m), .Y(ori_ori_n733_));
  OAI210     o0705(.A0(ori_ori_n733_), .A1(ori_ori_n690_), .B0(ori_ori_n231_), .Y(ori_ori_n734_));
  INV        o0706(.A(ori_ori_n734_), .Y(ori_ori_n735_));
  NO2        o0707(.A(ori_ori_n272_), .B(ori_ori_n75_), .Y(ori_ori_n736_));
  OAI210     o0708(.A0(ori_ori_n736_), .A1(ori_ori_n698_), .B0(ori_ori_n187_), .Y(ori_ori_n737_));
  NA2        o0709(.A(ori_ori_n500_), .B(ori_ori_n72_), .Y(ori_ori_n738_));
  NO2        o0710(.A(ori_ori_n342_), .B(ori_ori_n170_), .Y(ori_ori_n739_));
  AOI220     o0711(.A0(ori_ori_n739_), .A1(ori_ori_n276_), .B0(c), .B1(ori_ori_n174_), .Y(ori_ori_n740_));
  AOI220     o0712(.A0(ori_ori_n691_), .A1(ori_ori_n700_), .B0(ori_ori_n448_), .B1(ori_ori_n74_), .Y(ori_ori_n741_));
  NA4        o0713(.A(ori_ori_n741_), .B(ori_ori_n740_), .C(ori_ori_n738_), .D(ori_ori_n737_), .Y(ori_ori_n742_));
  OAI210     o0714(.A0(ori_ori_n264_), .A1(ori_ori_n263_), .B0(ori_ori_n88_), .Y(ori_ori_n743_));
  NA2        o0715(.A(ori_ori_n743_), .B(ori_ori_n400_), .Y(ori_ori_n744_));
  NA2        o0716(.A(ori_ori_n733_), .B(ori_ori_n689_), .Y(ori_ori_n745_));
  NO3        o0717(.A(ori_ori_n1029_), .B(ori_ori_n43_), .C(ori_ori_n39_), .Y(ori_ori_n746_));
  AOI220     o0718(.A0(ori_ori_n746_), .A1(ori_ori_n472_), .B0(ori_ori_n483_), .B1(ori_ori_n397_), .Y(ori_ori_n747_));
  NA3        o0719(.A(ori_ori_n747_), .B(ori_ori_n745_), .C(ori_ori_n744_), .Y(ori_ori_n748_));
  NO4        o0720(.A(ori_ori_n748_), .B(ori_ori_n742_), .C(ori_ori_n735_), .D(ori_ori_n730_), .Y(ori_ori_n749_));
  NAi31      o0721(.An(ori_ori_n110_), .B(ori_ori_n309_), .C(n), .Y(ori_ori_n750_));
  NO3        o0722(.A(ori_ori_n98_), .B(ori_ori_n243_), .C(ori_ori_n627_), .Y(ori_ori_n751_));
  NO2        o0723(.A(ori_ori_n751_), .B(ori_ori_n750_), .Y(ori_ori_n752_));
  NO2        o0724(.A(ori_ori_n207_), .B(ori_ori_n110_), .Y(ori_ori_n753_));
  AOI210     o0725(.A0(ori_ori_n753_), .A1(ori_ori_n370_), .B0(ori_ori_n752_), .Y(ori_ori_n754_));
  NA2        o0726(.A(ori_ori_n364_), .B(i), .Y(ori_ori_n755_));
  NA2        o0727(.A(ori_ori_n755_), .B(ori_ori_n754_), .Y(ori_ori_n756_));
  NA2        o0728(.A(ori_ori_n182_), .B(ori_ori_n133_), .Y(ori_ori_n757_));
  NO3        o0729(.A(ori_ori_n224_), .B(ori_ori_n326_), .C(ori_ori_n137_), .Y(ori_ori_n758_));
  NOi31      o0730(.An(ori_ori_n757_), .B(ori_ori_n758_), .C(ori_ori_n170_), .Y(ori_ori_n759_));
  NAi21      o0731(.An(ori_ori_n418_), .B(ori_ori_n739_), .Y(ori_ori_n760_));
  INV        o0732(.A(ori_ori_n760_), .Y(ori_ori_n761_));
  NA2        o0733(.A(ori_ori_n694_), .B(ori_ori_n685_), .Y(ori_ori_n762_));
  NA2        o0734(.A(ori_ori_n762_), .B(ori_ori_n467_), .Y(ori_ori_n763_));
  OAI210     o0735(.A0(ori_ori_n694_), .A1(ori_ori_n686_), .B0(ori_ori_n757_), .Y(ori_ori_n764_));
  NA3        o0736(.A(ori_ori_n728_), .B(ori_ori_n360_), .C(ori_ori_n40_), .Y(ori_ori_n765_));
  INV        o0737(.A(ori_ori_n233_), .Y(ori_ori_n766_));
  NA3        o0738(.A(ori_ori_n766_), .B(ori_ori_n765_), .C(ori_ori_n764_), .Y(ori_ori_n767_));
  OR2        o0739(.A(ori_ori_n767_), .B(ori_ori_n763_), .Y(ori_ori_n768_));
  NO4        o0740(.A(ori_ori_n768_), .B(ori_ori_n761_), .C(ori_ori_n759_), .D(ori_ori_n756_), .Y(ori_ori_n769_));
  NA4        o0741(.A(ori_ori_n769_), .B(ori_ori_n749_), .C(ori_ori_n720_), .D(ori_ori_n708_), .Y(ori13));
  AN2        o0742(.A(d), .B(c), .Y(ori_ori_n771_));
  NA2        o0743(.A(ori_ori_n771_), .B(ori_ori_n93_), .Y(ori_ori_n772_));
  NAi32      o0744(.An(f), .Bn(e), .C(c), .Y(ori_ori_n773_));
  NO3        o0745(.A(m), .B(i), .C(h), .Y(ori_ori_n774_));
  NA3        o0746(.A(k), .B(j), .C(i), .Y(ori_ori_n775_));
  NO2        o0747(.A(f), .B(c), .Y(ori_ori_n776_));
  NOi21      o0748(.An(ori_ori_n776_), .B(ori_ori_n325_), .Y(ori_ori_n777_));
  AN3        o0749(.A(g), .B(f), .C(c), .Y(ori_ori_n778_));
  NA3        o0750(.A(l), .B(k), .C(j), .Y(ori_ori_n779_));
  NA2        o0751(.A(i), .B(h), .Y(ori_ori_n780_));
  NO3        o0752(.A(ori_ori_n780_), .B(ori_ori_n779_), .C(ori_ori_n104_), .Y(ori_ori_n781_));
  NO3        o0753(.A(ori_ori_n111_), .B(ori_ori_n212_), .C(ori_ori_n170_), .Y(ori_ori_n782_));
  NA3        o0754(.A(c), .B(b), .C(a), .Y(ori_ori_n783_));
  NO2        o0755(.A(ori_ori_n393_), .B(ori_ori_n453_), .Y(ori_ori_n784_));
  NA3        o0756(.A(ori_ori_n72_), .B(g), .C(ori_ori_n169_), .Y(ori_ori_n785_));
  NA4        o0757(.A(ori_ori_n436_), .B(m), .C(ori_ori_n91_), .D(ori_ori_n169_), .Y(ori_ori_n786_));
  NA2        o0758(.A(ori_ori_n786_), .B(ori_ori_n785_), .Y(ori_ori_n787_));
  NO3        o0759(.A(ori_ori_n787_), .B(ori_ori_n784_), .C(ori_ori_n743_), .Y(ori_ori_n788_));
  NOi21      o0760(.An(ori_ori_n601_), .B(ori_ori_n632_), .Y(ori_ori_n789_));
  OAI220     o0761(.A0(ori_ori_n789_), .A1(ori_ori_n517_), .B0(ori_ori_n788_), .B1(ori_ori_n447_), .Y(ori_ori_n790_));
  NOi31      o0762(.An(m), .B(n), .C(f), .Y(ori_ori_n791_));
  NA2        o0763(.A(ori_ori_n791_), .B(ori_ori_n45_), .Y(ori_ori_n792_));
  NO2        o0764(.A(ori_ori_n71_), .B(g), .Y(ori_ori_n793_));
  NO3        o0765(.A(ori_ori_n790_), .B(ori_ori_n610_), .C(ori_ori_n428_), .Y(ori_ori_n794_));
  NA2        o0766(.A(c), .B(b), .Y(ori_ori_n795_));
  NO2        o0767(.A(ori_ori_n526_), .B(ori_ori_n795_), .Y(ori_ori_n796_));
  INV        o0768(.A(ori_ori_n306_), .Y(ori_ori_n797_));
  OAI210     o0769(.A0(ori_ori_n797_), .A1(ori_ori_n640_), .B0(ori_ori_n796_), .Y(ori_ori_n798_));
  NA3        o0770(.A(ori_ori_n313_), .B(ori_ori_n423_), .C(f), .Y(ori_ori_n799_));
  INV        o0771(.A(ori_ori_n799_), .Y(ori_ori_n800_));
  NA2        o0772(.A(k), .B(g), .Y(ori_ori_n801_));
  NAi21      o0773(.An(f), .B(d), .Y(ori_ori_n802_));
  NO2        o0774(.A(ori_ori_n802_), .B(ori_ori_n783_), .Y(ori_ori_n803_));
  INV        o0775(.A(ori_ori_n803_), .Y(ori_ori_n804_));
  AOI210     o0776(.A0(ori_ori_n801_), .A1(ori_ori_n214_), .B0(ori_ori_n804_), .Y(ori_ori_n805_));
  AOI210     o0777(.A0(ori_ori_n805_), .A1(ori_ori_n92_), .B0(ori_ori_n800_), .Y(ori_ori_n806_));
  NA2        o0778(.A(ori_ori_n425_), .B(ori_ori_n303_), .Y(ori_ori_n807_));
  NA2        o0779(.A(ori_ori_n329_), .B(ori_ori_n803_), .Y(ori_ori_n808_));
  NO2        o0780(.A(ori_ori_n267_), .B(ori_ori_n266_), .Y(ori_ori_n809_));
  NAi31      o0781(.An(ori_ori_n809_), .B(ori_ori_n808_), .C(ori_ori_n807_), .Y(ori_ori_n810_));
  INV        o0782(.A(ori_ori_n810_), .Y(ori_ori_n811_));
  NA4        o0783(.A(ori_ori_n811_), .B(ori_ori_n806_), .C(ori_ori_n798_), .D(ori_ori_n794_), .Y(ori00));
  NA2        o0784(.A(ori_ori_n666_), .B(ori_ori_n700_), .Y(ori_ori_n813_));
  NA2        o0785(.A(ori_ori_n813_), .B(ori_ori_n744_), .Y(ori_ori_n814_));
  NA2        o0786(.A(ori_ori_n378_), .B(f), .Y(ori_ori_n815_));
  OAI210     o0787(.A0(ori_ori_n751_), .A1(ori_ori_n36_), .B0(ori_ori_n485_), .Y(ori_ori_n816_));
  NA3        o0788(.A(ori_ori_n816_), .B(ori_ori_n202_), .C(n), .Y(ori_ori_n817_));
  AOI210     o0789(.A0(ori_ori_n817_), .A1(ori_ori_n815_), .B0(ori_ori_n772_), .Y(ori_ori_n818_));
  NO2        o0790(.A(ori_ori_n818_), .B(ori_ori_n814_), .Y(ori_ori_n819_));
  NA3        o0791(.A(d), .B(ori_ori_n50_), .C(b), .Y(ori_ori_n820_));
  INV        o0792(.A(ori_ori_n438_), .Y(ori_ori_n821_));
  NO2        o0793(.A(ori_ori_n821_), .B(ori_ori_n809_), .Y(ori_ori_n822_));
  NO4        o0794(.A(ori_ori_n361_), .B(ori_ori_n255_), .C(ori_ori_n795_), .D(ori_ori_n53_), .Y(ori_ori_n823_));
  NA3        o0795(.A(ori_ori_n277_), .B(ori_ori_n177_), .C(g), .Y(ori_ori_n824_));
  OR2        o0796(.A(ori_ori_n824_), .B(ori_ori_n820_), .Y(ori_ori_n825_));
  NO2        o0797(.A(h), .B(g), .Y(ori_ori_n826_));
  AOI220     o0798(.A0(ori_ori_n228_), .A1(ori_ori_n193_), .B0(ori_ori_n139_), .B1(ori_ori_n118_), .Y(ori_ori_n827_));
  NA2        o0799(.A(ori_ori_n827_), .B(ori_ori_n825_), .Y(ori_ori_n828_));
  NO2        o0800(.A(ori_ori_n828_), .B(ori_ori_n823_), .Y(ori_ori_n829_));
  AOI210     o0801(.A0(ori_ori_n193_), .A1(ori_ori_n247_), .B0(ori_ori_n440_), .Y(ori_ori_n830_));
  NA2        o0802(.A(ori_ori_n830_), .B(ori_ori_n123_), .Y(ori_ori_n831_));
  NO2        o0803(.A(ori_ori_n188_), .B(ori_ori_n143_), .Y(ori_ori_n832_));
  NA2        o0804(.A(ori_ori_n832_), .B(ori_ori_n313_), .Y(ori_ori_n833_));
  INV        o0805(.A(ori_ori_n833_), .Y(ori_ori_n834_));
  NO2        o0806(.A(ori_ori_n834_), .B(ori_ori_n831_), .Y(ori_ori_n835_));
  AN3        o0807(.A(ori_ori_n835_), .B(ori_ori_n829_), .C(ori_ori_n822_), .Y(ori_ori_n836_));
  NA2        o0808(.A(ori_ori_n400_), .B(ori_ori_n83_), .Y(ori_ori_n837_));
  NA3        o0809(.A(ori_ori_n791_), .B(ori_ori_n456_), .C(h), .Y(ori_ori_n838_));
  NA2        o0810(.A(ori_ori_n838_), .B(ori_ori_n837_), .Y(ori_ori_n839_));
  NA4        o0811(.A(ori_ori_n488_), .B(k), .C(ori_ori_n177_), .D(ori_ori_n131_), .Y(ori_ori_n840_));
  NA2        o0812(.A(ori_ori_n425_), .B(ori_ori_n303_), .Y(ori_ori_n841_));
  NO2        o0813(.A(ori_ori_n173_), .B(ori_ori_n170_), .Y(ori_ori_n842_));
  NA2        o0814(.A(n), .B(e), .Y(ori_ori_n843_));
  NO2        o0815(.A(ori_ori_n843_), .B(ori_ori_n116_), .Y(ori_ori_n844_));
  AOI220     o0816(.A0(ori_ori_n844_), .A1(ori_ori_n208_), .B0(ori_ori_n625_), .B1(ori_ori_n842_), .Y(ori_ori_n845_));
  NA2        o0817(.A(ori_ori_n845_), .B(ori_ori_n841_), .Y(ori_ori_n846_));
  NA2        o0818(.A(ori_ori_n844_), .B(ori_ori_n629_), .Y(ori_ori_n847_));
  AOI220     o0819(.A0(ori_ori_n712_), .A1(ori_ori_n437_), .B0(ori_ori_n488_), .B1(ori_ori_n190_), .Y(ori_ori_n848_));
  NA3        o0820(.A(ori_ori_n848_), .B(ori_ori_n847_), .C(ori_ori_n644_), .Y(ori_ori_n849_));
  NO4        o0821(.A(ori_ori_n849_), .B(ori_ori_n846_), .C(ori_ori_n216_), .D(ori_ori_n839_), .Y(ori_ori_n850_));
  NA2        o0822(.A(ori_ori_n620_), .B(ori_ori_n565_), .Y(ori_ori_n851_));
  NA4        o0823(.A(ori_ori_n851_), .B(ori_ori_n850_), .C(ori_ori_n836_), .D(ori_ori_n819_), .Y(ori01));
  NO2        o0824(.A(ori_ori_n355_), .B(ori_ori_n210_), .Y(ori_ori_n853_));
  NA2        o0825(.A(ori_ori_n288_), .B(i), .Y(ori_ori_n854_));
  NA3        o0826(.A(ori_ori_n854_), .B(ori_ori_n853_), .C(ori_ori_n762_), .Y(ori_ori_n855_));
  NA2        o0827(.A(ori_ori_n448_), .B(ori_ori_n74_), .Y(ori_ori_n856_));
  NA2        o0828(.A(ori_ori_n418_), .B(ori_ori_n206_), .Y(ori_ori_n857_));
  NA2        o0829(.A(ori_ori_n716_), .B(ori_ori_n857_), .Y(ori_ori_n858_));
  NA3        o0830(.A(ori_ori_n858_), .B(ori_ori_n856_), .C(ori_ori_n235_), .Y(ori_ori_n859_));
  NA2        o0831(.A(ori_ori_n533_), .B(ori_ori_n81_), .Y(ori_ori_n860_));
  INV        o0832(.A(ori_ori_n94_), .Y(ori_ori_n861_));
  OA220      o0833(.A0(ori_ori_n861_), .A1(ori_ori_n445_), .B0(ori_ori_n498_), .B1(ori_ori_n265_), .Y(ori_ori_n862_));
  NAi41      o0834(.An(ori_ori_n130_), .B(ori_ori_n862_), .C(ori_ori_n840_), .D(ori_ori_n665_), .Y(ori_ori_n863_));
  NO3        o0835(.A(ori_ori_n581_), .B(ori_ori_n506_), .C(ori_ori_n380_), .Y(ori_ori_n864_));
  NA3        o0836(.A(ori_ori_n533_), .B(ori_ori_n81_), .C(ori_ori_n169_), .Y(ori_ori_n865_));
  OR2        o0837(.A(ori_ori_n865_), .B(ori_ori_n503_), .Y(ori_ori_n866_));
  NA2        o0838(.A(ori_ori_n866_), .B(ori_ori_n864_), .Y(ori_ori_n867_));
  NO4        o0839(.A(ori_ori_n867_), .B(ori_ori_n863_), .C(ori_ori_n859_), .D(ori_ori_n855_), .Y(ori_ori_n868_));
  INV        o0840(.A(ori_ori_n824_), .Y(ori_ori_n869_));
  NA2        o0841(.A(ori_ori_n869_), .B(ori_ori_n397_), .Y(ori_ori_n870_));
  NA2        o0842(.A(ori_ori_n257_), .B(m), .Y(ori_ori_n871_));
  OR2        o0843(.A(ori_ori_n871_), .B(ori_ori_n234_), .Y(ori_ori_n872_));
  NA2        o0844(.A(ori_ori_n872_), .B(ori_ori_n870_), .Y(ori_ori_n873_));
  NA2        o0845(.A(ori_ori_n451_), .B(ori_ori_n94_), .Y(ori_ori_n874_));
  INV        o0846(.A(ori_ori_n874_), .Y(ori_ori_n875_));
  NO3        o0847(.A(ori_ori_n582_), .B(ori_ori_n875_), .C(ori_ori_n873_), .Y(ori_ori_n876_));
  NA3        o0848(.A(ori_ori_n454_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n877_));
  NO2        o0849(.A(ori_ori_n877_), .B(ori_ori_n163_), .Y(ori_ori_n878_));
  AOI210     o0850(.A0(ori_ori_n376_), .A1(ori_ori_n52_), .B0(ori_ori_n878_), .Y(ori_ori_n879_));
  OR2        o0851(.A(ori_ori_n860_), .B(ori_ori_n455_), .Y(ori_ori_n880_));
  NO2        o0852(.A(ori_ori_n865_), .B(ori_ori_n731_), .Y(ori_ori_n881_));
  NO2        o0853(.A(ori_ori_n165_), .B(ori_ori_n90_), .Y(ori_ori_n882_));
  NO2        o0854(.A(ori_ori_n882_), .B(ori_ori_n881_), .Y(ori_ori_n883_));
  NA4        o0855(.A(ori_ori_n883_), .B(ori_ori_n880_), .C(ori_ori_n879_), .D(ori_ori_n564_), .Y(ori_ori_n884_));
  NO2        o0856(.A(ori_ori_n722_), .B(ori_ori_n183_), .Y(ori_ori_n885_));
  NO2        o0857(.A(ori_ori_n723_), .B(ori_ori_n420_), .Y(ori_ori_n886_));
  OAI210     o0858(.A0(ori_ori_n886_), .A1(ori_ori_n885_), .B0(ori_ori_n243_), .Y(ori_ori_n887_));
  NA2        o0859(.A(ori_ori_n432_), .B(ori_ori_n430_), .Y(ori_ori_n888_));
  NO3        o0860(.A(ori_ori_n65_), .B(ori_ori_n220_), .C(ori_ori_n39_), .Y(ori_ori_n889_));
  NA2        o0861(.A(ori_ori_n889_), .B(ori_ori_n417_), .Y(ori_ori_n890_));
  NA2        o0862(.A(ori_ori_n890_), .B(ori_ori_n888_), .Y(ori_ori_n891_));
  OR2        o0863(.A(ori_ori_n824_), .B(ori_ori_n820_), .Y(ori_ori_n892_));
  NO2        o0864(.A(ori_ori_n265_), .B(ori_ori_n58_), .Y(ori_ori_n893_));
  INV        o0865(.A(ori_ori_n893_), .Y(ori_ori_n894_));
  NA2        o0866(.A(ori_ori_n889_), .B(ori_ori_n603_), .Y(ori_ori_n895_));
  NA4        o0867(.A(ori_ori_n895_), .B(ori_ori_n894_), .C(ori_ori_n892_), .D(ori_ori_n280_), .Y(ori_ori_n896_));
  NOi41      o0868(.An(ori_ori_n887_), .B(ori_ori_n896_), .C(ori_ori_n891_), .D(ori_ori_n884_), .Y(ori_ori_n897_));
  INV        o0869(.A(ori_ori_n105_), .Y(ori_ori_n898_));
  NO3        o0870(.A(ori_ori_n780_), .B(ori_ori_n138_), .C(ori_ori_n71_), .Y(ori_ori_n899_));
  AOI220     o0871(.A0(ori_ori_n899_), .A1(ori_ori_n898_), .B0(ori_ori_n889_), .B1(ori_ori_n726_), .Y(ori_ori_n900_));
  INV        o0872(.A(ori_ori_n900_), .Y(ori_ori_n901_));
  NO2        o0873(.A(ori_ori_n462_), .B(ori_ori_n461_), .Y(ori_ori_n902_));
  NO4        o0874(.A(ori_ori_n780_), .B(ori_ori_n902_), .C(ori_ori_n136_), .D(ori_ori_n71_), .Y(ori_ori_n903_));
  NO3        o0875(.A(ori_ori_n903_), .B(ori_ori_n901_), .C(ori_ori_n481_), .Y(ori_ori_n904_));
  NA4        o0876(.A(ori_ori_n904_), .B(ori_ori_n897_), .C(ori_ori_n876_), .D(ori_ori_n868_), .Y(ori06));
  NO2        o0877(.A(ori_ori_n179_), .B(ori_ori_n84_), .Y(ori_ori_n906_));
  OAI210     o0878(.A0(ori_ori_n906_), .A1(ori_ori_n899_), .B0(ori_ori_n276_), .Y(ori_ori_n907_));
  INV        o0879(.A(ori_ori_n602_), .Y(ori_ori_n908_));
  NA2        o0880(.A(ori_ori_n907_), .B(ori_ori_n887_), .Y(ori_ori_n909_));
  NO3        o0881(.A(ori_ori_n909_), .B(ori_ori_n891_), .C(ori_ori_n201_), .Y(ori_ori_n910_));
  NO2        o0882(.A(ori_ori_n220_), .B(ori_ori_n39_), .Y(ori_ori_n911_));
  AOI210     o0883(.A0(ori_ori_n911_), .A1(ori_ori_n727_), .B0(ori_ori_n885_), .Y(ori_ori_n912_));
  NA2        o0884(.A(ori_ori_n911_), .B(ori_ori_n421_), .Y(ori_ori_n913_));
  AOI210     o0885(.A0(ori_ori_n913_), .A1(ori_ori_n912_), .B0(ori_ori_n240_), .Y(ori_ori_n914_));
  NO2        o0886(.A(ori_ori_n382_), .B(ori_ori_n133_), .Y(ori_ori_n915_));
  NO2        o0887(.A(ori_ori_n457_), .B(ori_ori_n792_), .Y(ori_ori_n916_));
  NO2        o0888(.A(ori_ori_n916_), .B(ori_ori_n915_), .Y(ori_ori_n917_));
  INV        o0889(.A(ori_ori_n917_), .Y(ori_ori_n918_));
  AN2        o0890(.A(ori_ori_n712_), .B(ori_ori_n484_), .Y(ori_ori_n919_));
  NO3        o0891(.A(ori_ori_n919_), .B(ori_ori_n918_), .C(ori_ori_n914_), .Y(ori_ori_n920_));
  NO2        o0892(.A(ori_ori_n379_), .B(ori_ori_n382_), .Y(ori_ori_n921_));
  INV        o0893(.A(k), .Y(ori_ori_n922_));
  NO3        o0894(.A(ori_ori_n922_), .B(ori_ori_n453_), .C(j), .Y(ori_ori_n923_));
  NOi21      o0895(.An(ori_ori_n923_), .B(ori_ori_n503_), .Y(ori_ori_n924_));
  NO2        o0896(.A(ori_ori_n924_), .B(ori_ori_n921_), .Y(ori_ori_n925_));
  NA2        o0897(.A(ori_ori_n591_), .B(ori_ori_n590_), .Y(ori_ori_n926_));
  NAi31      o0898(.An(ori_ori_n558_), .B(ori_ori_n926_), .C(ori_ori_n162_), .Y(ori_ori_n927_));
  NA3        o0899(.A(ori_ori_n927_), .B(ori_ori_n925_), .C(ori_ori_n848_), .Y(ori_ori_n928_));
  OR3        o0900(.A(ori_ori_n908_), .B(ori_ori_n580_), .C(ori_ori_n406_), .Y(ori_ori_n929_));
  AOI210     o0901(.A0(ori_ori_n432_), .A1(ori_ori_n330_), .B0(ori_ori_n268_), .Y(ori_ori_n930_));
  NA2        o0902(.A(ori_ori_n923_), .B(ori_ori_n587_), .Y(ori_ori_n931_));
  NA3        o0903(.A(ori_ori_n931_), .B(ori_ori_n930_), .C(ori_ori_n929_), .Y(ori_ori_n932_));
  AN2        o0904(.A(ori_ori_n686_), .B(ori_ori_n685_), .Y(ori_ori_n933_));
  NO3        o0905(.A(ori_ori_n933_), .B(ori_ori_n650_), .C(ori_ori_n372_), .Y(ori_ori_n934_));
  NA2        o0906(.A(ori_ori_n934_), .B(ori_ori_n895_), .Y(ori_ori_n935_));
  NAi21      o0907(.An(j), .B(i), .Y(ori_ori_n936_));
  NO4        o0908(.A(ori_ori_n902_), .B(ori_ori_n936_), .C(ori_ori_n325_), .D(ori_ori_n185_), .Y(ori_ori_n937_));
  NO4        o0909(.A(ori_ori_n937_), .B(ori_ori_n935_), .C(ori_ori_n932_), .D(ori_ori_n928_), .Y(ori_ori_n938_));
  NA4        o0910(.A(ori_ori_n938_), .B(ori_ori_n920_), .C(ori_ori_n910_), .D(ori_ori_n904_), .Y(ori07));
  NAi32      o0911(.An(m), .Bn(b), .C(n), .Y(ori_ori_n940_));
  NO3        o0912(.A(ori_ori_n940_), .B(g), .C(f), .Y(ori_ori_n941_));
  NAi21      o0913(.An(f), .B(c), .Y(ori_ori_n942_));
  NOi31      o0914(.An(n), .B(m), .C(b), .Y(ori_ori_n943_));
  NO3        o0915(.A(ori_ori_n104_), .B(ori_ori_n332_), .C(h), .Y(ori_ori_n944_));
  NOi31      o0916(.An(i), .B(n), .C(h), .Y(ori_ori_n945_));
  NO2        o0917(.A(ori_ori_n773_), .B(ori_ori_n325_), .Y(ori_ori_n946_));
  NO2        o0918(.A(ori_ori_n775_), .B(ori_ori_n223_), .Y(ori_ori_n947_));
  NO2        o0919(.A(ori_ori_n946_), .B(ori_ori_n941_), .Y(ori_ori_n948_));
  NA3        o0920(.A(ori_ori_n521_), .B(ori_ori_n509_), .C(ori_ori_n91_), .Y(ori_ori_n949_));
  NO2        o0921(.A(l), .B(k), .Y(ori_ori_n950_));
  NO3        o0922(.A(ori_ori_n325_), .B(d), .C(c), .Y(ori_ori_n951_));
  NO2        o0923(.A(g), .B(c), .Y(ori_ori_n952_));
  NO2        o0924(.A(ori_ori_n335_), .B(a), .Y(ori_ori_n953_));
  NA2        o0925(.A(ori_ori_n953_), .B(ori_ori_n92_), .Y(ori_ori_n954_));
  NOi31      o0926(.An(m), .B(n), .C(b), .Y(ori_ori_n955_));
  NOi31      o0927(.An(f), .B(d), .C(c), .Y(ori_ori_n956_));
  NA2        o0928(.A(ori_ori_n956_), .B(ori_ori_n955_), .Y(ori_ori_n957_));
  NA2        o0929(.A(ori_ori_n778_), .B(ori_ori_n348_), .Y(ori_ori_n958_));
  NO2        o0930(.A(ori_ori_n958_), .B(ori_ori_n325_), .Y(ori_ori_n959_));
  NO3        o0931(.A(ori_ori_n37_), .B(i), .C(h), .Y(ori_ori_n960_));
  NO2        o0932(.A(ori_ori_n774_), .B(ori_ori_n959_), .Y(ori_ori_n961_));
  AN3        o0933(.A(ori_ori_n961_), .B(ori_ori_n957_), .C(ori_ori_n954_), .Y(ori_ori_n962_));
  NA2        o0934(.A(ori_ori_n943_), .B(ori_ori_n273_), .Y(ori_ori_n963_));
  INV        o0935(.A(ori_ori_n963_), .Y(ori_ori_n964_));
  INV        o0936(.A(ori_ori_n781_), .Y(ori_ori_n965_));
  NAi21      o0937(.An(ori_ori_n964_), .B(ori_ori_n965_), .Y(ori_ori_n966_));
  NO4        o0938(.A(ori_ori_n104_), .B(g), .C(f), .D(e), .Y(ori_ori_n967_));
  NA2        o0939(.A(ori_ori_n945_), .B(ori_ori_n950_), .Y(ori_ori_n968_));
  INV        o0940(.A(ori_ori_n968_), .Y(ori_ori_n969_));
  NA2        o0941(.A(ori_ori_n791_), .B(ori_ori_n301_), .Y(ori_ori_n970_));
  NO2        o0942(.A(ori_ori_n970_), .B(ori_ori_n318_), .Y(ori_ori_n971_));
  AO210      o0943(.A0(ori_ori_n971_), .A1(ori_ori_n93_), .B0(ori_ori_n969_), .Y(ori_ori_n972_));
  NO2        o0944(.A(ori_ori_n972_), .B(ori_ori_n966_), .Y(ori_ori_n973_));
  NA4        o0945(.A(ori_ori_n973_), .B(ori_ori_n962_), .C(ori_ori_n949_), .D(ori_ori_n948_), .Y(ori_ori_n974_));
  NO2        o0946(.A(ori_ori_n285_), .B(j), .Y(ori_ori_n975_));
  NA2        o0947(.A(ori_ori_n960_), .B(ori_ori_n791_), .Y(ori_ori_n976_));
  NA2        o0948(.A(ori_ori_n777_), .B(e), .Y(ori_ori_n977_));
  NA2        o0949(.A(ori_ori_n977_), .B(ori_ori_n976_), .Y(ori_ori_n978_));
  NA2        o0950(.A(ori_ori_n975_), .B(ori_ori_n127_), .Y(ori_ori_n979_));
  INV        o0951(.A(ori_ori_n979_), .Y(ori_ori_n980_));
  NO2        o0952(.A(ori_ori_n980_), .B(ori_ori_n978_), .Y(ori_ori_n981_));
  INV        o0953(.A(ori_ori_n43_), .Y(ori_ori_n982_));
  NA2        o0954(.A(ori_ori_n982_), .B(ori_ori_n826_), .Y(ori_ori_n983_));
  INV        o0955(.A(ori_ori_n983_), .Y(ori_ori_n984_));
  NO2        o0956(.A(ori_ori_n179_), .B(ori_ori_n138_), .Y(ori_ori_n985_));
  NO2        o0957(.A(ori_ori_n985_), .B(ori_ori_n984_), .Y(ori_ori_n986_));
  NA2        o0958(.A(c), .B(f), .Y(ori_ori_n987_));
  NO2        o0959(.A(ori_ori_n1027_), .B(ori_ori_n987_), .Y(ori_ori_n988_));
  NO2        o0960(.A(ori_ori_n936_), .B(ori_ori_n136_), .Y(ori_ori_n989_));
  NOi21      o0961(.An(d), .B(f), .Y(ori_ori_n990_));
  NA2        o0962(.A(h), .B(ori_ori_n989_), .Y(ori_ori_n991_));
  NA2        o0963(.A(h), .B(ori_ori_n407_), .Y(ori_ori_n992_));
  NA2        o0964(.A(ori_ori_n992_), .B(ori_ori_n991_), .Y(ori_ori_n993_));
  NO2        o0965(.A(ori_ori_n993_), .B(ori_ori_n988_), .Y(ori_ori_n994_));
  NA3        o0966(.A(ori_ori_n994_), .B(ori_ori_n986_), .C(ori_ori_n981_), .Y(ori_ori_n995_));
  NA2        o0967(.A(h), .B(ori_ori_n947_), .Y(ori_ori_n996_));
  OAI210     o0968(.A0(ori_ori_n967_), .A1(ori_ori_n943_), .B0(ori_ori_n654_), .Y(ori_ori_n997_));
  NA2        o0969(.A(ori_ori_n997_), .B(ori_ori_n996_), .Y(ori_ori_n998_));
  NA2        o0970(.A(ori_ori_n952_), .B(ori_ori_n990_), .Y(ori_ori_n999_));
  NO2        o0971(.A(ori_ori_n999_), .B(m), .Y(ori_ori_n1000_));
  NO2        o0972(.A(ori_ori_n120_), .B(ori_ori_n143_), .Y(ori_ori_n1001_));
  OAI210     o0973(.A0(ori_ori_n1001_), .A1(ori_ori_n89_), .B0(ori_ori_n955_), .Y(ori_ori_n1002_));
  INV        o0974(.A(ori_ori_n1002_), .Y(ori_ori_n1003_));
  NO3        o0975(.A(ori_ori_n1003_), .B(ori_ori_n1000_), .C(ori_ori_n998_), .Y(ori_ori_n1004_));
  NO2        o0976(.A(ori_ori_n942_), .B(e), .Y(ori_ori_n1005_));
  NA2        o0977(.A(ori_ori_n1005_), .B(ori_ori_n299_), .Y(ori_ori_n1006_));
  NA2        o0978(.A(ori_ori_n793_), .B(ori_ori_n477_), .Y(ori_ori_n1007_));
  BUFFER     o0979(.A(ori_ori_n104_), .Y(ori_ori_n1008_));
  OAI210     o0980(.A0(ori_ori_n1008_), .A1(ori_ori_n1006_), .B0(ori_ori_n1007_), .Y(ori_ori_n1009_));
  INV        o0981(.A(ori_ori_n1009_), .Y(ori_ori_n1010_));
  OR2        o0982(.A(h), .B(ori_ori_n405_), .Y(ori_ori_n1011_));
  NO2        o0983(.A(ori_ori_n1011_), .B(ori_ori_n136_), .Y(ori_ori_n1012_));
  NA2        o0984(.A(ori_ori_n782_), .B(ori_ori_n177_), .Y(ori_ori_n1013_));
  NO2        o0985(.A(ori_ori_n43_), .B(l), .Y(ori_ori_n1014_));
  INV        o0986(.A(ori_ori_n357_), .Y(ori_ori_n1015_));
  NA2        o0987(.A(ori_ori_n1015_), .B(ori_ori_n1014_), .Y(ori_ori_n1016_));
  NA2        o0988(.A(ori_ori_n1016_), .B(ori_ori_n1013_), .Y(ori_ori_n1017_));
  NO3        o0989(.A(ori_ori_n1017_), .B(ori_ori_n1012_), .C(ori_ori_n951_), .Y(ori_ori_n1018_));
  NA3        o0990(.A(ori_ori_n1018_), .B(ori_ori_n1010_), .C(ori_ori_n1004_), .Y(ori_ori_n1019_));
  NA3        o0991(.A(ori_ori_n715_), .B(ori_ori_n107_), .C(ori_ori_n40_), .Y(ori_ori_n1020_));
  NO2        o0992(.A(ori_ori_n970_), .B(d), .Y(ori_ori_n1021_));
  INV        o0993(.A(ori_ori_n1021_), .Y(ori_ori_n1022_));
  NA3        o0994(.A(ori_ori_n1022_), .B(ori_ori_n1028_), .C(ori_ori_n1020_), .Y(ori_ori_n1023_));
  OR4        o0995(.A(ori_ori_n1023_), .B(ori_ori_n1019_), .C(ori_ori_n995_), .D(ori_ori_n974_), .Y(ori04));
  INV        o0996(.A(ori_ori_n92_), .Y(ori_ori_n1027_));
  INV        o0997(.A(ori_ori_n944_), .Y(ori_ori_n1028_));
  INV        o0998(.A(j), .Y(ori_ori_n1029_));
  INV        o0999(.A(ori_ori_n225_), .Y(ori_ori_n1030_));
  INV        o1000(.A(ori_ori_n77_), .Y(ori_ori_n1031_));
  INV        o1001(.A(m), .Y(ori_ori_n1032_));
  INV        o1002(.A(g), .Y(ori_ori_n1033_));
  ZERO       o1003(.Y(ori02));
  ZERO       o1004(.Y(ori03));
  ZERO       o1005(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  NO3        m0023(.A(mai_mai_n48_), .B(mai_mai_n43_), .C(mai_mai_n39_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n32_), .Y(mai_mai_n53_));
  INV        m0025(.A(c), .Y(mai_mai_n54_));
  NA2        m0026(.A(e), .B(b), .Y(mai_mai_n55_));
  NO2        m0027(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  INV        m0028(.A(d), .Y(mai_mai_n57_));
  NAi21      m0029(.An(i), .B(h), .Y(mai_mai_n58_));
  NAi31      m0030(.An(i), .B(l), .C(j), .Y(mai_mai_n59_));
  NAi41      m0031(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n60_));
  NA2        m0032(.A(g), .B(f), .Y(mai_mai_n61_));
  NO2        m0033(.A(mai_mai_n61_), .B(mai_mai_n60_), .Y(mai_mai_n62_));
  NAi21      m0034(.An(i), .B(j), .Y(mai_mai_n63_));
  NAi32      m0035(.An(n), .Bn(k), .C(m), .Y(mai_mai_n64_));
  NO2        m0036(.A(mai_mai_n64_), .B(mai_mai_n63_), .Y(mai_mai_n65_));
  NAi31      m0037(.An(l), .B(m), .C(k), .Y(mai_mai_n66_));
  NAi41      m0038(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n67_));
  NA2        m0039(.A(mai_mai_n65_), .B(mai_mai_n62_), .Y(mai_mai_n68_));
  INV        m0040(.A(m), .Y(mai_mai_n69_));
  NOi21      m0041(.An(k), .B(l), .Y(mai_mai_n70_));
  NA2        m0042(.A(mai_mai_n70_), .B(mai_mai_n69_), .Y(mai_mai_n71_));
  AN4        m0043(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n72_));
  NOi31      m0044(.An(h), .B(g), .C(f), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  NAi32      m0046(.An(m), .Bn(k), .C(j), .Y(mai_mai_n75_));
  NOi32      m0047(.An(h), .Bn(g), .C(f), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n72_), .Y(mai_mai_n77_));
  OA220      m0049(.A0(mai_mai_n77_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .B1(mai_mai_n71_), .Y(mai_mai_n78_));
  NA2        m0050(.A(mai_mai_n78_), .B(mai_mai_n68_), .Y(mai_mai_n79_));
  INV        m0051(.A(n), .Y(mai_mai_n80_));
  NOi32      m0052(.An(e), .Bn(b), .C(d), .Y(mai_mai_n81_));
  NA2        m0053(.A(mai_mai_n81_), .B(mai_mai_n80_), .Y(mai_mai_n82_));
  INV        m0054(.A(j), .Y(mai_mai_n83_));
  AN3        m0055(.A(m), .B(k), .C(i), .Y(mai_mai_n84_));
  NA3        m0056(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(g), .Y(mai_mai_n85_));
  NAi32      m0057(.An(g), .Bn(f), .C(h), .Y(mai_mai_n86_));
  NAi31      m0058(.An(j), .B(m), .C(l), .Y(mai_mai_n87_));
  NA2        m0059(.A(m), .B(l), .Y(mai_mai_n88_));
  NAi31      m0060(.An(k), .B(j), .C(g), .Y(mai_mai_n89_));
  NO3        m0061(.A(mai_mai_n89_), .B(mai_mai_n88_), .C(f), .Y(mai_mai_n90_));
  AN2        m0062(.A(j), .B(g), .Y(mai_mai_n91_));
  NOi32      m0063(.An(m), .Bn(l), .C(i), .Y(mai_mai_n92_));
  NOi21      m0064(.An(g), .B(i), .Y(mai_mai_n93_));
  NOi32      m0065(.An(m), .Bn(j), .C(k), .Y(mai_mai_n94_));
  AOI220     m0066(.A0(mai_mai_n94_), .A1(mai_mai_n93_), .B0(mai_mai_n92_), .B1(mai_mai_n91_), .Y(mai_mai_n95_));
  NAi41      m0067(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n96_));
  AN2        m0068(.A(e), .B(b), .Y(mai_mai_n97_));
  NOi31      m0069(.An(c), .B(h), .C(f), .Y(mai_mai_n98_));
  NA2        m0070(.A(mai_mai_n98_), .B(mai_mai_n97_), .Y(mai_mai_n99_));
  NO2        m0071(.A(mai_mai_n99_), .B(mai_mai_n96_), .Y(mai_mai_n100_));
  NOi21      m0072(.An(i), .B(h), .Y(mai_mai_n101_));
  NA3        m0073(.A(mai_mai_n101_), .B(g), .C(mai_mai_n36_), .Y(mai_mai_n102_));
  INV        m0074(.A(a), .Y(mai_mai_n103_));
  NA2        m0075(.A(mai_mai_n97_), .B(mai_mai_n103_), .Y(mai_mai_n104_));
  INV        m0076(.A(l), .Y(mai_mai_n105_));
  NOi21      m0077(.An(m), .B(n), .Y(mai_mai_n106_));
  AN2        m0078(.A(k), .B(h), .Y(mai_mai_n107_));
  NO2        m0079(.A(mai_mai_n102_), .B(mai_mai_n82_), .Y(mai_mai_n108_));
  INV        m0080(.A(b), .Y(mai_mai_n109_));
  NA2        m0081(.A(l), .B(j), .Y(mai_mai_n110_));
  AN2        m0082(.A(k), .B(i), .Y(mai_mai_n111_));
  NA2        m0083(.A(mai_mai_n111_), .B(mai_mai_n110_), .Y(mai_mai_n112_));
  NA2        m0084(.A(g), .B(e), .Y(mai_mai_n113_));
  NOi32      m0085(.An(c), .Bn(a), .C(d), .Y(mai_mai_n114_));
  NA2        m0086(.A(mai_mai_n114_), .B(mai_mai_n106_), .Y(mai_mai_n115_));
  NO4        m0087(.A(mai_mai_n115_), .B(mai_mai_n113_), .C(mai_mai_n112_), .D(mai_mai_n109_), .Y(mai_mai_n116_));
  NO3        m0088(.A(mai_mai_n116_), .B(mai_mai_n108_), .C(mai_mai_n100_), .Y(mai_mai_n117_));
  OAI210     m0089(.A0(mai_mai_n95_), .A1(mai_mai_n82_), .B0(mai_mai_n117_), .Y(mai_mai_n118_));
  NOi31      m0090(.An(k), .B(m), .C(j), .Y(mai_mai_n119_));
  NOi31      m0091(.An(k), .B(m), .C(i), .Y(mai_mai_n120_));
  NOi32      m0092(.An(f), .Bn(b), .C(e), .Y(mai_mai_n121_));
  NAi21      m0093(.An(g), .B(h), .Y(mai_mai_n122_));
  NAi21      m0094(.An(m), .B(n), .Y(mai_mai_n123_));
  NAi21      m0095(.An(j), .B(k), .Y(mai_mai_n124_));
  NO3        m0096(.A(mai_mai_n124_), .B(mai_mai_n123_), .C(mai_mai_n122_), .Y(mai_mai_n125_));
  NAi41      m0097(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n126_));
  NAi31      m0098(.An(j), .B(k), .C(h), .Y(mai_mai_n127_));
  NO3        m0099(.A(mai_mai_n127_), .B(mai_mai_n126_), .C(mai_mai_n123_), .Y(mai_mai_n128_));
  AOI210     m0100(.A0(mai_mai_n125_), .A1(mai_mai_n121_), .B0(mai_mai_n128_), .Y(mai_mai_n129_));
  NO2        m0101(.A(k), .B(j), .Y(mai_mai_n130_));
  AN2        m0102(.A(k), .B(j), .Y(mai_mai_n131_));
  NAi21      m0103(.An(c), .B(b), .Y(mai_mai_n132_));
  NA2        m0104(.A(f), .B(d), .Y(mai_mai_n133_));
  NAi31      m0105(.An(f), .B(e), .C(b), .Y(mai_mai_n134_));
  NA2        m0106(.A(d), .B(b), .Y(mai_mai_n135_));
  NO2        m0107(.A(e), .B(mai_mai_n135_), .Y(mai_mai_n136_));
  NA2        m0108(.A(b), .B(a), .Y(mai_mai_n137_));
  NAi21      m0109(.An(e), .B(g), .Y(mai_mai_n138_));
  NAi21      m0110(.An(c), .B(d), .Y(mai_mai_n139_));
  NAi31      m0111(.An(l), .B(k), .C(h), .Y(mai_mai_n140_));
  INV        m0112(.A(mai_mai_n129_), .Y(mai_mai_n141_));
  NAi31      m0113(.An(e), .B(f), .C(b), .Y(mai_mai_n142_));
  NOi21      m0114(.An(h), .B(i), .Y(mai_mai_n143_));
  NOi21      m0115(.An(k), .B(m), .Y(mai_mai_n144_));
  NA3        m0116(.A(mai_mai_n144_), .B(mai_mai_n143_), .C(n), .Y(mai_mai_n145_));
  NOi21      m0117(.An(h), .B(g), .Y(mai_mai_n146_));
  NO2        m0118(.A(mai_mai_n133_), .B(mai_mai_n132_), .Y(mai_mai_n147_));
  NA2        m0119(.A(mai_mai_n147_), .B(mai_mai_n146_), .Y(mai_mai_n148_));
  NAi31      m0120(.An(l), .B(j), .C(h), .Y(mai_mai_n149_));
  NO2        m0121(.A(mai_mai_n149_), .B(mai_mai_n49_), .Y(mai_mai_n150_));
  NA2        m0122(.A(mai_mai_n150_), .B(mai_mai_n62_), .Y(mai_mai_n151_));
  NOi32      m0123(.An(n), .Bn(k), .C(m), .Y(mai_mai_n152_));
  NA2        m0124(.A(l), .B(i), .Y(mai_mai_n153_));
  NA2        m0125(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  OAI210     m0126(.A0(mai_mai_n154_), .A1(mai_mai_n148_), .B0(mai_mai_n151_), .Y(mai_mai_n155_));
  NA2        m0127(.A(j), .B(h), .Y(mai_mai_n156_));
  OR3        m0128(.A(n), .B(m), .C(k), .Y(mai_mai_n157_));
  NAi32      m0129(.An(m), .Bn(k), .C(n), .Y(mai_mai_n158_));
  NO2        m0130(.A(n), .B(m), .Y(mai_mai_n159_));
  NA2        m0131(.A(mai_mai_n159_), .B(mai_mai_n50_), .Y(mai_mai_n160_));
  NAi21      m0132(.An(f), .B(e), .Y(mai_mai_n161_));
  NA2        m0133(.A(d), .B(c), .Y(mai_mai_n162_));
  NO2        m0134(.A(mai_mai_n162_), .B(mai_mai_n161_), .Y(mai_mai_n163_));
  NOi21      m0135(.An(mai_mai_n163_), .B(mai_mai_n160_), .Y(mai_mai_n164_));
  NAi21      m0136(.An(d), .B(c), .Y(mai_mai_n165_));
  NAi31      m0137(.An(m), .B(n), .C(b), .Y(mai_mai_n166_));
  NA2        m0138(.A(k), .B(i), .Y(mai_mai_n167_));
  NAi21      m0139(.An(h), .B(f), .Y(mai_mai_n168_));
  NO2        m0140(.A(mai_mai_n168_), .B(mai_mai_n167_), .Y(mai_mai_n169_));
  NO2        m0141(.A(mai_mai_n166_), .B(mai_mai_n139_), .Y(mai_mai_n170_));
  NA2        m0142(.A(mai_mai_n170_), .B(mai_mai_n169_), .Y(mai_mai_n171_));
  NOi32      m0143(.An(f), .Bn(c), .C(d), .Y(mai_mai_n172_));
  NOi32      m0144(.An(f), .Bn(c), .C(e), .Y(mai_mai_n173_));
  NO2        m0145(.A(mai_mai_n173_), .B(mai_mai_n172_), .Y(mai_mai_n174_));
  NO3        m0146(.A(n), .B(m), .C(j), .Y(mai_mai_n175_));
  NA2        m0147(.A(mai_mai_n175_), .B(mai_mai_n107_), .Y(mai_mai_n176_));
  AO210      m0148(.A0(mai_mai_n176_), .A1(mai_mai_n160_), .B0(mai_mai_n174_), .Y(mai_mai_n177_));
  NAi31      m0149(.An(mai_mai_n164_), .B(mai_mai_n177_), .C(mai_mai_n171_), .Y(mai_mai_n178_));
  OR3        m0150(.A(mai_mai_n178_), .B(mai_mai_n155_), .C(mai_mai_n141_), .Y(mai_mai_n179_));
  NO4        m0151(.A(mai_mai_n179_), .B(mai_mai_n118_), .C(mai_mai_n79_), .D(mai_mai_n53_), .Y(mai_mai_n180_));
  NA3        m0152(.A(m), .B(mai_mai_n105_), .C(j), .Y(mai_mai_n181_));
  NAi31      m0153(.An(n), .B(h), .C(g), .Y(mai_mai_n182_));
  NO2        m0154(.A(mai_mai_n182_), .B(mai_mai_n181_), .Y(mai_mai_n183_));
  NOi32      m0155(.An(m), .Bn(k), .C(l), .Y(mai_mai_n184_));
  NA3        m0156(.A(mai_mai_n184_), .B(mai_mai_n83_), .C(g), .Y(mai_mai_n185_));
  NO2        m0157(.A(mai_mai_n185_), .B(n), .Y(mai_mai_n186_));
  NOi21      m0158(.An(k), .B(j), .Y(mai_mai_n187_));
  NA4        m0159(.A(mai_mai_n187_), .B(mai_mai_n106_), .C(i), .D(g), .Y(mai_mai_n188_));
  AN2        m0160(.A(i), .B(g), .Y(mai_mai_n189_));
  NA3        m0161(.A(mai_mai_n70_), .B(mai_mai_n189_), .C(mai_mai_n106_), .Y(mai_mai_n190_));
  NA2        m0162(.A(mai_mai_n190_), .B(mai_mai_n188_), .Y(mai_mai_n191_));
  INV        m0163(.A(mai_mai_n191_), .Y(mai_mai_n192_));
  NAi41      m0164(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n193_));
  INV        m0165(.A(mai_mai_n193_), .Y(mai_mai_n194_));
  INV        m0166(.A(f), .Y(mai_mai_n195_));
  INV        m0167(.A(g), .Y(mai_mai_n196_));
  NOi31      m0168(.An(i), .B(j), .C(h), .Y(mai_mai_n197_));
  NOi21      m0169(.An(l), .B(m), .Y(mai_mai_n198_));
  NA2        m0170(.A(mai_mai_n198_), .B(mai_mai_n197_), .Y(mai_mai_n199_));
  NO3        m0171(.A(mai_mai_n199_), .B(mai_mai_n196_), .C(mai_mai_n195_), .Y(mai_mai_n200_));
  NA2        m0172(.A(mai_mai_n200_), .B(mai_mai_n194_), .Y(mai_mai_n201_));
  OAI210     m0173(.A0(mai_mai_n192_), .A1(mai_mai_n32_), .B0(mai_mai_n201_), .Y(mai_mai_n202_));
  NOi21      m0174(.An(n), .B(m), .Y(mai_mai_n203_));
  NOi32      m0175(.An(l), .Bn(i), .C(j), .Y(mai_mai_n204_));
  NA2        m0176(.A(mai_mai_n204_), .B(mai_mai_n203_), .Y(mai_mai_n205_));
  OA220      m0177(.A0(mai_mai_n205_), .A1(mai_mai_n99_), .B0(mai_mai_n75_), .B1(mai_mai_n74_), .Y(mai_mai_n206_));
  NAi21      m0178(.An(j), .B(h), .Y(mai_mai_n207_));
  XN2        m0179(.A(i), .B(h), .Y(mai_mai_n208_));
  NA2        m0180(.A(mai_mai_n208_), .B(mai_mai_n207_), .Y(mai_mai_n209_));
  NOi31      m0181(.An(k), .B(n), .C(m), .Y(mai_mai_n210_));
  NOi31      m0182(.An(mai_mai_n210_), .B(mai_mai_n162_), .C(mai_mai_n161_), .Y(mai_mai_n211_));
  NA2        m0183(.A(mai_mai_n211_), .B(mai_mai_n209_), .Y(mai_mai_n212_));
  NAi31      m0184(.An(f), .B(e), .C(c), .Y(mai_mai_n213_));
  NO4        m0185(.A(mai_mai_n213_), .B(mai_mai_n157_), .C(mai_mai_n156_), .D(mai_mai_n57_), .Y(mai_mai_n214_));
  NA4        m0186(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n215_));
  NAi32      m0187(.An(m), .Bn(i), .C(k), .Y(mai_mai_n216_));
  NO3        m0188(.A(mai_mai_n216_), .B(mai_mai_n86_), .C(mai_mai_n215_), .Y(mai_mai_n217_));
  INV        m0189(.A(k), .Y(mai_mai_n218_));
  NO2        m0190(.A(mai_mai_n217_), .B(mai_mai_n214_), .Y(mai_mai_n219_));
  NAi21      m0191(.An(n), .B(a), .Y(mai_mai_n220_));
  NO2        m0192(.A(mai_mai_n220_), .B(mai_mai_n135_), .Y(mai_mai_n221_));
  NAi41      m0193(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n222_));
  NO2        m0194(.A(mai_mai_n222_), .B(e), .Y(mai_mai_n223_));
  NO3        m0195(.A(e), .B(mai_mai_n89_), .C(mai_mai_n88_), .Y(mai_mai_n224_));
  OAI210     m0196(.A0(mai_mai_n224_), .A1(mai_mai_n223_), .B0(mai_mai_n221_), .Y(mai_mai_n225_));
  AN4        m0197(.A(mai_mai_n225_), .B(mai_mai_n219_), .C(mai_mai_n212_), .D(mai_mai_n206_), .Y(mai_mai_n226_));
  OR2        m0198(.A(h), .B(g), .Y(mai_mai_n227_));
  NO2        m0199(.A(mai_mai_n227_), .B(mai_mai_n96_), .Y(mai_mai_n228_));
  NA2        m0200(.A(mai_mai_n228_), .B(mai_mai_n121_), .Y(mai_mai_n229_));
  NA2        m0201(.A(mai_mai_n144_), .B(mai_mai_n101_), .Y(mai_mai_n230_));
  NO2        m0202(.A(n), .B(a), .Y(mai_mai_n231_));
  NAi31      m0203(.An(mai_mai_n222_), .B(mai_mai_n231_), .C(mai_mai_n97_), .Y(mai_mai_n232_));
  NAi21      m0204(.An(h), .B(i), .Y(mai_mai_n233_));
  NA2        m0205(.A(mai_mai_n159_), .B(k), .Y(mai_mai_n234_));
  NO2        m0206(.A(mai_mai_n234_), .B(mai_mai_n233_), .Y(mai_mai_n235_));
  NA2        m0207(.A(mai_mai_n232_), .B(mai_mai_n229_), .Y(mai_mai_n236_));
  NOi21      m0208(.An(g), .B(e), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n67_), .B(mai_mai_n69_), .Y(mai_mai_n238_));
  NA2        m0210(.A(mai_mai_n238_), .B(mai_mai_n237_), .Y(mai_mai_n239_));
  NOi32      m0211(.An(l), .Bn(j), .C(i), .Y(mai_mai_n240_));
  AOI210     m0212(.A0(mai_mai_n70_), .A1(mai_mai_n83_), .B0(mai_mai_n240_), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n233_), .B(mai_mai_n44_), .Y(mai_mai_n242_));
  NAi21      m0214(.An(f), .B(g), .Y(mai_mai_n243_));
  NO2        m0215(.A(mai_mai_n243_), .B(mai_mai_n60_), .Y(mai_mai_n244_));
  NO2        m0216(.A(mai_mai_n64_), .B(mai_mai_n110_), .Y(mai_mai_n245_));
  AOI220     m0217(.A0(mai_mai_n245_), .A1(mai_mai_n244_), .B0(mai_mai_n242_), .B1(mai_mai_n62_), .Y(mai_mai_n246_));
  OAI210     m0218(.A0(mai_mai_n241_), .A1(mai_mai_n239_), .B0(mai_mai_n246_), .Y(mai_mai_n247_));
  NO3        m0219(.A(mai_mai_n124_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n248_));
  NOi41      m0220(.An(mai_mai_n226_), .B(mai_mai_n247_), .C(mai_mai_n236_), .D(mai_mai_n202_), .Y(mai_mai_n249_));
  NO4        m0221(.A(mai_mai_n183_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n250_));
  NO2        m0222(.A(mai_mai_n250_), .B(mai_mai_n104_), .Y(mai_mai_n251_));
  NA3        m0223(.A(mai_mai_n57_), .B(c), .C(b), .Y(mai_mai_n252_));
  NAi21      m0224(.An(h), .B(g), .Y(mai_mai_n253_));
  OR4        m0225(.A(mai_mai_n253_), .B(mai_mai_n252_), .C(mai_mai_n205_), .D(e), .Y(mai_mai_n254_));
  NO2        m0226(.A(mai_mai_n230_), .B(mai_mai_n243_), .Y(mai_mai_n255_));
  NAi31      m0227(.An(g), .B(k), .C(h), .Y(mai_mai_n256_));
  NO3        m0228(.A(mai_mai_n123_), .B(mai_mai_n256_), .C(l), .Y(mai_mai_n257_));
  NAi31      m0229(.An(e), .B(d), .C(a), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n257_), .B(mai_mai_n121_), .Y(mai_mai_n259_));
  NA2        m0231(.A(mai_mai_n259_), .B(mai_mai_n254_), .Y(mai_mai_n260_));
  NA3        m0232(.A(mai_mai_n144_), .B(mai_mai_n76_), .C(mai_mai_n72_), .Y(mai_mai_n261_));
  NA3        m0233(.A(mai_mai_n144_), .B(mai_mai_n143_), .C(mai_mai_n80_), .Y(mai_mai_n262_));
  BUFFER     m0234(.A(mai_mai_n261_), .Y(mai_mai_n263_));
  NA3        m0235(.A(e), .B(c), .C(b), .Y(mai_mai_n264_));
  NAi32      m0236(.An(k), .Bn(i), .C(j), .Y(mai_mai_n265_));
  NAi31      m0237(.An(h), .B(l), .C(i), .Y(mai_mai_n266_));
  NA3        m0238(.A(mai_mai_n266_), .B(mai_mai_n265_), .C(mai_mai_n149_), .Y(mai_mai_n267_));
  NOi21      m0239(.An(mai_mai_n267_), .B(mai_mai_n49_), .Y(mai_mai_n268_));
  NA2        m0240(.A(mai_mai_n244_), .B(mai_mai_n268_), .Y(mai_mai_n269_));
  NAi21      m0241(.An(l), .B(k), .Y(mai_mai_n270_));
  NO2        m0242(.A(mai_mai_n270_), .B(mai_mai_n49_), .Y(mai_mai_n271_));
  NOi21      m0243(.An(l), .B(j), .Y(mai_mai_n272_));
  NA2        m0244(.A(mai_mai_n146_), .B(mai_mai_n272_), .Y(mai_mai_n273_));
  NAi32      m0245(.An(j), .Bn(h), .C(i), .Y(mai_mai_n274_));
  NAi21      m0246(.An(m), .B(l), .Y(mai_mai_n275_));
  NO3        m0247(.A(mai_mai_n275_), .B(mai_mai_n274_), .C(mai_mai_n80_), .Y(mai_mai_n276_));
  NA2        m0248(.A(h), .B(g), .Y(mai_mai_n277_));
  NA2        m0249(.A(mai_mai_n152_), .B(mai_mai_n45_), .Y(mai_mai_n278_));
  NO2        m0250(.A(mai_mai_n278_), .B(mai_mai_n277_), .Y(mai_mai_n279_));
  OAI210     m0251(.A0(mai_mai_n279_), .A1(mai_mai_n276_), .B0(mai_mai_n147_), .Y(mai_mai_n280_));
  NA3        m0252(.A(mai_mai_n280_), .B(mai_mai_n269_), .C(mai_mai_n263_), .Y(mai_mai_n281_));
  NO2        m0253(.A(mai_mai_n99_), .B(mai_mai_n96_), .Y(mai_mai_n282_));
  NAi32      m0254(.An(n), .Bn(m), .C(l), .Y(mai_mai_n283_));
  NO2        m0255(.A(mai_mai_n283_), .B(mai_mai_n274_), .Y(mai_mai_n284_));
  NA2        m0256(.A(mai_mai_n284_), .B(mai_mai_n163_), .Y(mai_mai_n285_));
  NO2        m0257(.A(mai_mai_n115_), .B(mai_mai_n109_), .Y(mai_mai_n286_));
  NAi31      m0258(.An(k), .B(l), .C(j), .Y(mai_mai_n287_));
  OAI210     m0259(.A0(mai_mai_n270_), .A1(j), .B0(mai_mai_n287_), .Y(mai_mai_n288_));
  NOi21      m0260(.An(mai_mai_n288_), .B(mai_mai_n113_), .Y(mai_mai_n289_));
  NA2        m0261(.A(mai_mai_n289_), .B(mai_mai_n286_), .Y(mai_mai_n290_));
  NA2        m0262(.A(mai_mai_n290_), .B(mai_mai_n285_), .Y(mai_mai_n291_));
  NO4        m0263(.A(mai_mai_n291_), .B(mai_mai_n281_), .C(mai_mai_n260_), .D(mai_mai_n251_), .Y(mai_mai_n292_));
  NA2        m0264(.A(mai_mai_n235_), .B(mai_mai_n173_), .Y(mai_mai_n293_));
  NAi21      m0265(.An(m), .B(k), .Y(mai_mai_n294_));
  NO2        m0266(.A(mai_mai_n208_), .B(mai_mai_n294_), .Y(mai_mai_n295_));
  NAi41      m0267(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n296_));
  NO2        m0268(.A(mai_mai_n296_), .B(mai_mai_n138_), .Y(mai_mai_n297_));
  NA2        m0269(.A(mai_mai_n297_), .B(mai_mai_n295_), .Y(mai_mai_n298_));
  NAi31      m0270(.An(i), .B(l), .C(h), .Y(mai_mai_n299_));
  NO3        m0271(.A(mai_mai_n299_), .B(mai_mai_n138_), .C(mai_mai_n67_), .Y(mai_mai_n300_));
  NA2        m0272(.A(e), .B(c), .Y(mai_mai_n301_));
  NO3        m0273(.A(mai_mai_n301_), .B(n), .C(d), .Y(mai_mai_n302_));
  NOi21      m0274(.An(f), .B(h), .Y(mai_mai_n303_));
  NA2        m0275(.A(mai_mai_n303_), .B(mai_mai_n111_), .Y(mai_mai_n304_));
  NO2        m0276(.A(mai_mai_n304_), .B(mai_mai_n196_), .Y(mai_mai_n305_));
  NAi31      m0277(.An(d), .B(e), .C(b), .Y(mai_mai_n306_));
  NO2        m0278(.A(mai_mai_n123_), .B(mai_mai_n306_), .Y(mai_mai_n307_));
  NA2        m0279(.A(mai_mai_n307_), .B(mai_mai_n305_), .Y(mai_mai_n308_));
  NAi41      m0280(.An(mai_mai_n300_), .B(mai_mai_n308_), .C(mai_mai_n298_), .D(mai_mai_n293_), .Y(mai_mai_n309_));
  NO4        m0281(.A(mai_mai_n296_), .B(mai_mai_n75_), .C(e), .D(mai_mai_n196_), .Y(mai_mai_n310_));
  NA2        m0282(.A(mai_mai_n231_), .B(mai_mai_n97_), .Y(mai_mai_n311_));
  OR2        m0283(.A(mai_mai_n311_), .B(mai_mai_n185_), .Y(mai_mai_n312_));
  NOi31      m0284(.An(l), .B(n), .C(m), .Y(mai_mai_n313_));
  NAi21      m0285(.An(mai_mai_n310_), .B(mai_mai_n312_), .Y(mai_mai_n314_));
  NAi32      m0286(.An(m), .Bn(j), .C(k), .Y(mai_mai_n315_));
  NAi41      m0287(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n193_), .B(mai_mai_n316_), .Y(mai_mai_n317_));
  NOi31      m0289(.An(j), .B(m), .C(k), .Y(mai_mai_n318_));
  NO2        m0290(.A(mai_mai_n119_), .B(mai_mai_n318_), .Y(mai_mai_n319_));
  AN3        m0291(.A(h), .B(g), .C(f), .Y(mai_mai_n320_));
  NAi31      m0292(.An(mai_mai_n319_), .B(mai_mai_n320_), .C(mai_mai_n317_), .Y(mai_mai_n321_));
  NOi32      m0293(.An(m), .Bn(j), .C(l), .Y(mai_mai_n322_));
  NO2        m0294(.A(mai_mai_n322_), .B(mai_mai_n92_), .Y(mai_mai_n323_));
  NO2        m0295(.A(mai_mai_n275_), .B(mai_mai_n274_), .Y(mai_mai_n324_));
  NO2        m0296(.A(mai_mai_n199_), .B(g), .Y(mai_mai_n325_));
  INV        m0297(.A(mai_mai_n216_), .Y(mai_mai_n326_));
  NA3        m0298(.A(mai_mai_n326_), .B(mai_mai_n320_), .C(mai_mai_n194_), .Y(mai_mai_n327_));
  NA2        m0299(.A(mai_mai_n327_), .B(mai_mai_n321_), .Y(mai_mai_n328_));
  NA3        m0300(.A(h), .B(g), .C(f), .Y(mai_mai_n329_));
  NO2        m0301(.A(mai_mai_n329_), .B(mai_mai_n71_), .Y(mai_mai_n330_));
  NA2        m0302(.A(mai_mai_n316_), .B(mai_mai_n193_), .Y(mai_mai_n331_));
  NA2        m0303(.A(mai_mai_n146_), .B(e), .Y(mai_mai_n332_));
  NO2        m0304(.A(mai_mai_n332_), .B(mai_mai_n41_), .Y(mai_mai_n333_));
  AOI220     m0305(.A0(mai_mai_n333_), .A1(mai_mai_n286_), .B0(mai_mai_n331_), .B1(mai_mai_n330_), .Y(mai_mai_n334_));
  NOi32      m0306(.An(e), .Bn(b), .C(a), .Y(mai_mai_n335_));
  AN2        m0307(.A(l), .B(j), .Y(mai_mai_n336_));
  NA3        m0308(.A(mai_mai_n190_), .B(mai_mai_n188_), .C(mai_mai_n35_), .Y(mai_mai_n337_));
  NA2        m0309(.A(mai_mai_n337_), .B(mai_mai_n335_), .Y(mai_mai_n338_));
  NA2        m0310(.A(mai_mai_n189_), .B(k), .Y(mai_mai_n339_));
  NAi41      m0311(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n340_));
  NA2        m0312(.A(mai_mai_n51_), .B(mai_mai_n106_), .Y(mai_mai_n341_));
  NO2        m0313(.A(mai_mai_n341_), .B(mai_mai_n340_), .Y(mai_mai_n342_));
  NA2        m0314(.A(mai_mai_n342_), .B(b), .Y(mai_mai_n343_));
  NA3        m0315(.A(mai_mai_n343_), .B(mai_mai_n338_), .C(mai_mai_n334_), .Y(mai_mai_n344_));
  NO4        m0316(.A(mai_mai_n344_), .B(mai_mai_n328_), .C(mai_mai_n314_), .D(mai_mai_n309_), .Y(mai_mai_n345_));
  NA4        m0317(.A(mai_mai_n345_), .B(mai_mai_n292_), .C(mai_mai_n249_), .D(mai_mai_n180_), .Y(mai10));
  NA3        m0318(.A(m), .B(k), .C(i), .Y(mai_mai_n347_));
  NO3        m0319(.A(mai_mai_n347_), .B(j), .C(mai_mai_n196_), .Y(mai_mai_n348_));
  NOi21      m0320(.An(e), .B(f), .Y(mai_mai_n349_));
  NO4        m0321(.A(mai_mai_n139_), .B(mai_mai_n349_), .C(n), .D(mai_mai_n103_), .Y(mai_mai_n350_));
  NAi31      m0322(.An(b), .B(f), .C(c), .Y(mai_mai_n351_));
  INV        m0323(.A(mai_mai_n351_), .Y(mai_mai_n352_));
  NOi32      m0324(.An(k), .Bn(h), .C(j), .Y(mai_mai_n353_));
  NA2        m0325(.A(mai_mai_n353_), .B(mai_mai_n203_), .Y(mai_mai_n354_));
  NA2        m0326(.A(mai_mai_n145_), .B(mai_mai_n354_), .Y(mai_mai_n355_));
  AOI220     m0327(.A0(mai_mai_n355_), .A1(mai_mai_n352_), .B0(mai_mai_n350_), .B1(mai_mai_n348_), .Y(mai_mai_n356_));
  AN2        m0328(.A(j), .B(h), .Y(mai_mai_n357_));
  OR2        m0329(.A(m), .B(k), .Y(mai_mai_n358_));
  NO2        m0330(.A(mai_mai_n156_), .B(mai_mai_n358_), .Y(mai_mai_n359_));
  NA4        m0331(.A(n), .B(f), .C(c), .D(mai_mai_n109_), .Y(mai_mai_n360_));
  NOi32      m0332(.An(d), .Bn(a), .C(c), .Y(mai_mai_n361_));
  NA2        m0333(.A(mai_mai_n361_), .B(mai_mai_n161_), .Y(mai_mai_n362_));
  NAi21      m0334(.An(i), .B(g), .Y(mai_mai_n363_));
  NAi31      m0335(.An(k), .B(m), .C(j), .Y(mai_mai_n364_));
  NO2        m0336(.A(mai_mai_n360_), .B(mai_mai_n275_), .Y(mai_mai_n365_));
  NOi32      m0337(.An(f), .Bn(d), .C(c), .Y(mai_mai_n366_));
  AOI220     m0338(.A0(mai_mai_n366_), .A1(mai_mai_n284_), .B0(mai_mai_n365_), .B1(mai_mai_n197_), .Y(mai_mai_n367_));
  NA2        m0339(.A(mai_mai_n367_), .B(mai_mai_n356_), .Y(mai_mai_n368_));
  NO2        m0340(.A(mai_mai_n57_), .B(mai_mai_n109_), .Y(mai_mai_n369_));
  NA2        m0341(.A(mai_mai_n231_), .B(mai_mai_n369_), .Y(mai_mai_n370_));
  INV        m0342(.A(e), .Y(mai_mai_n371_));
  NA2        m0343(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n372_));
  OAI220     m0344(.A0(mai_mai_n372_), .A1(mai_mai_n181_), .B0(mai_mai_n185_), .B1(mai_mai_n371_), .Y(mai_mai_n373_));
  AN2        m0345(.A(g), .B(e), .Y(mai_mai_n374_));
  NA3        m0346(.A(mai_mai_n374_), .B(mai_mai_n184_), .C(i), .Y(mai_mai_n375_));
  INV        m0347(.A(mai_mai_n375_), .Y(mai_mai_n376_));
  NO2        m0348(.A(mai_mai_n376_), .B(mai_mai_n373_), .Y(mai_mai_n377_));
  NOi32      m0349(.An(h), .Bn(e), .C(g), .Y(mai_mai_n378_));
  NA3        m0350(.A(mai_mai_n378_), .B(mai_mai_n272_), .C(m), .Y(mai_mai_n379_));
  NOi21      m0351(.An(g), .B(h), .Y(mai_mai_n380_));
  AN3        m0352(.A(m), .B(l), .C(i), .Y(mai_mai_n381_));
  NA3        m0353(.A(mai_mai_n381_), .B(mai_mai_n380_), .C(e), .Y(mai_mai_n382_));
  AN3        m0354(.A(h), .B(g), .C(e), .Y(mai_mai_n383_));
  NA2        m0355(.A(mai_mai_n383_), .B(mai_mai_n92_), .Y(mai_mai_n384_));
  AN3        m0356(.A(mai_mai_n384_), .B(mai_mai_n382_), .C(mai_mai_n379_), .Y(mai_mai_n385_));
  AOI210     m0357(.A0(mai_mai_n385_), .A1(mai_mai_n377_), .B0(mai_mai_n370_), .Y(mai_mai_n386_));
  NA3        m0358(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n387_));
  NO2        m0359(.A(mai_mai_n387_), .B(mai_mai_n370_), .Y(mai_mai_n388_));
  NA3        m0360(.A(mai_mai_n361_), .B(mai_mai_n161_), .C(mai_mai_n80_), .Y(mai_mai_n389_));
  NAi31      m0361(.An(b), .B(c), .C(a), .Y(mai_mai_n390_));
  NO2        m0362(.A(mai_mai_n390_), .B(n), .Y(mai_mai_n391_));
  OAI210     m0363(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n392_));
  NO2        m0364(.A(mai_mai_n392_), .B(e), .Y(mai_mai_n393_));
  NA2        m0365(.A(mai_mai_n393_), .B(mai_mai_n391_), .Y(mai_mai_n394_));
  INV        m0366(.A(mai_mai_n394_), .Y(mai_mai_n395_));
  NO4        m0367(.A(mai_mai_n395_), .B(mai_mai_n388_), .C(mai_mai_n386_), .D(mai_mai_n368_), .Y(mai_mai_n396_));
  NA2        m0368(.A(i), .B(g), .Y(mai_mai_n397_));
  NO3        m0369(.A(mai_mai_n258_), .B(mai_mai_n397_), .C(c), .Y(mai_mai_n398_));
  NOi21      m0370(.An(a), .B(n), .Y(mai_mai_n399_));
  NA2        m0371(.A(d), .B(mai_mai_n399_), .Y(mai_mai_n400_));
  NA3        m0372(.A(i), .B(g), .C(f), .Y(mai_mai_n401_));
  OR2        m0373(.A(mai_mai_n401_), .B(mai_mai_n66_), .Y(mai_mai_n402_));
  NA2        m0374(.A(mai_mai_n398_), .B(mai_mai_n271_), .Y(mai_mai_n403_));
  OR2        m0375(.A(n), .B(m), .Y(mai_mai_n404_));
  NO2        m0376(.A(mai_mai_n162_), .B(e), .Y(mai_mai_n405_));
  INV        m0377(.A(mai_mai_n341_), .Y(mai_mai_n406_));
  NA3        m0378(.A(mai_mai_n406_), .B(mai_mai_n335_), .C(d), .Y(mai_mai_n407_));
  NO2        m0379(.A(mai_mai_n390_), .B(mai_mai_n49_), .Y(mai_mai_n408_));
  NAi21      m0380(.An(k), .B(j), .Y(mai_mai_n409_));
  NAi21      m0381(.An(e), .B(d), .Y(mai_mai_n410_));
  INV        m0382(.A(mai_mai_n410_), .Y(mai_mai_n411_));
  NO2        m0383(.A(mai_mai_n234_), .B(mai_mai_n195_), .Y(mai_mai_n412_));
  NA3        m0384(.A(mai_mai_n412_), .B(mai_mai_n411_), .C(mai_mai_n209_), .Y(mai_mai_n413_));
  NA2        m0385(.A(mai_mai_n413_), .B(mai_mai_n407_), .Y(mai_mai_n414_));
  NOi31      m0386(.An(n), .B(m), .C(k), .Y(mai_mai_n415_));
  AOI220     m0387(.A0(mai_mai_n415_), .A1(mai_mai_n357_), .B0(mai_mai_n203_), .B1(mai_mai_n50_), .Y(mai_mai_n416_));
  NAi31      m0388(.An(g), .B(f), .C(c), .Y(mai_mai_n417_));
  OR3        m0389(.A(mai_mai_n417_), .B(mai_mai_n416_), .C(e), .Y(mai_mai_n418_));
  NA2        m0390(.A(mai_mai_n418_), .B(mai_mai_n285_), .Y(mai_mai_n419_));
  NOi41      m0391(.An(mai_mai_n403_), .B(mai_mai_n419_), .C(mai_mai_n414_), .D(mai_mai_n247_), .Y(mai_mai_n420_));
  NOi32      m0392(.An(c), .Bn(a), .C(b), .Y(mai_mai_n421_));
  NA2        m0393(.A(mai_mai_n421_), .B(mai_mai_n106_), .Y(mai_mai_n422_));
  INV        m0394(.A(mai_mai_n256_), .Y(mai_mai_n423_));
  AN2        m0395(.A(e), .B(d), .Y(mai_mai_n424_));
  NA2        m0396(.A(mai_mai_n424_), .B(mai_mai_n423_), .Y(mai_mai_n425_));
  NO2        m0397(.A(mai_mai_n122_), .B(mai_mai_n41_), .Y(mai_mai_n426_));
  NO2        m0398(.A(mai_mai_n61_), .B(e), .Y(mai_mai_n427_));
  NOi31      m0399(.An(j), .B(k), .C(i), .Y(mai_mai_n428_));
  NOi21      m0400(.An(mai_mai_n149_), .B(mai_mai_n428_), .Y(mai_mai_n429_));
  NA4        m0401(.A(mai_mai_n299_), .B(mai_mai_n429_), .C(mai_mai_n241_), .D(mai_mai_n112_), .Y(mai_mai_n430_));
  NA2        m0402(.A(mai_mai_n430_), .B(mai_mai_n427_), .Y(mai_mai_n431_));
  AOI210     m0403(.A0(mai_mai_n431_), .A1(mai_mai_n425_), .B0(mai_mai_n422_), .Y(mai_mai_n432_));
  NO2        m0404(.A(mai_mai_n191_), .B(mai_mai_n186_), .Y(mai_mai_n433_));
  NOi21      m0405(.An(a), .B(b), .Y(mai_mai_n434_));
  NA3        m0406(.A(e), .B(d), .C(c), .Y(mai_mai_n435_));
  NAi21      m0407(.An(mai_mai_n435_), .B(mai_mai_n434_), .Y(mai_mai_n436_));
  NO2        m0408(.A(mai_mai_n389_), .B(mai_mai_n185_), .Y(mai_mai_n437_));
  NOi21      m0409(.An(mai_mai_n436_), .B(mai_mai_n437_), .Y(mai_mai_n438_));
  AOI210     m0410(.A0(mai_mai_n250_), .A1(mai_mai_n433_), .B0(mai_mai_n438_), .Y(mai_mai_n439_));
  NO4        m0411(.A(mai_mai_n168_), .B(mai_mai_n96_), .C(mai_mai_n54_), .D(b), .Y(mai_mai_n440_));
  OR2        m0412(.A(k), .B(j), .Y(mai_mai_n441_));
  NA2        m0413(.A(l), .B(k), .Y(mai_mai_n442_));
  INV        m0414(.A(mai_mai_n261_), .Y(mai_mai_n443_));
  NA2        m0415(.A(mai_mai_n361_), .B(mai_mai_n106_), .Y(mai_mai_n444_));
  NO4        m0416(.A(mai_mai_n444_), .B(mai_mai_n89_), .C(mai_mai_n105_), .D(e), .Y(mai_mai_n445_));
  NO3        m0417(.A(mai_mai_n445_), .B(mai_mai_n443_), .C(mai_mai_n300_), .Y(mai_mai_n446_));
  INV        m0418(.A(mai_mai_n446_), .Y(mai_mai_n447_));
  NO4        m0419(.A(mai_mai_n447_), .B(mai_mai_n440_), .C(mai_mai_n439_), .D(mai_mai_n432_), .Y(mai_mai_n448_));
  NA2        m0420(.A(mai_mai_n65_), .B(mai_mai_n62_), .Y(mai_mai_n449_));
  NOi21      m0421(.An(d), .B(e), .Y(mai_mai_n450_));
  NAi31      m0422(.An(j), .B(l), .C(i), .Y(mai_mai_n451_));
  OAI210     m0423(.A0(mai_mai_n451_), .A1(mai_mai_n123_), .B0(mai_mai_n96_), .Y(mai_mai_n452_));
  NO3        m0424(.A(mai_mai_n362_), .B(mai_mai_n323_), .C(mai_mai_n182_), .Y(mai_mai_n453_));
  NO3        m0425(.A(mai_mai_n453_), .B(mai_mai_n164_), .C(mai_mai_n282_), .Y(mai_mai_n454_));
  NA3        m0426(.A(mai_mai_n454_), .B(mai_mai_n449_), .C(mai_mai_n226_), .Y(mai_mai_n455_));
  OAI210     m0427(.A0(mai_mai_n120_), .A1(mai_mai_n119_), .B0(n), .Y(mai_mai_n456_));
  NO2        m0428(.A(mai_mai_n456_), .B(mai_mai_n122_), .Y(mai_mai_n457_));
  OA210      m0429(.A0(mai_mai_n228_), .A1(mai_mai_n457_), .B0(mai_mai_n173_), .Y(mai_mai_n458_));
  XO2        m0430(.A(i), .B(h), .Y(mai_mai_n459_));
  NA3        m0431(.A(mai_mai_n459_), .B(mai_mai_n144_), .C(n), .Y(mai_mai_n460_));
  NAi41      m0432(.An(mai_mai_n276_), .B(mai_mai_n460_), .C(mai_mai_n416_), .D(mai_mai_n354_), .Y(mai_mai_n461_));
  NOi32      m0433(.An(mai_mai_n461_), .Bn(mai_mai_n427_), .C(mai_mai_n252_), .Y(mai_mai_n462_));
  NAi31      m0434(.An(c), .B(f), .C(d), .Y(mai_mai_n463_));
  AOI210     m0435(.A0(mai_mai_n262_), .A1(mai_mai_n176_), .B0(mai_mai_n463_), .Y(mai_mai_n464_));
  NOi21      m0436(.An(mai_mai_n78_), .B(mai_mai_n464_), .Y(mai_mai_n465_));
  NA3        m0437(.A(mai_mai_n350_), .B(mai_mai_n92_), .C(mai_mai_n91_), .Y(mai_mai_n466_));
  NA2        m0438(.A(mai_mai_n210_), .B(mai_mai_n101_), .Y(mai_mai_n467_));
  AOI210     m0439(.A0(mai_mai_n467_), .A1(mai_mai_n160_), .B0(mai_mai_n463_), .Y(mai_mai_n468_));
  NOi21      m0440(.An(mai_mai_n466_), .B(mai_mai_n468_), .Y(mai_mai_n469_));
  AO220      m0441(.A0(mai_mai_n268_), .A1(mai_mai_n244_), .B0(mai_mai_n150_), .B1(mai_mai_n62_), .Y(mai_mai_n470_));
  NA3        m0442(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n471_));
  NO2        m0443(.A(mai_mai_n471_), .B(mai_mai_n400_), .Y(mai_mai_n472_));
  INV        m0444(.A(mai_mai_n472_), .Y(mai_mai_n473_));
  NAi41      m0445(.An(mai_mai_n470_), .B(mai_mai_n473_), .C(mai_mai_n469_), .D(mai_mai_n465_), .Y(mai_mai_n474_));
  NO4        m0446(.A(mai_mai_n474_), .B(mai_mai_n462_), .C(mai_mai_n458_), .D(mai_mai_n455_), .Y(mai_mai_n475_));
  NA4        m0447(.A(mai_mai_n475_), .B(mai_mai_n448_), .C(mai_mai_n420_), .D(mai_mai_n396_), .Y(mai11));
  NO2        m0448(.A(mai_mai_n67_), .B(f), .Y(mai_mai_n477_));
  NA2        m0449(.A(j), .B(g), .Y(mai_mai_n478_));
  NAi31      m0450(.An(i), .B(m), .C(l), .Y(mai_mai_n479_));
  NA3        m0451(.A(m), .B(k), .C(j), .Y(mai_mai_n480_));
  OAI220     m0452(.A0(mai_mai_n480_), .A1(mai_mai_n122_), .B0(mai_mai_n479_), .B1(mai_mai_n478_), .Y(mai_mai_n481_));
  NA2        m0453(.A(mai_mai_n481_), .B(mai_mai_n477_), .Y(mai_mai_n482_));
  NOi32      m0454(.An(e), .Bn(b), .C(f), .Y(mai_mai_n483_));
  NA2        m0455(.A(mai_mai_n240_), .B(mai_mai_n106_), .Y(mai_mai_n484_));
  NA2        m0456(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n485_));
  NO2        m0457(.A(mai_mai_n485_), .B(mai_mai_n278_), .Y(mai_mai_n486_));
  NAi31      m0458(.An(d), .B(e), .C(a), .Y(mai_mai_n487_));
  NO2        m0459(.A(mai_mai_n487_), .B(n), .Y(mai_mai_n488_));
  NA2        m0460(.A(mai_mai_n486_), .B(mai_mai_n483_), .Y(mai_mai_n489_));
  NAi41      m0461(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n490_));
  AN2        m0462(.A(mai_mai_n490_), .B(mai_mai_n340_), .Y(mai_mai_n491_));
  NA2        m0463(.A(j), .B(i), .Y(mai_mai_n492_));
  NAi31      m0464(.An(n), .B(m), .C(k), .Y(mai_mai_n493_));
  NO3        m0465(.A(mai_mai_n493_), .B(mai_mai_n492_), .C(mai_mai_n105_), .Y(mai_mai_n494_));
  NO4        m0466(.A(n), .B(d), .C(mai_mai_n109_), .D(a), .Y(mai_mai_n495_));
  NO2        m0467(.A(n), .B(mai_mai_n137_), .Y(mai_mai_n496_));
  NO2        m0468(.A(mai_mai_n496_), .B(mai_mai_n495_), .Y(mai_mai_n497_));
  NOi32      m0469(.An(g), .Bn(f), .C(i), .Y(mai_mai_n498_));
  AOI220     m0470(.A0(mai_mai_n498_), .A1(mai_mai_n94_), .B0(mai_mai_n481_), .B1(f), .Y(mai_mai_n499_));
  NO2        m0471(.A(mai_mai_n256_), .B(mai_mai_n49_), .Y(mai_mai_n500_));
  NO2        m0472(.A(mai_mai_n499_), .B(mai_mai_n497_), .Y(mai_mai_n501_));
  INV        m0473(.A(mai_mai_n501_), .Y(mai_mai_n502_));
  NA2        m0474(.A(mai_mai_n131_), .B(mai_mai_n34_), .Y(mai_mai_n503_));
  OAI220     m0475(.A0(mai_mai_n503_), .A1(m), .B0(mai_mai_n485_), .B1(mai_mai_n216_), .Y(mai_mai_n504_));
  NOi41      m0476(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n505_));
  NAi32      m0477(.An(e), .Bn(b), .C(c), .Y(mai_mai_n506_));
  OR2        m0478(.A(mai_mai_n506_), .B(mai_mai_n80_), .Y(mai_mai_n507_));
  AN2        m0479(.A(mai_mai_n316_), .B(mai_mai_n296_), .Y(mai_mai_n508_));
  NA2        m0480(.A(mai_mai_n508_), .B(mai_mai_n507_), .Y(mai_mai_n509_));
  AN2        m0481(.A(mai_mai_n509_), .B(mai_mai_n504_), .Y(mai_mai_n510_));
  OAI220     m0482(.A0(mai_mai_n364_), .A1(mai_mai_n363_), .B0(mai_mai_n479_), .B1(mai_mai_n478_), .Y(mai_mai_n511_));
  NAi31      m0483(.An(d), .B(c), .C(a), .Y(mai_mai_n512_));
  NO2        m0484(.A(mai_mai_n512_), .B(n), .Y(mai_mai_n513_));
  NA3        m0485(.A(mai_mai_n513_), .B(mai_mai_n511_), .C(e), .Y(mai_mai_n514_));
  NO3        m0486(.A(mai_mai_n59_), .B(mai_mai_n49_), .C(mai_mai_n196_), .Y(mai_mai_n515_));
  INV        m0487(.A(mai_mai_n213_), .Y(mai_mai_n516_));
  NA2        m0488(.A(mai_mai_n515_), .B(mai_mai_n516_), .Y(mai_mai_n517_));
  NA2        m0489(.A(mai_mai_n517_), .B(mai_mai_n514_), .Y(mai_mai_n518_));
  INV        m0490(.A(mai_mai_n391_), .Y(mai_mai_n519_));
  NA2        m0491(.A(mai_mai_n511_), .B(f), .Y(mai_mai_n520_));
  NAi32      m0492(.An(d), .Bn(a), .C(b), .Y(mai_mai_n521_));
  INV        m0493(.A(mai_mai_n89_), .Y(mai_mai_n522_));
  NO3        m0494(.A(mai_mai_n158_), .B(mai_mai_n156_), .C(g), .Y(mai_mai_n523_));
  NA2        m0495(.A(mai_mai_n523_), .B(mai_mai_n56_), .Y(mai_mai_n524_));
  OAI210     m0496(.A0(mai_mai_n520_), .A1(mai_mai_n519_), .B0(mai_mai_n524_), .Y(mai_mai_n525_));
  AN3        m0497(.A(j), .B(h), .C(g), .Y(mai_mai_n526_));
  NO2        m0498(.A(mai_mai_n135_), .B(c), .Y(mai_mai_n527_));
  NA3        m0499(.A(mai_mai_n527_), .B(mai_mai_n526_), .C(mai_mai_n415_), .Y(mai_mai_n528_));
  NA3        m0500(.A(f), .B(d), .C(b), .Y(mai_mai_n529_));
  INV        m0501(.A(mai_mai_n528_), .Y(mai_mai_n530_));
  NO4        m0502(.A(mai_mai_n530_), .B(mai_mai_n525_), .C(mai_mai_n518_), .D(mai_mai_n510_), .Y(mai_mai_n531_));
  AN4        m0503(.A(mai_mai_n531_), .B(mai_mai_n502_), .C(mai_mai_n489_), .D(mai_mai_n482_), .Y(mai_mai_n532_));
  INV        m0504(.A(k), .Y(mai_mai_n533_));
  NA3        m0505(.A(l), .B(mai_mai_n533_), .C(i), .Y(mai_mai_n534_));
  INV        m0506(.A(mai_mai_n534_), .Y(mai_mai_n535_));
  NAi32      m0507(.An(h), .Bn(f), .C(g), .Y(mai_mai_n536_));
  NAi41      m0508(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n537_));
  OAI210     m0509(.A0(mai_mai_n487_), .A1(n), .B0(mai_mai_n537_), .Y(mai_mai_n538_));
  NA2        m0510(.A(mai_mai_n538_), .B(m), .Y(mai_mai_n539_));
  NAi31      m0511(.An(h), .B(g), .C(f), .Y(mai_mai_n540_));
  NO3        m0512(.A(mai_mai_n536_), .B(mai_mai_n67_), .C(mai_mai_n69_), .Y(mai_mai_n541_));
  NO4        m0513(.A(mai_mai_n540_), .B(n), .C(mai_mai_n137_), .D(mai_mai_n69_), .Y(mai_mai_n542_));
  OR2        m0514(.A(mai_mai_n542_), .B(mai_mai_n541_), .Y(mai_mai_n543_));
  NAi31      m0515(.An(f), .B(h), .C(g), .Y(mai_mai_n544_));
  NO4        m0516(.A(mai_mai_n287_), .B(mai_mai_n544_), .C(mai_mai_n67_), .D(mai_mai_n69_), .Y(mai_mai_n545_));
  NOi41      m0517(.An(b), .B(mai_mai_n329_), .C(mai_mai_n64_), .D(mai_mai_n110_), .Y(mai_mai_n546_));
  OR2        m0518(.A(mai_mai_n546_), .B(mai_mai_n545_), .Y(mai_mai_n547_));
  NOi32      m0519(.An(d), .Bn(a), .C(e), .Y(mai_mai_n548_));
  NA2        m0520(.A(mai_mai_n548_), .B(mai_mai_n106_), .Y(mai_mai_n549_));
  NO2        m0521(.A(n), .B(c), .Y(mai_mai_n550_));
  NA3        m0522(.A(mai_mai_n550_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n551_));
  NA2        m0523(.A(mai_mai_n551_), .B(mai_mai_n549_), .Y(mai_mai_n552_));
  INV        m0524(.A(mai_mai_n503_), .Y(mai_mai_n553_));
  AOI210     m0525(.A0(mai_mai_n553_), .A1(mai_mai_n552_), .B0(mai_mai_n547_), .Y(mai_mai_n554_));
  INV        m0526(.A(mai_mai_n554_), .Y(mai_mai_n555_));
  AOI210     m0527(.A0(mai_mai_n543_), .A1(mai_mai_n535_), .B0(mai_mai_n555_), .Y(mai_mai_n556_));
  NO3        m0528(.A(mai_mai_n294_), .B(mai_mai_n58_), .C(n), .Y(mai_mai_n557_));
  INV        m0529(.A(mai_mai_n463_), .Y(mai_mai_n558_));
  NA2        m0530(.A(mai_mai_n417_), .B(mai_mai_n213_), .Y(mai_mai_n559_));
  NA2        m0531(.A(mai_mai_n70_), .B(mai_mai_n106_), .Y(mai_mai_n560_));
  NA2        m0532(.A(mai_mai_n559_), .B(mai_mai_n557_), .Y(mai_mai_n561_));
  NO2        m0533(.A(mai_mai_n561_), .B(mai_mai_n83_), .Y(mai_mai_n562_));
  NA3        m0534(.A(mai_mai_n505_), .B(mai_mai_n318_), .C(mai_mai_n46_), .Y(mai_mai_n563_));
  NOi32      m0535(.An(e), .Bn(c), .C(f), .Y(mai_mai_n564_));
  NOi21      m0536(.An(f), .B(g), .Y(mai_mai_n565_));
  NO2        m0537(.A(mai_mai_n565_), .B(mai_mai_n193_), .Y(mai_mai_n566_));
  NA2        m0538(.A(mai_mai_n566_), .B(mai_mai_n359_), .Y(mai_mai_n567_));
  NA2        m0539(.A(mai_mai_n567_), .B(mai_mai_n563_), .Y(mai_mai_n568_));
  NOi21      m0540(.An(j), .B(l), .Y(mai_mai_n569_));
  NAi21      m0541(.An(k), .B(h), .Y(mai_mai_n570_));
  NO2        m0542(.A(mai_mai_n570_), .B(mai_mai_n243_), .Y(mai_mai_n571_));
  NA2        m0543(.A(mai_mai_n571_), .B(mai_mai_n569_), .Y(mai_mai_n572_));
  OR2        m0544(.A(mai_mai_n572_), .B(mai_mai_n539_), .Y(mai_mai_n573_));
  NOi31      m0545(.An(m), .B(n), .C(k), .Y(mai_mai_n574_));
  NA2        m0546(.A(mai_mai_n569_), .B(mai_mai_n574_), .Y(mai_mai_n575_));
  NO2        m0547(.A(mai_mai_n258_), .B(mai_mai_n49_), .Y(mai_mai_n576_));
  NO2        m0548(.A(mai_mai_n487_), .B(mai_mai_n49_), .Y(mai_mai_n577_));
  INV        m0549(.A(mai_mai_n573_), .Y(mai_mai_n578_));
  NA2        m0550(.A(mai_mai_n101_), .B(mai_mai_n36_), .Y(mai_mai_n579_));
  NO2        m0551(.A(k), .B(mai_mai_n196_), .Y(mai_mai_n580_));
  NO2        m0552(.A(mai_mai_n483_), .B(mai_mai_n335_), .Y(mai_mai_n581_));
  NO2        m0553(.A(mai_mai_n581_), .B(n), .Y(mai_mai_n582_));
  NAi31      m0554(.An(mai_mai_n579_), .B(mai_mai_n582_), .C(mai_mai_n580_), .Y(mai_mai_n583_));
  NO2        m0555(.A(mai_mai_n485_), .B(mai_mai_n158_), .Y(mai_mai_n584_));
  NA3        m0556(.A(mai_mai_n506_), .B(mai_mai_n252_), .C(mai_mai_n134_), .Y(mai_mai_n585_));
  NA2        m0557(.A(mai_mai_n459_), .B(mai_mai_n144_), .Y(mai_mai_n586_));
  NO3        m0558(.A(mai_mai_n360_), .B(mai_mai_n586_), .C(mai_mai_n83_), .Y(mai_mai_n587_));
  AOI210     m0559(.A0(mai_mai_n585_), .A1(mai_mai_n584_), .B0(mai_mai_n587_), .Y(mai_mai_n588_));
  AN3        m0560(.A(f), .B(d), .C(b), .Y(mai_mai_n589_));
  OAI210     m0561(.A0(mai_mai_n589_), .A1(mai_mai_n121_), .B0(n), .Y(mai_mai_n590_));
  NA3        m0562(.A(mai_mai_n459_), .B(mai_mai_n144_), .C(mai_mai_n196_), .Y(mai_mai_n591_));
  AOI210     m0563(.A0(mai_mai_n590_), .A1(mai_mai_n215_), .B0(mai_mai_n591_), .Y(mai_mai_n592_));
  NAi31      m0564(.An(m), .B(n), .C(k), .Y(mai_mai_n593_));
  OR2        m0565(.A(mai_mai_n126_), .B(mai_mai_n58_), .Y(mai_mai_n594_));
  OAI210     m0566(.A0(mai_mai_n594_), .A1(mai_mai_n593_), .B0(mai_mai_n232_), .Y(mai_mai_n595_));
  OAI210     m0567(.A0(mai_mai_n595_), .A1(mai_mai_n592_), .B0(j), .Y(mai_mai_n596_));
  NA3        m0568(.A(mai_mai_n596_), .B(mai_mai_n588_), .C(mai_mai_n583_), .Y(mai_mai_n597_));
  NO4        m0569(.A(mai_mai_n597_), .B(mai_mai_n578_), .C(mai_mai_n568_), .D(mai_mai_n562_), .Y(mai_mai_n598_));
  NAi31      m0570(.An(g), .B(h), .C(f), .Y(mai_mai_n599_));
  OR3        m0571(.A(mai_mai_n599_), .B(mai_mai_n258_), .C(n), .Y(mai_mai_n600_));
  NA3        m0572(.A(mai_mai_n378_), .B(mai_mai_n114_), .C(mai_mai_n80_), .Y(mai_mai_n601_));
  NO3        m0573(.A(g), .B(mai_mai_n195_), .C(mai_mai_n54_), .Y(mai_mai_n602_));
  NAi21      m0574(.An(h), .B(j), .Y(mai_mai_n603_));
  NO2        m0575(.A(mai_mai_n467_), .B(mai_mai_n83_), .Y(mai_mai_n604_));
  OAI210     m0576(.A0(mai_mai_n604_), .A1(mai_mai_n359_), .B0(mai_mai_n602_), .Y(mai_mai_n605_));
  BUFFER     m0577(.A(mai_mai_n67_), .Y(mai_mai_n606_));
  NA2        m0578(.A(b), .B(mai_mai_n320_), .Y(mai_mai_n607_));
  OA220      m0579(.A0(mai_mai_n575_), .A1(mai_mai_n607_), .B0(mai_mai_n572_), .B1(mai_mai_n606_), .Y(mai_mai_n608_));
  NA3        m0580(.A(mai_mai_n477_), .B(mai_mai_n94_), .C(mai_mai_n93_), .Y(mai_mai_n609_));
  NA2        m0581(.A(h), .B(mai_mai_n37_), .Y(mai_mai_n610_));
  NA2        m0582(.A(mai_mai_n94_), .B(mai_mai_n46_), .Y(mai_mai_n611_));
  OAI220     m0583(.A0(mai_mai_n611_), .A1(mai_mai_n311_), .B0(mai_mai_n610_), .B1(mai_mai_n422_), .Y(mai_mai_n612_));
  AOI210     m0584(.A0(mai_mai_n521_), .A1(mai_mai_n390_), .B0(mai_mai_n49_), .Y(mai_mai_n613_));
  OAI220     m0585(.A0(mai_mai_n540_), .A1(mai_mai_n534_), .B0(mai_mai_n304_), .B1(mai_mai_n478_), .Y(mai_mai_n614_));
  AOI210     m0586(.A0(mai_mai_n614_), .A1(mai_mai_n613_), .B0(mai_mai_n612_), .Y(mai_mai_n615_));
  NA4        m0587(.A(mai_mai_n615_), .B(mai_mai_n609_), .C(mai_mai_n608_), .D(mai_mai_n605_), .Y(mai_mai_n616_));
  NO2        m0588(.A(mai_mai_n233_), .B(f), .Y(mai_mai_n617_));
  INV        m0589(.A(mai_mai_n58_), .Y(mai_mai_n618_));
  NO3        m0590(.A(mai_mai_n618_), .B(mai_mai_n617_), .C(mai_mai_n34_), .Y(mai_mai_n619_));
  NA2        m0591(.A(mai_mai_n307_), .B(mai_mai_n131_), .Y(mai_mai_n620_));
  NA2        m0592(.A(mai_mai_n1343_), .B(mai_mai_n483_), .Y(mai_mai_n621_));
  OR2        m0593(.A(mai_mai_n621_), .B(mai_mai_n503_), .Y(mai_mai_n622_));
  OAI210     m0594(.A0(mai_mai_n620_), .A1(mai_mai_n619_), .B0(mai_mai_n622_), .Y(mai_mai_n623_));
  NO2        m0595(.A(mai_mai_n366_), .B(mai_mai_n173_), .Y(mai_mai_n624_));
  NA2        m0596(.A(mai_mai_n624_), .B(mai_mai_n213_), .Y(mai_mai_n625_));
  NA3        m0597(.A(mai_mai_n625_), .B(mai_mai_n235_), .C(j), .Y(mai_mai_n626_));
  NA2        m0598(.A(mai_mai_n421_), .B(mai_mai_n80_), .Y(mai_mai_n627_));
  NO4        m0599(.A(mai_mai_n480_), .B(mai_mai_n627_), .C(mai_mai_n122_), .D(mai_mai_n195_), .Y(mai_mai_n628_));
  INV        m0600(.A(mai_mai_n628_), .Y(mai_mai_n629_));
  NA3        m0601(.A(mai_mai_n629_), .B(mai_mai_n626_), .C(mai_mai_n466_), .Y(mai_mai_n630_));
  NO3        m0602(.A(mai_mai_n630_), .B(mai_mai_n623_), .C(mai_mai_n616_), .Y(mai_mai_n631_));
  NA4        m0603(.A(mai_mai_n631_), .B(mai_mai_n598_), .C(mai_mai_n556_), .D(mai_mai_n532_), .Y(mai08));
  NO2        m0604(.A(k), .B(h), .Y(mai_mai_n633_));
  AO210      m0605(.A0(mai_mai_n233_), .A1(mai_mai_n409_), .B0(mai_mai_n633_), .Y(mai_mai_n634_));
  NO2        m0606(.A(mai_mai_n634_), .B(mai_mai_n275_), .Y(mai_mai_n635_));
  NA2        m0607(.A(mai_mai_n564_), .B(mai_mai_n80_), .Y(mai_mai_n636_));
  NA2        m0608(.A(mai_mai_n636_), .B(mai_mai_n417_), .Y(mai_mai_n637_));
  NA2        m0609(.A(mai_mai_n637_), .B(mai_mai_n635_), .Y(mai_mai_n638_));
  NA2        m0610(.A(mai_mai_n80_), .B(mai_mai_n103_), .Y(mai_mai_n639_));
  NO2        m0611(.A(mai_mai_n639_), .B(mai_mai_n55_), .Y(mai_mai_n640_));
  NA2        m0612(.A(mai_mai_n529_), .B(mai_mai_n215_), .Y(mai_mai_n641_));
  NA2        m0613(.A(mai_mai_n641_), .B(mai_mai_n325_), .Y(mai_mai_n642_));
  AOI210     m0614(.A0(mai_mai_n529_), .A1(mai_mai_n142_), .B0(mai_mai_n80_), .Y(mai_mai_n643_));
  NA4        m0615(.A(mai_mai_n198_), .B(mai_mai_n131_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n644_));
  AN2        m0616(.A(l), .B(k), .Y(mai_mai_n645_));
  NA4        m0617(.A(mai_mai_n645_), .B(mai_mai_n101_), .C(mai_mai_n69_), .D(mai_mai_n196_), .Y(mai_mai_n646_));
  OAI210     m0618(.A0(mai_mai_n644_), .A1(g), .B0(mai_mai_n646_), .Y(mai_mai_n647_));
  NA2        m0619(.A(mai_mai_n647_), .B(mai_mai_n643_), .Y(mai_mai_n648_));
  NA3        m0620(.A(mai_mai_n648_), .B(mai_mai_n642_), .C(mai_mai_n638_), .Y(mai_mai_n649_));
  AN2        m0621(.A(mai_mai_n488_), .B(mai_mai_n90_), .Y(mai_mai_n650_));
  INV        m0622(.A(mai_mai_n472_), .Y(mai_mai_n651_));
  NO2        m0623(.A(mai_mai_n38_), .B(mai_mai_n195_), .Y(mai_mai_n652_));
  NA2        m0624(.A(mai_mai_n566_), .B(mai_mai_n324_), .Y(mai_mai_n653_));
  NA2        m0625(.A(mai_mai_n653_), .B(mai_mai_n651_), .Y(mai_mai_n654_));
  NO2        m0626(.A(mai_mai_n491_), .B(mai_mai_n35_), .Y(mai_mai_n655_));
  OAI210     m0627(.A0(mai_mai_n506_), .A1(mai_mai_n47_), .B0(mai_mai_n594_), .Y(mai_mai_n656_));
  NO2        m0628(.A(mai_mai_n442_), .B(mai_mai_n123_), .Y(mai_mai_n657_));
  AOI210     m0629(.A0(mai_mai_n657_), .A1(mai_mai_n656_), .B0(mai_mai_n655_), .Y(mai_mai_n658_));
  INV        m0630(.A(mai_mai_n658_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n335_), .B(mai_mai_n43_), .Y(mai_mai_n660_));
  NA3        m0632(.A(mai_mai_n625_), .B(mai_mai_n313_), .C(mai_mai_n353_), .Y(mai_mai_n661_));
  NA2        m0633(.A(mai_mai_n645_), .B(mai_mai_n203_), .Y(mai_mai_n662_));
  NO2        m0634(.A(mai_mai_n662_), .B(mai_mai_n306_), .Y(mai_mai_n663_));
  AOI210     m0635(.A0(mai_mai_n663_), .A1(mai_mai_n617_), .B0(mai_mai_n445_), .Y(mai_mai_n664_));
  NA3        m0636(.A(m), .B(l), .C(k), .Y(mai_mai_n665_));
  AOI210     m0637(.A0(mai_mai_n601_), .A1(mai_mai_n600_), .B0(mai_mai_n665_), .Y(mai_mai_n666_));
  NO2        m0638(.A(mai_mai_n490_), .B(mai_mai_n253_), .Y(mai_mai_n667_));
  NOi21      m0639(.An(mai_mai_n667_), .B(mai_mai_n484_), .Y(mai_mai_n668_));
  NA4        m0640(.A(mai_mai_n106_), .B(l), .C(k), .D(mai_mai_n83_), .Y(mai_mai_n669_));
  NO2        m0641(.A(mai_mai_n668_), .B(mai_mai_n666_), .Y(mai_mai_n670_));
  NA4        m0642(.A(mai_mai_n670_), .B(mai_mai_n664_), .C(mai_mai_n661_), .D(mai_mai_n660_), .Y(mai_mai_n671_));
  NO4        m0643(.A(mai_mai_n671_), .B(mai_mai_n659_), .C(mai_mai_n654_), .D(mai_mai_n649_), .Y(mai_mai_n672_));
  NA2        m0644(.A(mai_mai_n566_), .B(mai_mai_n359_), .Y(mai_mai_n673_));
  NOi31      m0645(.An(g), .B(h), .C(f), .Y(mai_mai_n674_));
  NA2        m0646(.A(mai_mai_n577_), .B(mai_mai_n674_), .Y(mai_mai_n675_));
  NA3        m0647(.A(mai_mai_n675_), .B(mai_mai_n673_), .C(mai_mai_n232_), .Y(mai_mai_n676_));
  NOi21      m0648(.An(h), .B(j), .Y(mai_mai_n677_));
  NA2        m0649(.A(mai_mai_n677_), .B(f), .Y(mai_mai_n678_));
  NA2        m0650(.A(mai_mai_n676_), .B(l), .Y(mai_mai_n679_));
  NO2        m0651(.A(j), .B(i), .Y(mai_mai_n680_));
  NA2        m0652(.A(mai_mai_n680_), .B(mai_mai_n33_), .Y(mai_mai_n681_));
  NA2        m0653(.A(mai_mai_n383_), .B(mai_mai_n114_), .Y(mai_mai_n682_));
  OR2        m0654(.A(mai_mai_n682_), .B(mai_mai_n681_), .Y(mai_mai_n683_));
  NO3        m0655(.A(mai_mai_n139_), .B(mai_mai_n49_), .C(mai_mai_n103_), .Y(mai_mai_n684_));
  NO3        m0656(.A(n), .B(mai_mai_n137_), .C(mai_mai_n69_), .Y(mai_mai_n685_));
  NO3        m0657(.A(mai_mai_n442_), .B(mai_mai_n401_), .C(j), .Y(mai_mai_n686_));
  OAI210     m0658(.A0(mai_mai_n685_), .A1(mai_mai_n684_), .B0(mai_mai_n686_), .Y(mai_mai_n687_));
  OAI210     m0659(.A0(mai_mai_n675_), .A1(mai_mai_n59_), .B0(mai_mai_n687_), .Y(mai_mai_n688_));
  NA2        m0660(.A(k), .B(j), .Y(mai_mai_n689_));
  NO3        m0661(.A(mai_mai_n275_), .B(mai_mai_n689_), .C(mai_mai_n40_), .Y(mai_mai_n690_));
  AOI210     m0662(.A0(mai_mai_n483_), .A1(n), .B0(mai_mai_n505_), .Y(mai_mai_n691_));
  NA2        m0663(.A(mai_mai_n691_), .B(mai_mai_n508_), .Y(mai_mai_n692_));
  AN3        m0664(.A(mai_mai_n692_), .B(mai_mai_n690_), .C(mai_mai_n93_), .Y(mai_mai_n693_));
  NO2        m0665(.A(mai_mai_n275_), .B(mai_mai_n127_), .Y(mai_mai_n694_));
  NA2        m0666(.A(mai_mai_n694_), .B(mai_mai_n566_), .Y(mai_mai_n695_));
  NO2        m0667(.A(mai_mai_n665_), .B(mai_mai_n86_), .Y(mai_mai_n696_));
  NA2        m0668(.A(mai_mai_n696_), .B(mai_mai_n538_), .Y(mai_mai_n697_));
  NO2        m0669(.A(mai_mai_n540_), .B(mai_mai_n110_), .Y(mai_mai_n698_));
  OAI210     m0670(.A0(mai_mai_n698_), .A1(mai_mai_n686_), .B0(mai_mai_n613_), .Y(mai_mai_n699_));
  NA3        m0671(.A(mai_mai_n699_), .B(mai_mai_n697_), .C(mai_mai_n695_), .Y(mai_mai_n700_));
  OR3        m0672(.A(mai_mai_n700_), .B(mai_mai_n693_), .C(mai_mai_n688_), .Y(mai_mai_n701_));
  NA3        m0673(.A(mai_mai_n691_), .B(mai_mai_n508_), .C(mai_mai_n507_), .Y(mai_mai_n702_));
  NA4        m0674(.A(mai_mai_n702_), .B(mai_mai_n198_), .C(mai_mai_n409_), .D(mai_mai_n34_), .Y(mai_mai_n703_));
  OAI220     m0675(.A0(mai_mai_n644_), .A1(mai_mai_n636_), .B0(mai_mai_n311_), .B1(mai_mai_n38_), .Y(mai_mai_n704_));
  INV        m0676(.A(mai_mai_n704_), .Y(mai_mai_n705_));
  NA3        m0677(.A(mai_mai_n498_), .B(mai_mai_n272_), .C(h), .Y(mai_mai_n706_));
  NO2        m0678(.A(mai_mai_n87_), .B(mai_mai_n47_), .Y(mai_mai_n707_));
  NO2        m0679(.A(mai_mai_n706_), .B(mai_mai_n551_), .Y(mai_mai_n708_));
  AOI210     m0680(.A0(mai_mai_n707_), .A1(mai_mai_n582_), .B0(mai_mai_n708_), .Y(mai_mai_n709_));
  NA3        m0681(.A(mai_mai_n709_), .B(mai_mai_n705_), .C(mai_mai_n703_), .Y(mai_mai_n710_));
  OR2        m0682(.A(mai_mai_n696_), .B(mai_mai_n90_), .Y(mai_mai_n711_));
  NA2        m0683(.A(mai_mai_n711_), .B(mai_mai_n221_), .Y(mai_mai_n712_));
  OAI210     m0684(.A0(mai_mai_n665_), .A1(mai_mai_n599_), .B0(mai_mai_n471_), .Y(mai_mai_n713_));
  NA3        m0685(.A(mai_mai_n231_), .B(mai_mai_n57_), .C(b), .Y(mai_mai_n714_));
  AOI220     m0686(.A0(mai_mai_n550_), .A1(mai_mai_n29_), .B0(mai_mai_n421_), .B1(mai_mai_n80_), .Y(mai_mai_n715_));
  NA2        m0687(.A(mai_mai_n715_), .B(mai_mai_n714_), .Y(mai_mai_n716_));
  NO2        m0688(.A(mai_mai_n706_), .B(mai_mai_n444_), .Y(mai_mai_n717_));
  AOI210     m0689(.A0(mai_mai_n716_), .A1(mai_mai_n713_), .B0(mai_mai_n717_), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n718_), .B(mai_mai_n712_), .Y(mai_mai_n719_));
  NOi41      m0691(.An(mai_mai_n683_), .B(mai_mai_n719_), .C(mai_mai_n710_), .D(mai_mai_n701_), .Y(mai_mai_n720_));
  OR3        m0692(.A(mai_mai_n644_), .B(mai_mai_n215_), .C(g), .Y(mai_mai_n721_));
  NO3        m0693(.A(mai_mai_n319_), .B(mai_mai_n277_), .C(mai_mai_n105_), .Y(mai_mai_n722_));
  NA2        m0694(.A(mai_mai_n722_), .B(mai_mai_n692_), .Y(mai_mai_n723_));
  INV        m0695(.A(mai_mai_n46_), .Y(mai_mai_n724_));
  NO3        m0696(.A(mai_mai_n724_), .B(mai_mai_n681_), .C(mai_mai_n258_), .Y(mai_mai_n725_));
  INV        m0697(.A(mai_mai_n725_), .Y(mai_mai_n726_));
  NA4        m0698(.A(mai_mai_n726_), .B(mai_mai_n723_), .C(mai_mai_n721_), .D(mai_mai_n367_), .Y(mai_mai_n727_));
  OR2        m0699(.A(mai_mai_n599_), .B(mai_mai_n87_), .Y(mai_mai_n728_));
  NOi31      m0700(.An(b), .B(d), .C(a), .Y(mai_mai_n729_));
  NO2        m0701(.A(mai_mai_n729_), .B(mai_mai_n548_), .Y(mai_mai_n730_));
  NO2        m0702(.A(mai_mai_n730_), .B(n), .Y(mai_mai_n731_));
  NOi21      m0703(.An(mai_mai_n715_), .B(mai_mai_n731_), .Y(mai_mai_n732_));
  NO2        m0704(.A(mai_mai_n732_), .B(mai_mai_n728_), .Y(mai_mai_n733_));
  NO2        m0705(.A(mai_mai_n506_), .B(mai_mai_n80_), .Y(mai_mai_n734_));
  NO2        m0706(.A(mai_mai_n306_), .B(mai_mai_n110_), .Y(mai_mai_n735_));
  NOi21      m0707(.An(mai_mai_n735_), .B(mai_mai_n145_), .Y(mai_mai_n736_));
  AOI210     m0708(.A0(mai_mai_n722_), .A1(mai_mai_n734_), .B0(mai_mai_n736_), .Y(mai_mai_n737_));
  OAI210     m0709(.A0(mai_mai_n644_), .A1(mai_mai_n360_), .B0(mai_mai_n737_), .Y(mai_mai_n738_));
  NA2        m0710(.A(mai_mai_n694_), .B(mai_mai_n602_), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n114_), .B(mai_mai_n80_), .Y(mai_mai_n740_));
  AOI210     m0712(.A0(mai_mai_n387_), .A1(mai_mai_n379_), .B0(mai_mai_n740_), .Y(mai_mai_n741_));
  NA2        m0713(.A(mai_mai_n663_), .B(mai_mai_n34_), .Y(mai_mai_n742_));
  NAi21      m0714(.An(mai_mai_n669_), .B(mai_mai_n398_), .Y(mai_mai_n743_));
  NO2        m0715(.A(mai_mai_n253_), .B(i), .Y(mai_mai_n744_));
  OAI210     m0716(.A0(mai_mai_n542_), .A1(mai_mai_n541_), .B0(mai_mai_n336_), .Y(mai_mai_n745_));
  AN2        m0717(.A(mai_mai_n745_), .B(mai_mai_n743_), .Y(mai_mai_n746_));
  NAi41      m0718(.An(mai_mai_n741_), .B(mai_mai_n746_), .C(mai_mai_n742_), .D(mai_mai_n739_), .Y(mai_mai_n747_));
  NO4        m0719(.A(mai_mai_n747_), .B(mai_mai_n738_), .C(mai_mai_n733_), .D(mai_mai_n727_), .Y(mai_mai_n748_));
  NA4        m0720(.A(mai_mai_n748_), .B(mai_mai_n720_), .C(mai_mai_n679_), .D(mai_mai_n672_), .Y(mai09));
  INV        m0721(.A(mai_mai_n115_), .Y(mai_mai_n750_));
  NA2        m0722(.A(f), .B(e), .Y(mai_mai_n751_));
  NO2        m0723(.A(mai_mai_n208_), .B(mai_mai_n105_), .Y(mai_mai_n752_));
  NA4        m0724(.A(mai_mai_n287_), .B(mai_mai_n429_), .C(mai_mai_n241_), .D(mai_mai_n112_), .Y(mai_mai_n753_));
  AOI210     m0725(.A0(mai_mai_n753_), .A1(g), .B0(mai_mai_n426_), .Y(mai_mai_n754_));
  NO2        m0726(.A(mai_mai_n754_), .B(mai_mai_n751_), .Y(mai_mai_n755_));
  NA2        m0727(.A(mai_mai_n755_), .B(mai_mai_n750_), .Y(mai_mai_n756_));
  NO2        m0728(.A(mai_mai_n185_), .B(mai_mai_n195_), .Y(mai_mai_n757_));
  NA3        m0729(.A(m), .B(l), .C(i), .Y(mai_mai_n758_));
  OAI220     m0730(.A0(mai_mai_n540_), .A1(mai_mai_n758_), .B0(mai_mai_n329_), .B1(mai_mai_n479_), .Y(mai_mai_n759_));
  NA4        m0731(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(g), .D(f), .Y(mai_mai_n760_));
  NAi31      m0732(.An(mai_mai_n759_), .B(mai_mai_n760_), .C(mai_mai_n402_), .Y(mai_mai_n761_));
  OR2        m0733(.A(mai_mai_n761_), .B(mai_mai_n757_), .Y(mai_mai_n762_));
  NA3        m0734(.A(mai_mai_n728_), .B(mai_mai_n520_), .C(mai_mai_n471_), .Y(mai_mai_n763_));
  OA210      m0735(.A0(mai_mai_n763_), .A1(mai_mai_n762_), .B0(mai_mai_n731_), .Y(mai_mai_n764_));
  INV        m0736(.A(mai_mai_n316_), .Y(mai_mai_n765_));
  NO2        m0737(.A(mai_mai_n120_), .B(mai_mai_n119_), .Y(mai_mai_n766_));
  NOi31      m0738(.An(k), .B(m), .C(l), .Y(mai_mai_n767_));
  NO2        m0739(.A(mai_mai_n318_), .B(mai_mai_n767_), .Y(mai_mai_n768_));
  AOI210     m0740(.A0(mai_mai_n768_), .A1(mai_mai_n766_), .B0(mai_mai_n544_), .Y(mai_mai_n769_));
  NA2        m0741(.A(mai_mai_n714_), .B(mai_mai_n311_), .Y(mai_mai_n770_));
  NA2        m0742(.A(mai_mai_n320_), .B(mai_mai_n322_), .Y(mai_mai_n771_));
  OAI210     m0743(.A0(mai_mai_n185_), .A1(mai_mai_n195_), .B0(mai_mai_n771_), .Y(mai_mai_n772_));
  AOI220     m0744(.A0(mai_mai_n772_), .A1(mai_mai_n770_), .B0(mai_mai_n769_), .B1(mai_mai_n765_), .Y(mai_mai_n773_));
  NA2        m0745(.A(mai_mai_n153_), .B(mai_mai_n107_), .Y(mai_mai_n774_));
  NA3        m0746(.A(mai_mai_n774_), .B(mai_mai_n634_), .C(mai_mai_n127_), .Y(mai_mai_n775_));
  NA3        m0747(.A(mai_mai_n775_), .B(mai_mai_n170_), .C(mai_mai_n31_), .Y(mai_mai_n776_));
  NA4        m0748(.A(mai_mai_n776_), .B(mai_mai_n773_), .C(mai_mai_n567_), .D(mai_mai_n78_), .Y(mai_mai_n777_));
  NO2        m0749(.A(mai_mai_n536_), .B(mai_mai_n451_), .Y(mai_mai_n778_));
  NA2        m0750(.A(mai_mai_n778_), .B(mai_mai_n170_), .Y(mai_mai_n779_));
  NOi21      m0751(.An(f), .B(d), .Y(mai_mai_n780_));
  NA2        m0752(.A(mai_mai_n780_), .B(m), .Y(mai_mai_n781_));
  NOi32      m0753(.An(g), .Bn(f), .C(d), .Y(mai_mai_n782_));
  NA4        m0754(.A(mai_mai_n782_), .B(mai_mai_n550_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n783_));
  NA3        m0755(.A(mai_mai_n287_), .B(mai_mai_n241_), .C(mai_mai_n112_), .Y(mai_mai_n784_));
  AN2        m0756(.A(f), .B(d), .Y(mai_mai_n785_));
  NA3        m0757(.A(mai_mai_n434_), .B(mai_mai_n785_), .C(mai_mai_n80_), .Y(mai_mai_n786_));
  NO3        m0758(.A(mai_mai_n786_), .B(mai_mai_n69_), .C(mai_mai_n196_), .Y(mai_mai_n787_));
  NO2        m0759(.A(mai_mai_n265_), .B(mai_mai_n54_), .Y(mai_mai_n788_));
  NA2        m0760(.A(mai_mai_n784_), .B(mai_mai_n787_), .Y(mai_mai_n789_));
  NAi31      m0761(.An(mai_mai_n443_), .B(mai_mai_n789_), .C(mai_mai_n779_), .Y(mai_mai_n790_));
  NO4        m0762(.A(mai_mai_n565_), .B(mai_mai_n123_), .C(mai_mai_n306_), .D(mai_mai_n140_), .Y(mai_mai_n791_));
  NO2        m0763(.A(mai_mai_n593_), .B(mai_mai_n306_), .Y(mai_mai_n792_));
  AN2        m0764(.A(mai_mai_n792_), .B(mai_mai_n617_), .Y(mai_mai_n793_));
  NO3        m0765(.A(mai_mai_n793_), .B(mai_mai_n791_), .C(mai_mai_n217_), .Y(mai_mai_n794_));
  NA2        m0766(.A(mai_mai_n548_), .B(mai_mai_n80_), .Y(mai_mai_n795_));
  NO2        m0767(.A(mai_mai_n771_), .B(mai_mai_n795_), .Y(mai_mai_n796_));
  NA3        m0768(.A(mai_mai_n144_), .B(mai_mai_n101_), .C(g), .Y(mai_mai_n797_));
  OAI220     m0769(.A0(mai_mai_n786_), .A1(mai_mai_n392_), .B0(mai_mai_n316_), .B1(mai_mai_n797_), .Y(mai_mai_n798_));
  NOi41      m0770(.An(mai_mai_n206_), .B(mai_mai_n798_), .C(mai_mai_n796_), .D(mai_mai_n282_), .Y(mai_mai_n799_));
  NA2        m0771(.A(c), .B(mai_mai_n109_), .Y(mai_mai_n800_));
  NO2        m0772(.A(mai_mai_n800_), .B(mai_mai_n371_), .Y(mai_mai_n801_));
  NA3        m0773(.A(mai_mai_n801_), .B(mai_mai_n461_), .C(f), .Y(mai_mai_n802_));
  OR2        m0774(.A(mai_mai_n599_), .B(mai_mai_n493_), .Y(mai_mai_n803_));
  INV        m0775(.A(mai_mai_n803_), .Y(mai_mai_n804_));
  NA2        m0776(.A(mai_mai_n730_), .B(mai_mai_n104_), .Y(mai_mai_n805_));
  NA2        m0777(.A(mai_mai_n805_), .B(mai_mai_n804_), .Y(mai_mai_n806_));
  NA4        m0778(.A(mai_mai_n806_), .B(mai_mai_n802_), .C(mai_mai_n799_), .D(mai_mai_n794_), .Y(mai_mai_n807_));
  NO4        m0779(.A(mai_mai_n807_), .B(mai_mai_n790_), .C(mai_mai_n777_), .D(mai_mai_n764_), .Y(mai_mai_n808_));
  NO2        m0780(.A(mai_mai_n392_), .B(mai_mai_n751_), .Y(mai_mai_n809_));
  NA2        m0781(.A(mai_mai_n809_), .B(mai_mai_n513_), .Y(mai_mai_n810_));
  INV        m0782(.A(mai_mai_n810_), .Y(mai_mai_n811_));
  NA2        m0783(.A(e), .B(d), .Y(mai_mai_n812_));
  OAI220     m0784(.A0(mai_mai_n812_), .A1(c), .B0(mai_mai_n301_), .B1(d), .Y(mai_mai_n813_));
  NA3        m0785(.A(mai_mai_n813_), .B(mai_mai_n412_), .C(mai_mai_n459_), .Y(mai_mai_n814_));
  AOI210     m0786(.A0(mai_mai_n467_), .A1(mai_mai_n160_), .B0(mai_mai_n213_), .Y(mai_mai_n815_));
  AOI210     m0787(.A0(mai_mai_n566_), .A1(mai_mai_n324_), .B0(mai_mai_n815_), .Y(mai_mai_n816_));
  NA2        m0788(.A(mai_mai_n265_), .B(mai_mai_n149_), .Y(mai_mai_n817_));
  NA2        m0789(.A(mai_mai_n787_), .B(mai_mai_n817_), .Y(mai_mai_n818_));
  NA3        m0790(.A(mai_mai_n152_), .B(mai_mai_n81_), .C(mai_mai_n34_), .Y(mai_mai_n819_));
  NA4        m0791(.A(mai_mai_n819_), .B(mai_mai_n818_), .C(mai_mai_n816_), .D(mai_mai_n814_), .Y(mai_mai_n820_));
  NO2        m0792(.A(mai_mai_n820_), .B(mai_mai_n811_), .Y(mai_mai_n821_));
  NA2        m0793(.A(mai_mai_n765_), .B(mai_mai_n31_), .Y(mai_mai_n822_));
  OR2        m0794(.A(mai_mai_n822_), .B(mai_mai_n199_), .Y(mai_mai_n823_));
  OAI220     m0795(.A0(mai_mai_n565_), .A1(mai_mai_n58_), .B0(mai_mai_n277_), .B1(j), .Y(mai_mai_n824_));
  AOI220     m0796(.A0(mai_mai_n824_), .A1(mai_mai_n792_), .B0(mai_mai_n557_), .B1(mai_mai_n564_), .Y(mai_mai_n825_));
  INV        m0797(.A(mai_mai_n825_), .Y(mai_mai_n826_));
  OAI210     m0798(.A0(mai_mai_n752_), .A1(mai_mai_n817_), .B0(mai_mai_n782_), .Y(mai_mai_n827_));
  NO2        m0799(.A(mai_mai_n827_), .B(mai_mai_n551_), .Y(mai_mai_n828_));
  AOI210     m0800(.A0(mai_mai_n111_), .A1(mai_mai_n110_), .B0(mai_mai_n240_), .Y(mai_mai_n829_));
  NO2        m0801(.A(mai_mai_n829_), .B(mai_mai_n783_), .Y(mai_mai_n830_));
  AO210      m0802(.A0(mai_mai_n770_), .A1(mai_mai_n759_), .B0(mai_mai_n830_), .Y(mai_mai_n831_));
  NOi31      m0803(.An(mai_mai_n496_), .B(mai_mai_n781_), .C(mai_mai_n273_), .Y(mai_mai_n832_));
  NO4        m0804(.A(mai_mai_n832_), .B(mai_mai_n831_), .C(mai_mai_n828_), .D(mai_mai_n826_), .Y(mai_mai_n833_));
  AN2        m0805(.A(mai_mai_n412_), .B(mai_mai_n677_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n834_), .B(mai_mai_n813_), .Y(mai_mai_n835_));
  NA2        m0807(.A(mai_mai_n763_), .B(mai_mai_n640_), .Y(mai_mai_n836_));
  AN4        m0808(.A(mai_mai_n836_), .B(mai_mai_n835_), .C(mai_mai_n833_), .D(mai_mai_n823_), .Y(mai_mai_n837_));
  NA4        m0809(.A(mai_mai_n837_), .B(mai_mai_n821_), .C(mai_mai_n808_), .D(mai_mai_n756_), .Y(mai12));
  NO4        m0810(.A(mai_mai_n404_), .B(mai_mai_n233_), .C(mai_mai_n533_), .D(mai_mai_n196_), .Y(mai_mai_n839_));
  NO2        m0811(.A(mai_mai_n410_), .B(mai_mai_n109_), .Y(mai_mai_n840_));
  NO2        m0812(.A(mai_mai_n599_), .B(mai_mai_n347_), .Y(mai_mai_n841_));
  INV        m0813(.A(mai_mai_n403_), .Y(mai_mai_n842_));
  AOI210     m0814(.A0(mai_mai_n216_), .A1(mai_mai_n315_), .B0(mai_mai_n182_), .Y(mai_mai_n843_));
  OR2        m0815(.A(mai_mai_n843_), .B(mai_mai_n839_), .Y(mai_mai_n844_));
  NA2        m0816(.A(mai_mai_n844_), .B(mai_mai_n366_), .Y(mai_mai_n845_));
  NO2        m0817(.A(mai_mai_n579_), .B(mai_mai_n243_), .Y(mai_mai_n846_));
  NO2        m0818(.A(mai_mai_n540_), .B(mai_mai_n758_), .Y(mai_mai_n847_));
  NO2        m0819(.A(mai_mai_n139_), .B(mai_mai_n220_), .Y(mai_mai_n848_));
  INV        m0820(.A(mai_mai_n845_), .Y(mai_mai_n849_));
  OR2        m0821(.A(mai_mai_n302_), .B(mai_mai_n840_), .Y(mai_mai_n850_));
  NA2        m0822(.A(mai_mai_n850_), .B(mai_mai_n330_), .Y(mai_mai_n851_));
  NO3        m0823(.A(mai_mai_n123_), .B(mai_mai_n140_), .C(mai_mai_n196_), .Y(mai_mai_n852_));
  NA2        m0824(.A(mai_mai_n852_), .B(mai_mai_n483_), .Y(mai_mai_n853_));
  NA2        m0825(.A(mai_mai_n853_), .B(mai_mai_n851_), .Y(mai_mai_n854_));
  NO3        m0826(.A(mai_mai_n601_), .B(mai_mai_n87_), .C(mai_mai_n45_), .Y(mai_mai_n855_));
  NO4        m0827(.A(mai_mai_n855_), .B(mai_mai_n854_), .C(mai_mai_n849_), .D(mai_mai_n842_), .Y(mai_mai_n856_));
  NA2        m0828(.A(mai_mai_n506_), .B(mai_mai_n134_), .Y(mai_mai_n857_));
  NOi21      m0829(.An(mai_mai_n34_), .B(mai_mai_n593_), .Y(mai_mai_n858_));
  NA2        m0830(.A(mai_mai_n858_), .B(mai_mai_n857_), .Y(mai_mai_n859_));
  OAI210     m0831(.A0(mai_mai_n232_), .A1(mai_mai_n45_), .B0(mai_mai_n859_), .Y(mai_mai_n860_));
  NA2        m0832(.A(mai_mai_n398_), .B(mai_mai_n245_), .Y(mai_mai_n861_));
  NO3        m0833(.A(mai_mai_n740_), .B(mai_mai_n85_), .C(mai_mai_n371_), .Y(mai_mai_n862_));
  NA2        m0834(.A(mai_mai_n861_), .B(mai_mai_n298_), .Y(mai_mai_n863_));
  NO2        m0835(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n864_));
  NO2        m0836(.A(mai_mai_n456_), .B(mai_mai_n277_), .Y(mai_mai_n865_));
  INV        m0837(.A(mai_mai_n865_), .Y(mai_mai_n866_));
  NO2        m0838(.A(mai_mai_n866_), .B(mai_mai_n134_), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n574_), .B(mai_mai_n336_), .Y(mai_mai_n868_));
  INV        m0840(.A(mai_mai_n338_), .Y(mai_mai_n869_));
  NO4        m0841(.A(mai_mai_n869_), .B(mai_mai_n867_), .C(mai_mai_n863_), .D(mai_mai_n860_), .Y(mai_mai_n870_));
  NA2        m0842(.A(mai_mai_n324_), .B(g), .Y(mai_mai_n871_));
  NA2        m0843(.A(mai_mai_n146_), .B(i), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n873_));
  OAI220     m0845(.A0(mai_mai_n873_), .A1(mai_mai_n181_), .B0(mai_mai_n872_), .B1(mai_mai_n87_), .Y(mai_mai_n874_));
  AOI210     m0846(.A0(mai_mai_n381_), .A1(mai_mai_n37_), .B0(mai_mai_n874_), .Y(mai_mai_n875_));
  NO2        m0847(.A(mai_mai_n134_), .B(mai_mai_n80_), .Y(mai_mai_n876_));
  OR2        m0848(.A(mai_mai_n876_), .B(mai_mai_n505_), .Y(mai_mai_n877_));
  NA2        m0849(.A(mai_mai_n506_), .B(mai_mai_n351_), .Y(mai_mai_n878_));
  AOI210     m0850(.A0(mai_mai_n878_), .A1(n), .B0(mai_mai_n877_), .Y(mai_mai_n879_));
  OAI220     m0851(.A0(mai_mai_n879_), .A1(mai_mai_n871_), .B0(mai_mai_n875_), .B1(mai_mai_n311_), .Y(mai_mai_n880_));
  NO2        m0852(.A(mai_mai_n599_), .B(mai_mai_n451_), .Y(mai_mai_n881_));
  NA3        m0853(.A(mai_mai_n320_), .B(mai_mai_n569_), .C(i), .Y(mai_mai_n882_));
  OAI210     m0854(.A0(mai_mai_n401_), .A1(mai_mai_n287_), .B0(mai_mai_n882_), .Y(mai_mai_n883_));
  OAI220     m0855(.A0(mai_mai_n883_), .A1(mai_mai_n881_), .B0(mai_mai_n613_), .B1(mai_mai_n685_), .Y(mai_mai_n884_));
  OR3        m0856(.A(mai_mai_n287_), .B(mai_mai_n397_), .C(f), .Y(mai_mai_n885_));
  NA3        m0857(.A(mai_mai_n569_), .B(mai_mai_n76_), .C(i), .Y(mai_mai_n886_));
  OR2        m0858(.A(mai_mai_n885_), .B(mai_mai_n539_), .Y(mai_mai_n887_));
  NA2        m0859(.A(mai_mai_n627_), .B(mai_mai_n795_), .Y(mai_mai_n888_));
  NA2        m0860(.A(mai_mai_n760_), .B(mai_mai_n402_), .Y(mai_mai_n889_));
  NA2        m0861(.A(mai_mai_n204_), .B(mai_mai_n73_), .Y(mai_mai_n890_));
  NA3        m0862(.A(mai_mai_n890_), .B(mai_mai_n886_), .C(mai_mai_n885_), .Y(mai_mai_n891_));
  AOI220     m0863(.A0(mai_mai_n891_), .A1(mai_mai_n238_), .B0(mai_mai_n889_), .B1(mai_mai_n888_), .Y(mai_mai_n892_));
  NA3        m0864(.A(mai_mai_n892_), .B(mai_mai_n887_), .C(mai_mai_n884_), .Y(mai_mai_n893_));
  NO2        m0865(.A(mai_mai_n347_), .B(mai_mai_n86_), .Y(mai_mai_n894_));
  OAI210     m0866(.A0(mai_mai_n894_), .A1(mai_mai_n846_), .B0(mai_mai_n221_), .Y(mai_mai_n895_));
  NO2        m0867(.A(mai_mai_n416_), .B(mai_mai_n196_), .Y(mai_mai_n896_));
  AOI220     m0868(.A0(mai_mai_n896_), .A1(mai_mai_n352_), .B0(mai_mai_n850_), .B1(mai_mai_n200_), .Y(mai_mai_n897_));
  NA2        m0869(.A(mai_mai_n841_), .B(mai_mai_n848_), .Y(mai_mai_n898_));
  NA3        m0870(.A(mai_mai_n898_), .B(mai_mai_n897_), .C(mai_mai_n895_), .Y(mai_mai_n899_));
  OAI210     m0871(.A0(mai_mai_n889_), .A1(mai_mai_n847_), .B0(mai_mai_n495_), .Y(mai_mai_n900_));
  AOI210     m0872(.A0(mai_mai_n382_), .A1(mai_mai_n375_), .B0(mai_mai_n740_), .Y(mai_mai_n901_));
  INV        m0873(.A(mai_mai_n901_), .Y(mai_mai_n902_));
  NA2        m0874(.A(mai_mai_n584_), .B(mai_mai_n483_), .Y(mai_mai_n903_));
  NA3        m0875(.A(mai_mai_n903_), .B(mai_mai_n902_), .C(mai_mai_n900_), .Y(mai_mai_n904_));
  NO4        m0876(.A(mai_mai_n904_), .B(mai_mai_n899_), .C(mai_mai_n893_), .D(mai_mai_n880_), .Y(mai_mai_n905_));
  NAi31      m0877(.An(mai_mai_n132_), .B(mai_mai_n383_), .C(n), .Y(mai_mai_n906_));
  NO3        m0878(.A(mai_mai_n119_), .B(mai_mai_n318_), .C(mai_mai_n767_), .Y(mai_mai_n907_));
  NO2        m0879(.A(mai_mai_n907_), .B(mai_mai_n906_), .Y(mai_mai_n908_));
  NO3        m0880(.A(mai_mai_n253_), .B(mai_mai_n132_), .C(mai_mai_n371_), .Y(mai_mai_n909_));
  AOI210     m0881(.A0(mai_mai_n909_), .A1(mai_mai_n452_), .B0(mai_mai_n908_), .Y(mai_mai_n910_));
  INV        m0882(.A(mai_mai_n910_), .Y(mai_mai_n911_));
  INV        m0883(.A(mai_mai_n213_), .Y(mai_mai_n912_));
  NAi21      m0884(.An(mai_mai_n506_), .B(mai_mai_n896_), .Y(mai_mai_n913_));
  NO3        m0885(.A(mai_mai_n401_), .B(mai_mai_n287_), .C(mai_mai_n69_), .Y(mai_mai_n914_));
  AOI220     m0886(.A0(mai_mai_n914_), .A1(mai_mai_n399_), .B0(mai_mai_n440_), .B1(g), .Y(mai_mai_n915_));
  NA2        m0887(.A(mai_mai_n915_), .B(mai_mai_n913_), .Y(mai_mai_n916_));
  NO2        m0888(.A(mai_mai_n906_), .B(mai_mai_n216_), .Y(mai_mai_n917_));
  NO3        m0889(.A(n), .B(mai_mai_n137_), .C(mai_mai_n195_), .Y(mai_mai_n918_));
  OAI210     m0890(.A0(mai_mai_n918_), .A1(mai_mai_n477_), .B0(mai_mai_n348_), .Y(mai_mai_n919_));
  OAI220     m0891(.A0(mai_mai_n841_), .A1(mai_mai_n847_), .B0(mai_mai_n496_), .B1(mai_mai_n391_), .Y(mai_mai_n920_));
  NA3        m0892(.A(mai_mai_n920_), .B(mai_mai_n919_), .C(mai_mai_n563_), .Y(mai_mai_n921_));
  OAI210     m0893(.A0(mai_mai_n843_), .A1(mai_mai_n839_), .B0(mai_mai_n912_), .Y(mai_mai_n922_));
  AOI210     m0894(.A0(mai_mai_n350_), .A1(mai_mai_n348_), .B0(mai_mai_n310_), .Y(mai_mai_n923_));
  NA3        m0895(.A(mai_mai_n923_), .B(mai_mai_n922_), .C(mai_mai_n254_), .Y(mai_mai_n924_));
  OR3        m0896(.A(mai_mai_n924_), .B(mai_mai_n921_), .C(mai_mai_n917_), .Y(mai_mai_n925_));
  NO3        m0897(.A(mai_mai_n925_), .B(mai_mai_n916_), .C(mai_mai_n911_), .Y(mai_mai_n926_));
  NA4        m0898(.A(mai_mai_n926_), .B(mai_mai_n905_), .C(mai_mai_n870_), .D(mai_mai_n856_), .Y(mai13));
  AN2        m0899(.A(c), .B(b), .Y(mai_mai_n928_));
  NA3        m0900(.A(mai_mai_n231_), .B(mai_mai_n928_), .C(m), .Y(mai_mai_n929_));
  NA2        m0901(.A(mai_mai_n450_), .B(f), .Y(mai_mai_n930_));
  NO3        m0902(.A(mai_mai_n930_), .B(mai_mai_n929_), .C(mai_mai_n534_), .Y(mai_mai_n931_));
  NAi32      m0903(.An(d), .Bn(c), .C(e), .Y(mai_mai_n932_));
  NA2        m0904(.A(mai_mai_n131_), .B(mai_mai_n45_), .Y(mai_mai_n933_));
  NO4        m0905(.A(mai_mai_n933_), .B(mai_mai_n932_), .C(mai_mai_n540_), .D(mai_mai_n283_), .Y(mai_mai_n934_));
  NA2        m0906(.A(mai_mai_n374_), .B(mai_mai_n195_), .Y(mai_mai_n935_));
  AN2        m0907(.A(d), .B(c), .Y(mai_mai_n936_));
  NA2        m0908(.A(mai_mai_n936_), .B(mai_mai_n109_), .Y(mai_mai_n937_));
  NO4        m0909(.A(mai_mai_n937_), .B(mai_mai_n935_), .C(mai_mai_n158_), .D(mai_mai_n153_), .Y(mai_mai_n938_));
  NA2        m0910(.A(mai_mai_n450_), .B(c), .Y(mai_mai_n939_));
  NO4        m0911(.A(mai_mai_n933_), .B(mai_mai_n536_), .C(mai_mai_n939_), .D(mai_mai_n283_), .Y(mai_mai_n940_));
  OR2        m0912(.A(mai_mai_n938_), .B(mai_mai_n940_), .Y(mai_mai_n941_));
  OR3        m0913(.A(mai_mai_n941_), .B(mai_mai_n934_), .C(mai_mai_n931_), .Y(mai_mai_n942_));
  NAi32      m0914(.An(f), .Bn(e), .C(c), .Y(mai_mai_n943_));
  NO2        m0915(.A(mai_mai_n943_), .B(mai_mai_n135_), .Y(mai_mai_n944_));
  NA2        m0916(.A(mai_mai_n944_), .B(g), .Y(mai_mai_n945_));
  OR2        m0917(.A(mai_mai_n207_), .B(mai_mai_n158_), .Y(mai_mai_n946_));
  NO2        m0918(.A(mai_mai_n946_), .B(mai_mai_n945_), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n939_), .B(mai_mai_n283_), .Y(mai_mai_n948_));
  NA2        m0920(.A(mai_mai_n571_), .B(mai_mai_n1342_), .Y(mai_mai_n949_));
  NOi21      m0921(.An(mai_mai_n948_), .B(mai_mai_n949_), .Y(mai_mai_n950_));
  NO2        m0922(.A(mai_mai_n689_), .B(mai_mai_n105_), .Y(mai_mai_n951_));
  NOi41      m0923(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n952_));
  NA2        m0924(.A(mai_mai_n952_), .B(mai_mai_n951_), .Y(mai_mai_n953_));
  NO2        m0925(.A(mai_mai_n953_), .B(mai_mai_n945_), .Y(mai_mai_n954_));
  NA3        m0926(.A(k), .B(j), .C(i), .Y(mai_mai_n955_));
  NO3        m0927(.A(mai_mai_n955_), .B(mai_mai_n283_), .C(mai_mai_n86_), .Y(mai_mai_n956_));
  BUFFER     m0928(.A(mai_mai_n956_), .Y(mai_mai_n957_));
  OR4        m0929(.A(mai_mai_n957_), .B(mai_mai_n954_), .C(mai_mai_n950_), .D(mai_mai_n947_), .Y(mai_mai_n958_));
  NA3        m0930(.A(mai_mai_n424_), .B(mai_mai_n313_), .C(mai_mai_n54_), .Y(mai_mai_n959_));
  NO2        m0931(.A(mai_mai_n959_), .B(mai_mai_n949_), .Y(mai_mai_n960_));
  NO3        m0932(.A(mai_mai_n959_), .B(mai_mai_n536_), .C(mai_mai_n409_), .Y(mai_mai_n961_));
  NO2        m0933(.A(f), .B(c), .Y(mai_mai_n962_));
  NOi21      m0934(.An(mai_mai_n962_), .B(mai_mai_n404_), .Y(mai_mai_n963_));
  NA2        m0935(.A(mai_mai_n963_), .B(mai_mai_n57_), .Y(mai_mai_n964_));
  NO3        m0936(.A(k), .B(mai_mai_n227_), .C(l), .Y(mai_mai_n965_));
  NOi31      m0937(.An(mai_mai_n965_), .B(mai_mai_n964_), .C(j), .Y(mai_mai_n966_));
  OR3        m0938(.A(mai_mai_n966_), .B(mai_mai_n961_), .C(mai_mai_n960_), .Y(mai_mai_n967_));
  OR3        m0939(.A(mai_mai_n967_), .B(mai_mai_n958_), .C(mai_mai_n942_), .Y(mai02));
  OR2        m0940(.A(l), .B(k), .Y(mai_mai_n969_));
  OR3        m0941(.A(h), .B(g), .C(f), .Y(mai_mai_n970_));
  OR3        m0942(.A(n), .B(m), .C(i), .Y(mai_mai_n971_));
  NO4        m0943(.A(mai_mai_n971_), .B(mai_mai_n970_), .C(mai_mai_n969_), .D(e), .Y(mai_mai_n972_));
  NO2        m0944(.A(mai_mai_n956_), .B(mai_mai_n934_), .Y(mai_mai_n973_));
  AN3        m0945(.A(g), .B(f), .C(c), .Y(mai_mai_n974_));
  NA2        m0946(.A(mai_mai_n974_), .B(mai_mai_n424_), .Y(mai_mai_n975_));
  OR2        m0947(.A(mai_mai_n955_), .B(mai_mai_n283_), .Y(mai_mai_n976_));
  OR2        m0948(.A(mai_mai_n976_), .B(mai_mai_n975_), .Y(mai_mai_n977_));
  NO3        m0949(.A(mai_mai_n959_), .B(mai_mai_n933_), .C(mai_mai_n536_), .Y(mai_mai_n978_));
  NO2        m0950(.A(mai_mai_n978_), .B(mai_mai_n947_), .Y(mai_mai_n979_));
  NA3        m0951(.A(l), .B(k), .C(j), .Y(mai_mai_n980_));
  NA2        m0952(.A(i), .B(h), .Y(mai_mai_n981_));
  NO3        m0953(.A(mai_mai_n981_), .B(mai_mai_n980_), .C(mai_mai_n123_), .Y(mai_mai_n982_));
  NO3        m0954(.A(mai_mai_n133_), .B(mai_mai_n264_), .C(mai_mai_n196_), .Y(mai_mai_n983_));
  AOI210     m0955(.A0(mai_mai_n983_), .A1(mai_mai_n982_), .B0(mai_mai_n950_), .Y(mai_mai_n984_));
  NA3        m0956(.A(c), .B(b), .C(a), .Y(mai_mai_n985_));
  NO3        m0957(.A(mai_mai_n985_), .B(mai_mai_n812_), .C(mai_mai_n195_), .Y(mai_mai_n986_));
  NO2        m0958(.A(mai_mai_n277_), .B(mai_mai_n49_), .Y(mai_mai_n987_));
  AOI210     m0959(.A0(mai_mai_n987_), .A1(mai_mai_n986_), .B0(mai_mai_n960_), .Y(mai_mai_n988_));
  AN4        m0960(.A(mai_mai_n988_), .B(mai_mai_n984_), .C(mai_mai_n979_), .D(mai_mai_n977_), .Y(mai_mai_n989_));
  NO2        m0961(.A(mai_mai_n937_), .B(mai_mai_n935_), .Y(mai_mai_n990_));
  NA2        m0962(.A(mai_mai_n953_), .B(mai_mai_n946_), .Y(mai_mai_n991_));
  AOI210     m0963(.A0(mai_mai_n991_), .A1(mai_mai_n990_), .B0(mai_mai_n931_), .Y(mai_mai_n992_));
  NAi41      m0964(.An(mai_mai_n972_), .B(mai_mai_n992_), .C(mai_mai_n989_), .D(mai_mai_n973_), .Y(mai03));
  NA4        m0965(.A(mai_mai_n526_), .B(m), .C(mai_mai_n105_), .D(mai_mai_n195_), .Y(mai_mai_n994_));
  INV        m0966(.A(mai_mai_n994_), .Y(mai_mai_n995_));
  NO3        m0967(.A(mai_mai_n772_), .B(mai_mai_n761_), .C(mai_mai_n652_), .Y(mai_mai_n996_));
  OAI220     m0968(.A0(mai_mai_n996_), .A1(mai_mai_n627_), .B0(mai_mai_n994_), .B1(mai_mai_n537_), .Y(mai_mai_n997_));
  NOi31      m0969(.An(i), .B(k), .C(j), .Y(mai_mai_n998_));
  NA4        m0970(.A(mai_mai_n998_), .B(e), .C(mai_mai_n320_), .D(mai_mai_n313_), .Y(mai_mai_n999_));
  OAI210     m0971(.A0(mai_mai_n740_), .A1(mai_mai_n384_), .B0(mai_mai_n999_), .Y(mai_mai_n1000_));
  NOi31      m0972(.An(m), .B(n), .C(f), .Y(mai_mai_n1001_));
  NA2        m0973(.A(mai_mai_n1001_), .B(mai_mai_n51_), .Y(mai_mai_n1002_));
  NA2        m0974(.A(c), .B(a), .Y(mai_mai_n1003_));
  OAI220     m0975(.A0(mai_mai_n1003_), .A1(mai_mai_n1002_), .B0(mai_mai_n803_), .B1(mai_mai_n390_), .Y(mai_mai_n1004_));
  NA2        m0976(.A(mai_mai_n459_), .B(l), .Y(mai_mai_n1005_));
  NOi31      m0977(.An(mai_mai_n782_), .B(mai_mai_n929_), .C(mai_mai_n1005_), .Y(mai_mai_n1006_));
  NO4        m0978(.A(mai_mai_n1006_), .B(mai_mai_n1004_), .C(mai_mai_n1000_), .D(mai_mai_n901_), .Y(mai_mai_n1007_));
  INV        m0979(.A(mai_mai_n264_), .Y(mai_mai_n1008_));
  INV        m0980(.A(mai_mai_n934_), .Y(mai_mai_n1009_));
  NO2        m0981(.A(mai_mai_n981_), .B(mai_mai_n442_), .Y(mai_mai_n1010_));
  NO2        m0982(.A(mai_mai_n83_), .B(g), .Y(mai_mai_n1011_));
  AOI210     m0983(.A0(mai_mai_n1011_), .A1(mai_mai_n1010_), .B0(mai_mai_n965_), .Y(mai_mai_n1012_));
  OR2        m0984(.A(mai_mai_n1012_), .B(mai_mai_n964_), .Y(mai_mai_n1013_));
  NA3        m0985(.A(mai_mai_n1013_), .B(mai_mai_n1009_), .C(mai_mai_n1007_), .Y(mai_mai_n1014_));
  NO4        m0986(.A(mai_mai_n1014_), .B(mai_mai_n997_), .C(mai_mai_n741_), .D(mai_mai_n518_), .Y(mai_mai_n1015_));
  NA2        m0987(.A(c), .B(b), .Y(mai_mai_n1016_));
  NO2        m0988(.A(mai_mai_n639_), .B(mai_mai_n1016_), .Y(mai_mai_n1017_));
  OAI210     m0989(.A0(mai_mai_n781_), .A1(mai_mai_n754_), .B0(mai_mai_n377_), .Y(mai_mai_n1018_));
  NA2        m0990(.A(mai_mai_n1018_), .B(mai_mai_n1017_), .Y(mai_mai_n1019_));
  NAi21      m0991(.An(mai_mai_n385_), .B(mai_mai_n1017_), .Y(mai_mai_n1020_));
  OAI210     m0992(.A0(mai_mai_n500_), .A1(mai_mai_n39_), .B0(mai_mai_n1008_), .Y(mai_mai_n1021_));
  NA2        m0993(.A(mai_mai_n1021_), .B(mai_mai_n1020_), .Y(mai_mai_n1022_));
  NA2        m0994(.A(mai_mai_n267_), .B(g), .Y(mai_mai_n1023_));
  NAi21      m0995(.An(f), .B(d), .Y(mai_mai_n1024_));
  NO2        m0996(.A(mai_mai_n1024_), .B(mai_mai_n985_), .Y(mai_mai_n1025_));
  INV        m0997(.A(mai_mai_n1025_), .Y(mai_mai_n1026_));
  NO2        m0998(.A(mai_mai_n1023_), .B(mai_mai_n1026_), .Y(mai_mai_n1027_));
  AOI210     m0999(.A0(mai_mai_n1027_), .A1(mai_mai_n106_), .B0(mai_mai_n1022_), .Y(mai_mai_n1028_));
  INV        m1000(.A(mai_mai_n426_), .Y(mai_mai_n1029_));
  NO2        m1001(.A(mai_mai_n162_), .B(mai_mai_n220_), .Y(mai_mai_n1030_));
  NA2        m1002(.A(mai_mai_n1030_), .B(m), .Y(mai_mai_n1031_));
  NA3        m1003(.A(mai_mai_n829_), .B(mai_mai_n1005_), .C(mai_mai_n429_), .Y(mai_mai_n1032_));
  OAI210     m1004(.A0(mai_mai_n1032_), .A1(mai_mai_n288_), .B0(mai_mai_n427_), .Y(mai_mai_n1033_));
  AOI210     m1005(.A0(mai_mai_n1033_), .A1(mai_mai_n1029_), .B0(mai_mai_n1031_), .Y(mai_mai_n1034_));
  NA2        m1006(.A(mai_mai_n143_), .B(mai_mai_n33_), .Y(mai_mai_n1035_));
  AOI210     m1007(.A0(mai_mai_n868_), .A1(mai_mai_n1035_), .B0(mai_mai_n196_), .Y(mai_mai_n1036_));
  OAI210     m1008(.A0(mai_mai_n1036_), .A1(mai_mai_n406_), .B0(mai_mai_n1025_), .Y(mai_mai_n1037_));
  NO2        m1009(.A(mai_mai_n341_), .B(mai_mai_n340_), .Y(mai_mai_n1038_));
  AOI210     m1010(.A0(mai_mai_n1030_), .A1(mai_mai_n393_), .B0(mai_mai_n862_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n1039_), .B(mai_mai_n1037_), .Y(mai_mai_n1040_));
  NO2        m1012(.A(mai_mai_n1040_), .B(mai_mai_n1034_), .Y(mai_mai_n1041_));
  NA4        m1013(.A(mai_mai_n1041_), .B(mai_mai_n1028_), .C(mai_mai_n1019_), .D(mai_mai_n1015_), .Y(mai00));
  NO2        m1014(.A(mai_mai_n276_), .B(mai_mai_n257_), .Y(mai_mai_n1043_));
  NO2        m1015(.A(mai_mai_n1043_), .B(mai_mai_n529_), .Y(mai_mai_n1044_));
  AOI210     m1016(.A0(mai_mai_n809_), .A1(mai_mai_n848_), .B0(mai_mai_n1000_), .Y(mai_mai_n1045_));
  NO3        m1017(.A(mai_mai_n978_), .B(mai_mai_n862_), .C(mai_mai_n650_), .Y(mai_mai_n1046_));
  NA3        m1018(.A(mai_mai_n1046_), .B(mai_mai_n1045_), .C(mai_mai_n902_), .Y(mai_mai_n1047_));
  NA2        m1019(.A(mai_mai_n461_), .B(f), .Y(mai_mai_n1048_));
  OAI210     m1020(.A0(mai_mai_n907_), .A1(mai_mai_n40_), .B0(mai_mai_n586_), .Y(mai_mai_n1049_));
  NA3        m1021(.A(mai_mai_n1049_), .B(mai_mai_n237_), .C(n), .Y(mai_mai_n1050_));
  AOI210     m1022(.A0(mai_mai_n1050_), .A1(mai_mai_n1048_), .B0(mai_mai_n937_), .Y(mai_mai_n1051_));
  NO4        m1023(.A(mai_mai_n1051_), .B(mai_mai_n1047_), .C(mai_mai_n1044_), .D(mai_mai_n958_), .Y(mai_mai_n1052_));
  NA3        m1024(.A(mai_mai_n152_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1053_));
  NA3        m1025(.A(d), .B(mai_mai_n54_), .C(b), .Y(mai_mai_n1054_));
  NOi31      m1026(.An(n), .B(m), .C(i), .Y(mai_mai_n1055_));
  NA3        m1027(.A(mai_mai_n1055_), .B(mai_mai_n589_), .C(mai_mai_n51_), .Y(mai_mai_n1056_));
  OAI210     m1028(.A0(mai_mai_n1054_), .A1(mai_mai_n1053_), .B0(mai_mai_n1056_), .Y(mai_mai_n1057_));
  INV        m1029(.A(mai_mai_n528_), .Y(mai_mai_n1058_));
  NO4        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1057_), .C(mai_mai_n1038_), .D(mai_mai_n832_), .Y(mai_mai_n1059_));
  NA3        m1031(.A(mai_mai_n353_), .B(mai_mai_n203_), .C(g), .Y(mai_mai_n1060_));
  OR2        m1032(.A(mai_mai_n354_), .B(mai_mai_n126_), .Y(mai_mai_n1061_));
  NO2        m1033(.A(h), .B(g), .Y(mai_mai_n1062_));
  NA4        m1034(.A(mai_mai_n452_), .B(mai_mai_n424_), .C(mai_mai_n1062_), .D(mai_mai_n928_), .Y(mai_mai_n1063_));
  NA2        m1035(.A(mai_mai_n852_), .B(mai_mai_n527_), .Y(mai_mai_n1064_));
  NA3        m1036(.A(mai_mai_n1064_), .B(mai_mai_n1063_), .C(mai_mai_n1061_), .Y(mai_mai_n1065_));
  NO2        m1037(.A(mai_mai_n1065_), .B(mai_mai_n247_), .Y(mai_mai_n1066_));
  NO2        m1038(.A(mai_mai_n222_), .B(mai_mai_n161_), .Y(mai_mai_n1067_));
  NA2        m1039(.A(mai_mai_n1067_), .B(mai_mai_n391_), .Y(mai_mai_n1068_));
  NA3        m1040(.A(mai_mai_n159_), .B(mai_mai_n105_), .C(g), .Y(mai_mai_n1069_));
  NOi31      m1041(.An(mai_mai_n788_), .B(mai_mai_n1345_), .C(mai_mai_n1069_), .Y(mai_mai_n1070_));
  NAi31      m1042(.An(mai_mai_n166_), .B(mai_mai_n778_), .C(mai_mai_n424_), .Y(mai_mai_n1071_));
  NAi31      m1043(.An(mai_mai_n1070_), .B(mai_mai_n1071_), .C(mai_mai_n1068_), .Y(mai_mai_n1072_));
  NO2        m1044(.A(mai_mai_n256_), .B(mai_mai_n69_), .Y(mai_mai_n1073_));
  NO3        m1045(.A(mai_mai_n390_), .B(mai_mai_n751_), .C(n), .Y(mai_mai_n1074_));
  AOI210     m1046(.A0(mai_mai_n1074_), .A1(mai_mai_n1073_), .B0(mai_mai_n972_), .Y(mai_mai_n1075_));
  NAi31      m1047(.An(mai_mai_n940_), .B(mai_mai_n1075_), .C(mai_mai_n68_), .Y(mai_mai_n1076_));
  NO4        m1048(.A(mai_mai_n1076_), .B(mai_mai_n1072_), .C(mai_mai_n300_), .D(mai_mai_n470_), .Y(mai_mai_n1077_));
  AN3        m1049(.A(mai_mai_n1077_), .B(mai_mai_n1066_), .C(mai_mai_n1059_), .Y(mai_mai_n1078_));
  NA2        m1050(.A(mai_mai_n514_), .B(mai_mai_n225_), .Y(mai_mai_n1079_));
  NA2        m1051(.A(mai_mai_n995_), .B(mai_mai_n488_), .Y(mai_mai_n1080_));
  INV        m1052(.A(mai_mai_n1080_), .Y(mai_mai_n1081_));
  OAI210     m1053(.A0(mai_mai_n422_), .A1(mai_mai_n113_), .B0(mai_mai_n783_), .Y(mai_mai_n1082_));
  NA2        m1054(.A(mai_mai_n1082_), .B(mai_mai_n1032_), .Y(mai_mai_n1083_));
  OR3        m1055(.A(mai_mai_n937_), .B(mai_mai_n253_), .C(mai_mai_n205_), .Y(mai_mai_n1084_));
  NO2        m1056(.A(mai_mai_n199_), .B(mai_mai_n196_), .Y(mai_mai_n1085_));
  NA2        m1057(.A(n), .B(e), .Y(mai_mai_n1086_));
  NO2        m1058(.A(mai_mai_n1086_), .B(mai_mai_n135_), .Y(mai_mai_n1087_));
  AOI220     m1059(.A0(mai_mai_n1087_), .A1(mai_mai_n255_), .B0(mai_mai_n765_), .B1(mai_mai_n1085_), .Y(mai_mai_n1088_));
  OAI210     m1060(.A0(mai_mai_n333_), .A1(mai_mai_n289_), .B0(mai_mai_n408_), .Y(mai_mai_n1089_));
  NA4        m1061(.A(mai_mai_n1089_), .B(mai_mai_n1088_), .C(mai_mai_n1084_), .D(mai_mai_n1083_), .Y(mai_mai_n1090_));
  AOI210     m1062(.A0(mai_mai_n1087_), .A1(mai_mai_n769_), .B0(mai_mai_n741_), .Y(mai_mai_n1091_));
  AOI220     m1063(.A0(mai_mai_n858_), .A1(mai_mai_n527_), .B0(mai_mai_n589_), .B1(mai_mai_n228_), .Y(mai_mai_n1092_));
  NO2        m1064(.A(mai_mai_n63_), .B(h), .Y(mai_mai_n1093_));
  NO3        m1065(.A(mai_mai_n937_), .B(mai_mai_n935_), .C(mai_mai_n662_), .Y(mai_mai_n1094_));
  NO2        m1066(.A(mai_mai_n969_), .B(mai_mai_n123_), .Y(mai_mai_n1095_));
  AN2        m1067(.A(mai_mai_n1095_), .B(mai_mai_n983_), .Y(mai_mai_n1096_));
  OAI210     m1068(.A0(mai_mai_n1096_), .A1(mai_mai_n1094_), .B0(mai_mai_n1093_), .Y(mai_mai_n1097_));
  NA3        m1069(.A(mai_mai_n1097_), .B(mai_mai_n1092_), .C(mai_mai_n1091_), .Y(mai_mai_n1098_));
  NO4        m1070(.A(mai_mai_n1098_), .B(mai_mai_n1090_), .C(mai_mai_n1081_), .D(mai_mai_n1079_), .Y(mai_mai_n1099_));
  NA2        m1071(.A(mai_mai_n755_), .B(mai_mai_n684_), .Y(mai_mai_n1100_));
  NA4        m1072(.A(mai_mai_n1100_), .B(mai_mai_n1099_), .C(mai_mai_n1078_), .D(mai_mai_n1052_), .Y(mai01));
  NO3        m1073(.A(mai_mai_n725_), .B(mai_mai_n717_), .C(mai_mai_n437_), .Y(mai_mai_n1102_));
  NA2        m1074(.A(mai_mai_n1102_), .B(mai_mai_n919_), .Y(mai_mai_n1103_));
  NA2        m1075(.A(mai_mai_n506_), .B(mai_mai_n252_), .Y(mai_mai_n1104_));
  NA2        m1076(.A(mai_mai_n865_), .B(mai_mai_n1104_), .Y(mai_mai_n1105_));
  NA3        m1077(.A(mai_mai_n1105_), .B(mai_mai_n825_), .C(mai_mai_n312_), .Y(mai_mai_n1106_));
  NA2        m1078(.A(mai_mai_n645_), .B(mai_mai_n91_), .Y(mai_mai_n1107_));
  NO2        m1079(.A(mai_mai_n1107_), .B(i), .Y(mai_mai_n1108_));
  NA2        m1080(.A(mai_mai_n1108_), .B(mai_mai_n576_), .Y(mai_mai_n1109_));
  INV        m1081(.A(mai_mai_n1109_), .Y(mai_mai_n1110_));
  NO2        m1082(.A(mai_mai_n612_), .B(mai_mai_n464_), .Y(mai_mai_n1111_));
  OR2        m1083(.A(mai_mai_n176_), .B(mai_mai_n174_), .Y(mai_mai_n1112_));
  NA3        m1084(.A(mai_mai_n1112_), .B(mai_mai_n1111_), .C(mai_mai_n129_), .Y(mai_mai_n1113_));
  NO4        m1085(.A(mai_mai_n1113_), .B(mai_mai_n1110_), .C(mai_mai_n1106_), .D(mai_mai_n1103_), .Y(mai_mai_n1114_));
  NA2        m1086(.A(mai_mai_n1060_), .B(mai_mai_n188_), .Y(mai_mai_n1115_));
  OAI210     m1087(.A0(mai_mai_n1115_), .A1(mai_mai_n279_), .B0(mai_mai_n483_), .Y(mai_mai_n1116_));
  NA2        m1088(.A(mai_mai_n491_), .B(mai_mai_n362_), .Y(mai_mai_n1117_));
  NA2        m1089(.A(mai_mai_n515_), .B(mai_mai_n1117_), .Y(mai_mai_n1118_));
  AOI210     m1090(.A0(mai_mai_n185_), .A1(mai_mai_n85_), .B0(mai_mai_n195_), .Y(mai_mai_n1119_));
  OAI210     m1091(.A0(mai_mai_n731_), .A1(mai_mai_n391_), .B0(mai_mai_n1119_), .Y(mai_mai_n1120_));
  AN2        m1092(.A(m), .B(k), .Y(mai_mai_n1121_));
  NA2        m1093(.A(mai_mai_n34_), .B(mai_mai_n1121_), .Y(mai_mai_n1122_));
  OR2        m1094(.A(mai_mai_n1122_), .B(mai_mai_n311_), .Y(mai_mai_n1123_));
  NA4        m1095(.A(mai_mai_n1123_), .B(mai_mai_n1120_), .C(mai_mai_n1118_), .D(mai_mai_n1116_), .Y(mai_mai_n1124_));
  AOI210     m1096(.A0(mai_mai_n543_), .A1(mai_mai_n111_), .B0(mai_mai_n547_), .Y(mai_mai_n1125_));
  INV        m1097(.A(mai_mai_n1125_), .Y(mai_mai_n1126_));
  NA2        m1098(.A(mai_mai_n262_), .B(mai_mai_n176_), .Y(mai_mai_n1127_));
  NA2        m1099(.A(mai_mai_n1127_), .B(mai_mai_n602_), .Y(mai_mai_n1128_));
  NO3        m1100(.A(mai_mai_n740_), .B(mai_mai_n185_), .C(mai_mai_n371_), .Y(mai_mai_n1129_));
  NO2        m1101(.A(mai_mai_n1129_), .B(mai_mai_n862_), .Y(mai_mai_n1130_));
  OAI210     m1102(.A0(mai_mai_n1108_), .A1(mai_mai_n305_), .B0(mai_mai_n613_), .Y(mai_mai_n1131_));
  NA4        m1103(.A(mai_mai_n1131_), .B(mai_mai_n1130_), .C(mai_mai_n1128_), .D(mai_mai_n709_), .Y(mai_mai_n1132_));
  NO3        m1104(.A(mai_mai_n1132_), .B(mai_mai_n1126_), .C(mai_mai_n1124_), .Y(mai_mai_n1133_));
  NA2        m1105(.A(mai_mai_n457_), .B(mai_mai_n56_), .Y(mai_mai_n1134_));
  INV        m1106(.A(mai_mai_n1057_), .Y(mai_mai_n1135_));
  NA3        m1107(.A(mai_mai_n1135_), .B(mai_mai_n1134_), .C(mai_mai_n683_), .Y(mai_mai_n1136_));
  NO2        m1108(.A(mai_mai_n872_), .B(mai_mai_n215_), .Y(mai_mai_n1137_));
  NO2        m1109(.A(mai_mai_n873_), .B(mai_mai_n508_), .Y(mai_mai_n1138_));
  OAI210     m1110(.A0(mai_mai_n1138_), .A1(mai_mai_n1137_), .B0(mai_mai_n318_), .Y(mai_mai_n1139_));
  NO3        m1111(.A(mai_mai_n75_), .B(mai_mai_n277_), .C(mai_mai_n45_), .Y(mai_mai_n1140_));
  NA2        m1112(.A(mai_mai_n1140_), .B(mai_mai_n505_), .Y(mai_mai_n1141_));
  NA2        m1113(.A(mai_mai_n1141_), .B(mai_mai_n608_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n1140_), .B(mai_mai_n734_), .Y(mai_mai_n1143_));
  NA2        m1115(.A(mai_mai_n1143_), .B(mai_mai_n356_), .Y(mai_mai_n1144_));
  NOi41      m1116(.An(mai_mai_n1139_), .B(mai_mai_n1144_), .C(mai_mai_n1142_), .D(mai_mai_n1136_), .Y(mai_mai_n1145_));
  NO2        m1117(.A(mai_mai_n122_), .B(mai_mai_n45_), .Y(mai_mai_n1146_));
  NO2        m1118(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1147_));
  AO220      m1119(.A0(mai_mai_n1147_), .A1(mai_mai_n566_), .B0(mai_mai_n1146_), .B1(mai_mai_n643_), .Y(mai_mai_n1148_));
  NA2        m1120(.A(mai_mai_n1148_), .B(mai_mai_n318_), .Y(mai_mai_n1149_));
  NA2        m1121(.A(mai_mai_n1140_), .B(mai_mai_n876_), .Y(mai_mai_n1150_));
  NA2        m1122(.A(mai_mai_n1150_), .B(mai_mai_n1149_), .Y(mai_mai_n1151_));
  NO2        m1123(.A(mai_mai_n559_), .B(mai_mai_n558_), .Y(mai_mai_n1152_));
  NO2        m1124(.A(mai_mai_n1151_), .B(mai_mai_n578_), .Y(mai_mai_n1153_));
  NA4        m1125(.A(mai_mai_n1153_), .B(mai_mai_n1145_), .C(mai_mai_n1133_), .D(mai_mai_n1114_), .Y(mai06));
  OR2        m1126(.A(mai_mai_n1344_), .B(mai_mai_n803_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n1155_), .B(mai_mai_n1139_), .Y(mai_mai_n1156_));
  NO3        m1128(.A(mai_mai_n1156_), .B(mai_mai_n1142_), .C(mai_mai_n236_), .Y(mai_mai_n1157_));
  NO2        m1129(.A(mai_mai_n277_), .B(mai_mai_n45_), .Y(mai_mai_n1158_));
  AOI210     m1130(.A0(mai_mai_n1158_), .A1(mai_mai_n877_), .B0(mai_mai_n1137_), .Y(mai_mai_n1159_));
  AOI210     m1131(.A0(mai_mai_n1158_), .A1(mai_mai_n509_), .B0(mai_mai_n1148_), .Y(mai_mai_n1160_));
  AOI210     m1132(.A0(mai_mai_n1160_), .A1(mai_mai_n1159_), .B0(mai_mai_n315_), .Y(mai_mai_n1161_));
  OAI210     m1133(.A0(mai_mai_n85_), .A1(mai_mai_n40_), .B0(mai_mai_n611_), .Y(mai_mai_n1162_));
  NA2        m1134(.A(mai_mai_n1162_), .B(mai_mai_n582_), .Y(mai_mai_n1163_));
  OAI210     m1135(.A0(mai_mai_n417_), .A1(mai_mai_n230_), .B0(mai_mai_n819_), .Y(mai_mai_n1164_));
  NO2        m1136(.A(mai_mai_n1164_), .B(mai_mai_n128_), .Y(mai_mai_n1165_));
  OR2        m1137(.A(mai_mai_n546_), .B(mai_mai_n545_), .Y(mai_mai_n1166_));
  INV        m1138(.A(mai_mai_n1166_), .Y(mai_mai_n1167_));
  NA3        m1139(.A(mai_mai_n1167_), .B(mai_mai_n1165_), .C(mai_mai_n1163_), .Y(mai_mai_n1168_));
  NO2        m1140(.A(mai_mai_n678_), .B(mai_mai_n339_), .Y(mai_mai_n1169_));
  NO2        m1141(.A(mai_mai_n613_), .B(mai_mai_n685_), .Y(mai_mai_n1170_));
  NOi21      m1142(.An(mai_mai_n1169_), .B(mai_mai_n1170_), .Y(mai_mai_n1171_));
  AN2        m1143(.A(mai_mai_n858_), .B(mai_mai_n585_), .Y(mai_mai_n1172_));
  NO4        m1144(.A(mai_mai_n1172_), .B(mai_mai_n1171_), .C(mai_mai_n1168_), .D(mai_mai_n1161_), .Y(mai_mai_n1173_));
  NO2        m1145(.A(mai_mai_n724_), .B(mai_mai_n258_), .Y(mai_mai_n1174_));
  OAI220     m1146(.A0(mai_mai_n669_), .A1(mai_mai_n47_), .B0(mai_mai_n207_), .B1(mai_mai_n560_), .Y(mai_mai_n1175_));
  OAI210     m1147(.A0(mai_mai_n258_), .A1(c), .B0(mai_mai_n581_), .Y(mai_mai_n1176_));
  AOI220     m1148(.A0(mai_mai_n1176_), .A1(mai_mai_n1175_), .B0(mai_mai_n1174_), .B1(mai_mai_n248_), .Y(mai_mai_n1177_));
  NO3        m1149(.A(mai_mai_n227_), .B(mai_mai_n96_), .C(mai_mai_n264_), .Y(mai_mai_n1178_));
  OAI220     m1150(.A0(mai_mai_n636_), .A1(mai_mai_n230_), .B0(mai_mai_n463_), .B1(mai_mai_n467_), .Y(mai_mai_n1179_));
  NO3        m1151(.A(mai_mai_n1179_), .B(mai_mai_n1178_), .C(mai_mai_n1004_), .Y(mai_mai_n1180_));
  NA3        m1152(.A(mai_mai_n715_), .B(mai_mai_n714_), .C(mai_mai_n400_), .Y(mai_mai_n1181_));
  NAi31      m1153(.An(mai_mai_n678_), .B(mai_mai_n1181_), .C(mai_mai_n184_), .Y(mai_mai_n1182_));
  NA4        m1154(.A(mai_mai_n1182_), .B(mai_mai_n1180_), .C(mai_mai_n1177_), .D(mai_mai_n1092_), .Y(mai_mai_n1183_));
  OR2        m1155(.A(mai_mai_n706_), .B(mai_mai_n493_), .Y(mai_mai_n1184_));
  OR3        m1156(.A(mai_mai_n340_), .B(mai_mai_n207_), .C(mai_mai_n560_), .Y(mai_mai_n1185_));
  NA2        m1157(.A(mai_mai_n522_), .B(mai_mai_n408_), .Y(mai_mai_n1186_));
  NA3        m1158(.A(mai_mai_n1186_), .B(mai_mai_n1185_), .C(mai_mai_n1184_), .Y(mai_mai_n1187_));
  NA2        m1159(.A(mai_mai_n1169_), .B(mai_mai_n684_), .Y(mai_mai_n1188_));
  NO2        m1160(.A(mai_mai_n793_), .B(mai_mai_n440_), .Y(mai_mai_n1189_));
  NA3        m1161(.A(mai_mai_n1189_), .B(mai_mai_n1188_), .C(mai_mai_n1143_), .Y(mai_mai_n1190_));
  NAi21      m1162(.An(j), .B(i), .Y(mai_mai_n1191_));
  NO4        m1163(.A(mai_mai_n1152_), .B(mai_mai_n1191_), .C(mai_mai_n404_), .D(mai_mai_n218_), .Y(mai_mai_n1192_));
  NO4        m1164(.A(mai_mai_n1192_), .B(mai_mai_n1190_), .C(mai_mai_n1187_), .D(mai_mai_n1183_), .Y(mai_mai_n1193_));
  NA4        m1165(.A(mai_mai_n1193_), .B(mai_mai_n1173_), .C(mai_mai_n1157_), .D(mai_mai_n1153_), .Y(mai07));
  NOi21      m1166(.An(j), .B(k), .Y(mai_mai_n1195_));
  NA4        m1167(.A(mai_mai_n159_), .B(mai_mai_n101_), .C(mai_mai_n1195_), .D(f), .Y(mai_mai_n1196_));
  NAi32      m1168(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1197_));
  NO3        m1169(.A(mai_mai_n1197_), .B(g), .C(f), .Y(mai_mai_n1198_));
  OAI210     m1170(.A0(mai_mai_n299_), .A1(mai_mai_n441_), .B0(mai_mai_n1198_), .Y(mai_mai_n1199_));
  NAi21      m1171(.An(f), .B(c), .Y(mai_mai_n1200_));
  OR2        m1172(.A(e), .B(d), .Y(mai_mai_n1201_));
  OAI220     m1173(.A0(mai_mai_n1201_), .A1(mai_mai_n1200_), .B0(mai_mai_n570_), .B1(mai_mai_n301_), .Y(mai_mai_n1202_));
  NA3        m1174(.A(mai_mai_n1202_), .B(mai_mai_n1342_), .C(mai_mai_n159_), .Y(mai_mai_n1203_));
  NOi31      m1175(.An(n), .B(m), .C(b), .Y(mai_mai_n1204_));
  NO3        m1176(.A(mai_mai_n123_), .B(mai_mai_n409_), .C(h), .Y(mai_mai_n1205_));
  NA3        m1177(.A(mai_mai_n1203_), .B(mai_mai_n1199_), .C(mai_mai_n1196_), .Y(mai_mai_n1206_));
  NA2        m1178(.A(mai_mai_n83_), .B(mai_mai_n45_), .Y(mai_mai_n1207_));
  NO2        m1179(.A(mai_mai_n943_), .B(mai_mai_n404_), .Y(mai_mai_n1208_));
  NA3        m1180(.A(mai_mai_n1208_), .B(mai_mai_n1207_), .C(mai_mai_n196_), .Y(mai_mai_n1209_));
  NA2        m1181(.A(mai_mai_n494_), .B(mai_mai_n76_), .Y(mai_mai_n1210_));
  NA2        m1182(.A(mai_mai_n1093_), .B(mai_mai_n271_), .Y(mai_mai_n1211_));
  NA3        m1183(.A(mai_mai_n1211_), .B(mai_mai_n1210_), .C(mai_mai_n1209_), .Y(mai_mai_n1212_));
  NO2        m1184(.A(mai_mai_n1212_), .B(mai_mai_n1206_), .Y(mai_mai_n1213_));
  NO3        m1185(.A(e), .B(d), .C(c), .Y(mai_mai_n1214_));
  NA2        m1186(.A(mai_mai_n1339_), .B(mai_mai_n1214_), .Y(mai_mai_n1215_));
  NO2        m1187(.A(mai_mai_n1215_), .B(mai_mai_n196_), .Y(mai_mai_n1216_));
  NA3        m1188(.A(mai_mai_n633_), .B(mai_mai_n1343_), .C(mai_mai_n105_), .Y(mai_mai_n1217_));
  NO2        m1189(.A(mai_mai_n1217_), .B(mai_mai_n45_), .Y(mai_mai_n1218_));
  NO2        m1190(.A(l), .B(k), .Y(mai_mai_n1219_));
  NOi41      m1191(.An(mai_mai_n498_), .B(mai_mai_n1219_), .C(mai_mai_n435_), .D(mai_mai_n404_), .Y(mai_mai_n1220_));
  NO3        m1192(.A(mai_mai_n404_), .B(d), .C(c), .Y(mai_mai_n1221_));
  NO3        m1193(.A(mai_mai_n1220_), .B(mai_mai_n1218_), .C(mai_mai_n1216_), .Y(mai_mai_n1222_));
  NO2        m1194(.A(k), .B(l), .Y(mai_mai_n1223_));
  NO2        m1195(.A(g), .B(c), .Y(mai_mai_n1224_));
  NA3        m1196(.A(mai_mai_n1224_), .B(mai_mai_n133_), .C(mai_mai_n167_), .Y(mai_mai_n1225_));
  NO2        m1197(.A(mai_mai_n1225_), .B(mai_mai_n1223_), .Y(mai_mai_n1226_));
  NA2        m1198(.A(mai_mai_n1226_), .B(mai_mai_n159_), .Y(mai_mai_n1227_));
  NO2        m1199(.A(mai_mai_n410_), .B(a), .Y(mai_mai_n1228_));
  NA3        m1200(.A(mai_mai_n1228_), .B(mai_mai_n1341_), .C(mai_mai_n106_), .Y(mai_mai_n1229_));
  NO2        m1201(.A(i), .B(h), .Y(mai_mai_n1230_));
  NA2        m1202(.A(mai_mai_n1230_), .B(mai_mai_n203_), .Y(mai_mai_n1231_));
  NA2        m1203(.A(mai_mai_n1024_), .B(h), .Y(mai_mai_n1232_));
  NA2        m1204(.A(mai_mai_n130_), .B(mai_mai_n203_), .Y(mai_mai_n1233_));
  AOI210     m1205(.A0(mai_mai_n237_), .A1(mai_mai_n109_), .B0(mai_mai_n483_), .Y(mai_mai_n1234_));
  OAI220     m1206(.A0(mai_mai_n1234_), .A1(mai_mai_n1231_), .B0(mai_mai_n1233_), .B1(mai_mai_n1232_), .Y(mai_mai_n1235_));
  NO2        m1207(.A(mai_mai_n681_), .B(mai_mai_n168_), .Y(mai_mai_n1236_));
  NOi31      m1208(.An(m), .B(n), .C(b), .Y(mai_mai_n1237_));
  NOi31      m1209(.An(f), .B(d), .C(c), .Y(mai_mai_n1238_));
  NA2        m1210(.A(mai_mai_n1238_), .B(mai_mai_n1237_), .Y(mai_mai_n1239_));
  INV        m1211(.A(mai_mai_n1239_), .Y(mai_mai_n1240_));
  NO3        m1212(.A(mai_mai_n1240_), .B(mai_mai_n1236_), .C(mai_mai_n1235_), .Y(mai_mai_n1241_));
  NA2        m1213(.A(mai_mai_n974_), .B(mai_mai_n424_), .Y(mai_mai_n1242_));
  NO4        m1214(.A(mai_mai_n1242_), .B(mai_mai_n951_), .C(mai_mai_n404_), .D(mai_mai_n45_), .Y(mai_mai_n1243_));
  OAI210     m1215(.A0(mai_mai_n162_), .A1(mai_mai_n478_), .B0(mai_mai_n952_), .Y(mai_mai_n1244_));
  INV        m1216(.A(mai_mai_n1244_), .Y(mai_mai_n1245_));
  NO2        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1243_), .Y(mai_mai_n1246_));
  AN4        m1218(.A(mai_mai_n1246_), .B(mai_mai_n1241_), .C(mai_mai_n1229_), .D(mai_mai_n1227_), .Y(mai_mai_n1247_));
  NA2        m1219(.A(mai_mai_n1204_), .B(mai_mai_n349_), .Y(mai_mai_n1248_));
  NA2        m1220(.A(mai_mai_n982_), .B(mai_mai_n1242_), .Y(mai_mai_n1249_));
  NO4        m1221(.A(mai_mai_n123_), .B(g), .C(f), .D(e), .Y(mai_mai_n1250_));
  NA2        m1222(.A(mai_mai_n272_), .B(h), .Y(mai_mai_n1251_));
  OR2        m1223(.A(e), .B(a), .Y(mai_mai_n1252_));
  OR3        m1224(.A(mai_mai_n493_), .B(mai_mai_n492_), .C(mai_mai_n105_), .Y(mai_mai_n1253_));
  NA2        m1225(.A(mai_mai_n1001_), .B(mai_mai_n371_), .Y(mai_mai_n1254_));
  NA4        m1226(.A(mai_mai_n1249_), .B(mai_mai_n1247_), .C(mai_mai_n1222_), .D(mai_mai_n1213_), .Y(mai_mai_n1255_));
  NAi31      m1227(.An(mai_mai_n1230_), .B(mai_mai_n963_), .C(mai_mai_n153_), .Y(mai_mai_n1256_));
  INV        m1228(.A(mai_mai_n1256_), .Y(mai_mai_n1257_));
  NO3        m1229(.A(mai_mai_n678_), .B(mai_mai_n157_), .C(mai_mai_n374_), .Y(mai_mai_n1258_));
  NO2        m1230(.A(mai_mai_n1258_), .B(mai_mai_n1257_), .Y(mai_mai_n1259_));
  OR2        m1231(.A(n), .B(i), .Y(mai_mai_n1260_));
  OAI210     m1232(.A0(mai_mai_n1260_), .A1(mai_mai_n962_), .B0(mai_mai_n49_), .Y(mai_mai_n1261_));
  AOI220     m1233(.A0(mai_mai_n1261_), .A1(mai_mai_n1062_), .B0(mai_mai_n744_), .B1(mai_mai_n175_), .Y(mai_mai_n1262_));
  INV        m1234(.A(mai_mai_n1262_), .Y(mai_mai_n1263_));
  OAI220     m1235(.A0(mai_mai_n603_), .A1(g), .B0(mai_mai_n207_), .B1(c), .Y(mai_mai_n1264_));
  INV        m1236(.A(mai_mai_n1264_), .Y(mai_mai_n1265_));
  NO2        m1237(.A(mai_mai_n1265_), .B(mai_mai_n158_), .Y(mai_mai_n1266_));
  NO3        m1238(.A(mai_mai_n1253_), .B(mai_mai_n424_), .C(mai_mai_n329_), .Y(mai_mai_n1267_));
  NO3        m1239(.A(mai_mai_n1267_), .B(mai_mai_n1266_), .C(mai_mai_n1263_), .Y(mai_mai_n1268_));
  NO2        m1240(.A(mai_mai_n971_), .B(h), .Y(mai_mai_n1269_));
  NA3        m1241(.A(mai_mai_n1269_), .B(d), .C(mai_mai_n935_), .Y(mai_mai_n1270_));
  NO2        m1242(.A(mai_mai_n1270_), .B(c), .Y(mai_mai_n1271_));
  NOi21      m1243(.An(d), .B(f), .Y(mai_mai_n1272_));
  NO2        m1244(.A(mai_mai_n1201_), .B(f), .Y(mai_mai_n1273_));
  INV        m1245(.A(mai_mai_n1271_), .Y(mai_mai_n1274_));
  NA3        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1268_), .C(mai_mai_n1259_), .Y(mai_mai_n1275_));
  OAI210     m1247(.A0(mai_mai_n1250_), .A1(mai_mai_n1204_), .B0(mai_mai_n800_), .Y(mai_mai_n1276_));
  NO2        m1248(.A(mai_mai_n932_), .B(mai_mai_n123_), .Y(mai_mai_n1277_));
  NA2        m1249(.A(mai_mai_n1277_), .B(mai_mai_n565_), .Y(mai_mai_n1278_));
  NA2        m1250(.A(mai_mai_n1278_), .B(mai_mai_n1276_), .Y(mai_mai_n1279_));
  NA2        m1251(.A(mai_mai_n1224_), .B(mai_mai_n1272_), .Y(mai_mai_n1280_));
  NO2        m1252(.A(mai_mai_n1280_), .B(m), .Y(mai_mai_n1281_));
  NO2        m1253(.A(mai_mai_n139_), .B(mai_mai_n161_), .Y(mai_mai_n1282_));
  OAI210     m1254(.A0(mai_mai_n1282_), .A1(mai_mai_n103_), .B0(mai_mai_n1237_), .Y(mai_mai_n1283_));
  INV        m1255(.A(mai_mai_n1283_), .Y(mai_mai_n1284_));
  NO3        m1256(.A(mai_mai_n1284_), .B(mai_mai_n1281_), .C(mai_mai_n1279_), .Y(mai_mai_n1285_));
  NO2        m1257(.A(mai_mai_n1200_), .B(e), .Y(mai_mai_n1286_));
  OAI210     m1258(.A0(mai_mai_n1273_), .A1(mai_mai_n1011_), .B0(mai_mai_n574_), .Y(mai_mai_n1287_));
  NO2        m1259(.A(mai_mai_n1287_), .B(mai_mai_n405_), .Y(mai_mai_n1288_));
  INV        m1260(.A(mai_mai_n1288_), .Y(mai_mai_n1289_));
  NO2        m1261(.A(mai_mai_n161_), .B(c), .Y(mai_mai_n1290_));
  OAI210     m1262(.A0(mai_mai_n1290_), .A1(mai_mai_n1286_), .B0(mai_mai_n159_), .Y(mai_mai_n1291_));
  AOI220     m1263(.A0(mai_mai_n1291_), .A1(mai_mai_n964_), .B0(mai_mai_n485_), .B1(mai_mai_n339_), .Y(mai_mai_n1292_));
  NA2        m1264(.A(mai_mai_n492_), .B(g), .Y(mai_mai_n1293_));
  NA2        m1265(.A(mai_mai_n1293_), .B(mai_mai_n1221_), .Y(mai_mai_n1294_));
  NO2        m1266(.A(mai_mai_n1252_), .B(f), .Y(mai_mai_n1295_));
  NA2        m1267(.A(mai_mai_n1011_), .B(a), .Y(mai_mai_n1296_));
  OAI220     m1268(.A0(mai_mai_n1296_), .A1(mai_mai_n64_), .B0(mai_mai_n1294_), .B1(mai_mai_n195_), .Y(mai_mai_n1297_));
  NA2        m1269(.A(mai_mai_n1295_), .B(mai_mai_n1207_), .Y(mai_mai_n1298_));
  OAI220     m1270(.A0(mai_mai_n1298_), .A1(mai_mai_n49_), .B0(mai_mai_n1340_), .B1(mai_mai_n157_), .Y(mai_mai_n1299_));
  NA4        m1271(.A(mai_mai_n983_), .B(mai_mai_n980_), .C(mai_mai_n203_), .D(mai_mai_n63_), .Y(mai_mai_n1300_));
  NA2        m1272(.A(mai_mai_n1205_), .B(mai_mai_n162_), .Y(mai_mai_n1301_));
  NO2        m1273(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1302_));
  OAI210     m1274(.A0(mai_mai_n1252_), .A1(mai_mai_n780_), .B0(mai_mai_n441_), .Y(mai_mai_n1303_));
  OAI210     m1275(.A0(mai_mai_n1303_), .A1(mai_mai_n986_), .B0(mai_mai_n1302_), .Y(mai_mai_n1304_));
  NO2        m1276(.A(m), .B(i), .Y(mai_mai_n1305_));
  NA3        m1277(.A(mai_mai_n1304_), .B(mai_mai_n1301_), .C(mai_mai_n1300_), .Y(mai_mai_n1306_));
  NO4        m1278(.A(mai_mai_n1306_), .B(mai_mai_n1299_), .C(mai_mai_n1297_), .D(mai_mai_n1292_), .Y(mai_mai_n1307_));
  NA3        m1279(.A(mai_mai_n1307_), .B(mai_mai_n1289_), .C(mai_mai_n1285_), .Y(mai_mai_n1308_));
  NA3        m1280(.A(mai_mai_n864_), .B(mai_mai_n130_), .C(mai_mai_n46_), .Y(mai_mai_n1309_));
  AOI210     m1281(.A0(mai_mai_n136_), .A1(c), .B0(mai_mai_n1309_), .Y(mai_mai_n1310_));
  INV        m1282(.A(mai_mai_n165_), .Y(mai_mai_n1311_));
  NA2        m1283(.A(mai_mai_n1311_), .B(mai_mai_n1269_), .Y(mai_mai_n1312_));
  AO210      m1284(.A0(mai_mai_n124_), .A1(l), .B0(mai_mai_n1248_), .Y(mai_mai_n1313_));
  NA2        m1285(.A(mai_mai_n1313_), .B(mai_mai_n1312_), .Y(mai_mai_n1314_));
  NO2        m1286(.A(mai_mai_n1314_), .B(mai_mai_n1310_), .Y(mai_mai_n1315_));
  NO4        m1287(.A(mai_mai_n207_), .B(mai_mai_n166_), .C(mai_mai_n237_), .D(k), .Y(mai_mai_n1316_));
  NOi21      m1288(.An(mai_mai_n1205_), .B(e), .Y(mai_mai_n1317_));
  NO2        m1289(.A(mai_mai_n1317_), .B(mai_mai_n1316_), .Y(mai_mai_n1318_));
  AN2        m1290(.A(mai_mai_n983_), .B(mai_mai_n969_), .Y(mai_mai_n1319_));
  AOI220     m1291(.A0(mai_mai_n1305_), .A1(mai_mai_n580_), .B0(mai_mai_n1342_), .B1(mai_mai_n144_), .Y(mai_mai_n1320_));
  NOi31      m1292(.An(mai_mai_n30_), .B(mai_mai_n1320_), .C(n), .Y(mai_mai_n1321_));
  AOI210     m1293(.A0(mai_mai_n1319_), .A1(mai_mai_n1055_), .B0(mai_mai_n1321_), .Y(mai_mai_n1322_));
  NA2        m1294(.A(mai_mai_n57_), .B(a), .Y(mai_mai_n1323_));
  NO2        m1295(.A(mai_mai_n1254_), .B(mai_mai_n1323_), .Y(mai_mai_n1324_));
  INV        m1296(.A(mai_mai_n1324_), .Y(mai_mai_n1325_));
  NA4        m1297(.A(mai_mai_n1325_), .B(mai_mai_n1322_), .C(mai_mai_n1318_), .D(mai_mai_n1315_), .Y(mai_mai_n1326_));
  OR4        m1298(.A(mai_mai_n1326_), .B(mai_mai_n1308_), .C(mai_mai_n1275_), .D(mai_mai_n1255_), .Y(mai04));
  NOi31      m1299(.An(mai_mai_n1250_), .B(mai_mai_n1251_), .C(mai_mai_n937_), .Y(mai_mai_n1328_));
  NA2        m1300(.A(mai_mai_n1273_), .B(mai_mai_n744_), .Y(mai_mai_n1329_));
  NO2        m1301(.A(mai_mai_n1329_), .B(mai_mai_n929_), .Y(mai_mai_n1330_));
  OR3        m1302(.A(mai_mai_n1330_), .B(mai_mai_n1328_), .C(mai_mai_n954_), .Y(mai_mai_n1331_));
  NO2        m1303(.A(mai_mai_n1207_), .B(mai_mai_n86_), .Y(mai_mai_n1332_));
  AOI210     m1304(.A0(mai_mai_n1332_), .A1(mai_mai_n948_), .B0(mai_mai_n1070_), .Y(mai_mai_n1333_));
  NA2        m1305(.A(mai_mai_n1333_), .B(mai_mai_n1097_), .Y(mai_mai_n1334_));
  NO4        m1306(.A(mai_mai_n1334_), .B(mai_mai_n1331_), .C(mai_mai_n961_), .D(mai_mai_n942_), .Y(mai_mai_n1335_));
  NA4        m1307(.A(mai_mai_n1335_), .B(mai_mai_n1013_), .C(mai_mai_n999_), .D(mai_mai_n989_), .Y(mai05));
  INV        m1308(.A(m), .Y(mai_mai_n1339_));
  INV        m1309(.A(mai_mai_n98_), .Y(mai_mai_n1340_));
  INV        m1310(.A(i), .Y(mai_mai_n1341_));
  INV        m1311(.A(j), .Y(mai_mai_n1342_));
  INV        m1312(.A(m), .Y(mai_mai_n1343_));
  INV        m1313(.A(b), .Y(mai_mai_n1344_));
  INV        m1314(.A(f), .Y(mai_mai_n1345_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(g), .Y(men_men_n50_));
  INV        u0022(.A(men_men_n50_), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n49_), .Y(men_men_n52_));
  NO3        u0024(.A(men_men_n52_), .B(men_men_n43_), .C(men_men_n39_), .Y(men_men_n53_));
  NO2        u0025(.A(men_men_n53_), .B(men_men_n32_), .Y(men_men_n54_));
  INV        u0026(.A(c), .Y(men_men_n55_));
  NA2        u0027(.A(e), .B(b), .Y(men_men_n56_));
  INV        u0028(.A(men_men_n56_), .Y(men_men_n57_));
  INV        u0029(.A(d), .Y(men_men_n58_));
  NA2        u0030(.A(g), .B(men_men_n58_), .Y(men_men_n59_));
  NAi21      u0031(.An(i), .B(h), .Y(men_men_n60_));
  NAi31      u0032(.An(i), .B(l), .C(j), .Y(men_men_n61_));
  NO2        u0033(.A(men_men_n60_), .B(men_men_n44_), .Y(men_men_n62_));
  NAi31      u0034(.An(men_men_n59_), .B(men_men_n62_), .C(men_men_n57_), .Y(men_men_n63_));
  NAi41      u0035(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n64_));
  NA2        u0036(.A(g), .B(f), .Y(men_men_n65_));
  NO2        u0037(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NAi21      u0038(.An(i), .B(j), .Y(men_men_n67_));
  NAi32      u0039(.An(n), .Bn(k), .C(m), .Y(men_men_n68_));
  NO2        u0040(.A(men_men_n68_), .B(men_men_n67_), .Y(men_men_n69_));
  NAi31      u0041(.An(l), .B(m), .C(k), .Y(men_men_n70_));
  NAi41      u0042(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n71_));
  NA2        u0043(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n72_));
  INV        u0044(.A(m), .Y(men_men_n73_));
  NOi21      u0045(.An(k), .B(l), .Y(men_men_n74_));
  AN4        u0046(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n75_));
  NOi31      u0047(.An(h), .B(g), .C(f), .Y(men_men_n76_));
  NOi32      u0048(.An(h), .Bn(g), .C(f), .Y(men_men_n77_));
  NA2        u0049(.A(men_men_n72_), .B(men_men_n63_), .Y(men_men_n78_));
  INV        u0050(.A(n), .Y(men_men_n79_));
  NOi32      u0051(.An(e), .Bn(b), .C(d), .Y(men_men_n80_));
  NA2        u0052(.A(men_men_n80_), .B(men_men_n79_), .Y(men_men_n81_));
  INV        u0053(.A(j), .Y(men_men_n82_));
  AN3        u0054(.A(m), .B(k), .C(i), .Y(men_men_n83_));
  NA3        u0055(.A(men_men_n83_), .B(men_men_n82_), .C(g), .Y(men_men_n84_));
  NO2        u0056(.A(men_men_n84_), .B(f), .Y(men_men_n85_));
  NAi32      u0057(.An(g), .Bn(f), .C(h), .Y(men_men_n86_));
  NAi31      u0058(.An(j), .B(m), .C(l), .Y(men_men_n87_));
  NO2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  NA2        u0060(.A(m), .B(l), .Y(men_men_n89_));
  NAi31      u0061(.An(k), .B(j), .C(g), .Y(men_men_n90_));
  NO3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(f), .Y(men_men_n91_));
  AN2        u0063(.A(j), .B(g), .Y(men_men_n92_));
  NOi32      u0064(.An(m), .Bn(l), .C(i), .Y(men_men_n93_));
  NOi21      u0065(.An(g), .B(i), .Y(men_men_n94_));
  NOi32      u0066(.An(m), .Bn(j), .C(k), .Y(men_men_n95_));
  AOI220     u0067(.A0(men_men_n95_), .A1(men_men_n94_), .B0(men_men_n93_), .B1(men_men_n92_), .Y(men_men_n96_));
  NO2        u0068(.A(men_men_n96_), .B(f), .Y(men_men_n97_));
  NO4        u0069(.A(men_men_n97_), .B(men_men_n91_), .C(men_men_n88_), .D(men_men_n85_), .Y(men_men_n98_));
  NAi41      u0070(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n99_));
  AN2        u0071(.A(e), .B(b), .Y(men_men_n100_));
  NOi31      u0072(.An(c), .B(h), .C(f), .Y(men_men_n101_));
  NA2        u0073(.A(men_men_n101_), .B(men_men_n100_), .Y(men_men_n102_));
  NO2        u0074(.A(men_men_n102_), .B(men_men_n99_), .Y(men_men_n103_));
  NOi21      u0075(.An(g), .B(f), .Y(men_men_n104_));
  NOi21      u0076(.An(i), .B(h), .Y(men_men_n105_));
  NA3        u0077(.A(men_men_n105_), .B(men_men_n104_), .C(men_men_n36_), .Y(men_men_n106_));
  INV        u0078(.A(a), .Y(men_men_n107_));
  NA2        u0079(.A(men_men_n100_), .B(men_men_n107_), .Y(men_men_n108_));
  INV        u0080(.A(l), .Y(men_men_n109_));
  NOi21      u0081(.An(m), .B(n), .Y(men_men_n110_));
  AN2        u0082(.A(k), .B(h), .Y(men_men_n111_));
  NO2        u0083(.A(men_men_n106_), .B(men_men_n81_), .Y(men_men_n112_));
  INV        u0084(.A(b), .Y(men_men_n113_));
  NA2        u0085(.A(l), .B(j), .Y(men_men_n114_));
  AN2        u0086(.A(k), .B(i), .Y(men_men_n115_));
  NA2        u0087(.A(men_men_n115_), .B(men_men_n114_), .Y(men_men_n116_));
  NA2        u0088(.A(g), .B(e), .Y(men_men_n117_));
  NOi32      u0089(.An(c), .Bn(a), .C(d), .Y(men_men_n118_));
  NA2        u0090(.A(men_men_n118_), .B(men_men_n110_), .Y(men_men_n119_));
  NO4        u0091(.A(men_men_n119_), .B(men_men_n117_), .C(men_men_n116_), .D(men_men_n113_), .Y(men_men_n120_));
  NO3        u0092(.A(men_men_n120_), .B(men_men_n112_), .C(men_men_n103_), .Y(men_men_n121_));
  OAI210     u0093(.A0(men_men_n98_), .A1(men_men_n81_), .B0(men_men_n121_), .Y(men_men_n122_));
  NOi31      u0094(.An(k), .B(m), .C(j), .Y(men_men_n123_));
  NA3        u0095(.A(men_men_n123_), .B(men_men_n76_), .C(men_men_n75_), .Y(men_men_n124_));
  NOi31      u0096(.An(k), .B(m), .C(i), .Y(men_men_n125_));
  NA3        u0097(.A(men_men_n125_), .B(men_men_n77_), .C(men_men_n75_), .Y(men_men_n126_));
  NA2        u0098(.A(men_men_n126_), .B(men_men_n124_), .Y(men_men_n127_));
  NOi32      u0099(.An(f), .Bn(b), .C(e), .Y(men_men_n128_));
  NAi21      u0100(.An(g), .B(h), .Y(men_men_n129_));
  NAi21      u0101(.An(m), .B(n), .Y(men_men_n130_));
  NAi21      u0102(.An(j), .B(k), .Y(men_men_n131_));
  NO3        u0103(.A(men_men_n131_), .B(men_men_n130_), .C(men_men_n129_), .Y(men_men_n132_));
  NAi41      u0104(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n133_));
  NAi31      u0105(.An(j), .B(k), .C(h), .Y(men_men_n134_));
  NO3        u0106(.A(men_men_n134_), .B(men_men_n133_), .C(men_men_n130_), .Y(men_men_n135_));
  AOI210     u0107(.A0(men_men_n132_), .A1(men_men_n128_), .B0(men_men_n135_), .Y(men_men_n136_));
  NO2        u0108(.A(k), .B(j), .Y(men_men_n137_));
  NO2        u0109(.A(men_men_n137_), .B(men_men_n130_), .Y(men_men_n138_));
  AN2        u0110(.A(k), .B(j), .Y(men_men_n139_));
  NAi21      u0111(.An(c), .B(b), .Y(men_men_n140_));
  NA2        u0112(.A(f), .B(d), .Y(men_men_n141_));
  NO4        u0113(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n139_), .D(men_men_n129_), .Y(men_men_n142_));
  NA2        u0114(.A(h), .B(c), .Y(men_men_n143_));
  NAi31      u0115(.An(f), .B(e), .C(b), .Y(men_men_n144_));
  NA2        u0116(.A(men_men_n142_), .B(men_men_n138_), .Y(men_men_n145_));
  NA2        u0117(.A(d), .B(b), .Y(men_men_n146_));
  NAi21      u0118(.An(e), .B(f), .Y(men_men_n147_));
  NO2        u0119(.A(men_men_n147_), .B(men_men_n146_), .Y(men_men_n148_));
  NA2        u0120(.A(b), .B(a), .Y(men_men_n149_));
  NAi21      u0121(.An(c), .B(d), .Y(men_men_n150_));
  NAi31      u0122(.An(l), .B(k), .C(h), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n130_), .B(men_men_n151_), .Y(men_men_n152_));
  NA2        u0124(.A(men_men_n152_), .B(men_men_n148_), .Y(men_men_n153_));
  NAi41      u0125(.An(men_men_n127_), .B(men_men_n153_), .C(men_men_n145_), .D(men_men_n136_), .Y(men_men_n154_));
  NAi31      u0126(.An(e), .B(f), .C(b), .Y(men_men_n155_));
  NOi21      u0127(.An(g), .B(d), .Y(men_men_n156_));
  NO2        u0128(.A(men_men_n156_), .B(men_men_n155_), .Y(men_men_n157_));
  NOi21      u0129(.An(h), .B(i), .Y(men_men_n158_));
  NOi21      u0130(.An(k), .B(m), .Y(men_men_n159_));
  NA3        u0131(.A(men_men_n159_), .B(men_men_n158_), .C(n), .Y(men_men_n160_));
  NOi21      u0132(.An(men_men_n157_), .B(men_men_n160_), .Y(men_men_n161_));
  NOi21      u0133(.An(h), .B(g), .Y(men_men_n162_));
  NO2        u0134(.A(men_men_n141_), .B(men_men_n140_), .Y(men_men_n163_));
  NA2        u0135(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  NAi31      u0136(.An(l), .B(j), .C(h), .Y(men_men_n165_));
  NO2        u0137(.A(men_men_n165_), .B(men_men_n49_), .Y(men_men_n166_));
  NA2        u0138(.A(men_men_n166_), .B(men_men_n66_), .Y(men_men_n167_));
  NOi32      u0139(.An(n), .Bn(k), .C(m), .Y(men_men_n168_));
  NA2        u0140(.A(l), .B(i), .Y(men_men_n169_));
  NA2        u0141(.A(men_men_n169_), .B(men_men_n168_), .Y(men_men_n170_));
  OAI210     u0142(.A0(men_men_n170_), .A1(men_men_n164_), .B0(men_men_n167_), .Y(men_men_n171_));
  NAi31      u0143(.An(d), .B(f), .C(c), .Y(men_men_n172_));
  NAi31      u0144(.An(e), .B(f), .C(c), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  NA2        u0146(.A(j), .B(h), .Y(men_men_n175_));
  OR3        u0147(.A(n), .B(m), .C(k), .Y(men_men_n176_));
  NO2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  NAi32      u0149(.An(m), .Bn(k), .C(n), .Y(men_men_n178_));
  NO2        u0150(.A(men_men_n178_), .B(men_men_n175_), .Y(men_men_n179_));
  AOI220     u0151(.A0(men_men_n179_), .A1(men_men_n157_), .B0(men_men_n177_), .B1(men_men_n174_), .Y(men_men_n180_));
  NO2        u0152(.A(n), .B(m), .Y(men_men_n181_));
  NAi21      u0153(.An(f), .B(e), .Y(men_men_n182_));
  NA2        u0154(.A(d), .B(c), .Y(men_men_n183_));
  NAi31      u0155(.An(m), .B(n), .C(b), .Y(men_men_n184_));
  NAi21      u0156(.An(h), .B(f), .Y(men_men_n185_));
  NO2        u0157(.A(men_men_n184_), .B(men_men_n150_), .Y(men_men_n186_));
  NOi32      u0158(.An(f), .Bn(c), .C(d), .Y(men_men_n187_));
  NOi32      u0159(.An(f), .Bn(c), .C(e), .Y(men_men_n188_));
  NO2        u0160(.A(men_men_n188_), .B(men_men_n187_), .Y(men_men_n189_));
  NO3        u0161(.A(n), .B(m), .C(j), .Y(men_men_n190_));
  NA2        u0162(.A(men_men_n190_), .B(men_men_n111_), .Y(men_men_n191_));
  OR2        u0163(.A(men_men_n191_), .B(men_men_n189_), .Y(men_men_n192_));
  NA2        u0164(.A(men_men_n192_), .B(men_men_n180_), .Y(men_men_n193_));
  OR4        u0165(.A(men_men_n193_), .B(men_men_n171_), .C(men_men_n161_), .D(men_men_n154_), .Y(men_men_n194_));
  NO4        u0166(.A(men_men_n194_), .B(men_men_n122_), .C(men_men_n78_), .D(men_men_n54_), .Y(men_men_n195_));
  NA3        u0167(.A(m), .B(men_men_n109_), .C(j), .Y(men_men_n196_));
  NAi31      u0168(.An(n), .B(h), .C(g), .Y(men_men_n197_));
  NO2        u0169(.A(men_men_n197_), .B(men_men_n196_), .Y(men_men_n198_));
  NOi32      u0170(.An(m), .Bn(k), .C(l), .Y(men_men_n199_));
  NA3        u0171(.A(men_men_n199_), .B(men_men_n82_), .C(g), .Y(men_men_n200_));
  NO2        u0172(.A(men_men_n200_), .B(n), .Y(men_men_n201_));
  NOi21      u0173(.An(k), .B(j), .Y(men_men_n202_));
  NA4        u0174(.A(men_men_n202_), .B(men_men_n110_), .C(i), .D(g), .Y(men_men_n203_));
  AN2        u0175(.A(i), .B(g), .Y(men_men_n204_));
  NA3        u0176(.A(men_men_n74_), .B(men_men_n204_), .C(men_men_n110_), .Y(men_men_n205_));
  NA2        u0177(.A(men_men_n205_), .B(men_men_n203_), .Y(men_men_n206_));
  NO3        u0178(.A(men_men_n206_), .B(men_men_n201_), .C(men_men_n198_), .Y(men_men_n207_));
  NAi41      u0179(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n208_));
  INV        u0180(.A(men_men_n208_), .Y(men_men_n209_));
  INV        u0181(.A(f), .Y(men_men_n210_));
  INV        u0182(.A(g), .Y(men_men_n211_));
  NOi31      u0183(.An(i), .B(j), .C(h), .Y(men_men_n212_));
  NOi21      u0184(.An(l), .B(m), .Y(men_men_n213_));
  NA2        u0185(.A(men_men_n213_), .B(men_men_n212_), .Y(men_men_n214_));
  NO2        u0186(.A(men_men_n207_), .B(men_men_n32_), .Y(men_men_n215_));
  NOi21      u0187(.An(n), .B(m), .Y(men_men_n216_));
  NOi32      u0188(.An(l), .Bn(i), .C(j), .Y(men_men_n217_));
  NA2        u0189(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n218_));
  OR2        u0190(.A(men_men_n218_), .B(men_men_n102_), .Y(men_men_n219_));
  NAi21      u0191(.An(j), .B(h), .Y(men_men_n220_));
  XN2        u0192(.A(i), .B(h), .Y(men_men_n221_));
  NA2        u0193(.A(men_men_n221_), .B(men_men_n220_), .Y(men_men_n222_));
  NOi31      u0194(.An(k), .B(n), .C(m), .Y(men_men_n223_));
  NOi31      u0195(.An(men_men_n223_), .B(men_men_n183_), .C(men_men_n182_), .Y(men_men_n224_));
  NA2        u0196(.A(men_men_n224_), .B(men_men_n222_), .Y(men_men_n225_));
  NAi31      u0197(.An(f), .B(e), .C(c), .Y(men_men_n226_));
  NO4        u0198(.A(men_men_n226_), .B(men_men_n176_), .C(men_men_n175_), .D(men_men_n58_), .Y(men_men_n227_));
  NA4        u0199(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n228_));
  NAi32      u0200(.An(m), .Bn(i), .C(k), .Y(men_men_n229_));
  NO3        u0201(.A(men_men_n229_), .B(men_men_n86_), .C(men_men_n228_), .Y(men_men_n230_));
  INV        u0202(.A(k), .Y(men_men_n231_));
  NO2        u0203(.A(men_men_n230_), .B(men_men_n227_), .Y(men_men_n232_));
  NAi21      u0204(.An(n), .B(a), .Y(men_men_n233_));
  NO2        u0205(.A(men_men_n233_), .B(men_men_n146_), .Y(men_men_n234_));
  NAi41      u0206(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n235_));
  NO2        u0207(.A(men_men_n235_), .B(e), .Y(men_men_n236_));
  NO3        u0208(.A(men_men_n147_), .B(men_men_n90_), .C(men_men_n89_), .Y(men_men_n237_));
  OAI210     u0209(.A0(men_men_n237_), .A1(men_men_n236_), .B0(men_men_n234_), .Y(men_men_n238_));
  AN4        u0210(.A(men_men_n238_), .B(men_men_n232_), .C(men_men_n225_), .D(men_men_n219_), .Y(men_men_n239_));
  OR2        u0211(.A(h), .B(g), .Y(men_men_n240_));
  NAi41      u0212(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n241_));
  NO2        u0213(.A(men_men_n241_), .B(men_men_n210_), .Y(men_men_n242_));
  NA2        u0214(.A(men_men_n159_), .B(men_men_n105_), .Y(men_men_n243_));
  NAi21      u0215(.An(men_men_n243_), .B(men_men_n242_), .Y(men_men_n244_));
  NO2        u0216(.A(n), .B(a), .Y(men_men_n245_));
  NAi31      u0217(.An(men_men_n235_), .B(men_men_n245_), .C(men_men_n100_), .Y(men_men_n246_));
  AN2        u0218(.A(men_men_n246_), .B(men_men_n244_), .Y(men_men_n247_));
  NAi21      u0219(.An(h), .B(i), .Y(men_men_n248_));
  NA2        u0220(.A(men_men_n181_), .B(k), .Y(men_men_n249_));
  NO2        u0221(.A(men_men_n249_), .B(men_men_n248_), .Y(men_men_n250_));
  NA2        u0222(.A(men_men_n250_), .B(men_men_n187_), .Y(men_men_n251_));
  NA2        u0223(.A(men_men_n251_), .B(men_men_n247_), .Y(men_men_n252_));
  NO2        u0224(.A(men_men_n71_), .B(men_men_n73_), .Y(men_men_n253_));
  NOi32      u0225(.An(l), .Bn(j), .C(i), .Y(men_men_n254_));
  AOI210     u0226(.A0(men_men_n74_), .A1(men_men_n82_), .B0(men_men_n254_), .Y(men_men_n255_));
  NO2        u0227(.A(men_men_n248_), .B(men_men_n44_), .Y(men_men_n256_));
  NAi21      u0228(.An(f), .B(g), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n257_), .B(men_men_n64_), .Y(men_men_n258_));
  NO2        u0230(.A(men_men_n68_), .B(men_men_n114_), .Y(men_men_n259_));
  AOI220     u0231(.A0(men_men_n259_), .A1(men_men_n258_), .B0(men_men_n256_), .B1(men_men_n66_), .Y(men_men_n260_));
  INV        u0232(.A(men_men_n260_), .Y(men_men_n261_));
  NO3        u0233(.A(men_men_n131_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n262_));
  NOi41      u0234(.An(men_men_n239_), .B(men_men_n261_), .C(men_men_n252_), .D(men_men_n215_), .Y(men_men_n263_));
  NO4        u0235(.A(men_men_n198_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n264_));
  NO2        u0236(.A(men_men_n264_), .B(men_men_n108_), .Y(men_men_n265_));
  NA2        u0237(.A(c), .B(b), .Y(men_men_n266_));
  NAi21      u0238(.An(h), .B(g), .Y(men_men_n267_));
  OR4        u0239(.A(men_men_n267_), .B(men_men_n266_), .C(men_men_n218_), .D(e), .Y(men_men_n268_));
  NAi31      u0240(.An(g), .B(k), .C(h), .Y(men_men_n269_));
  NO3        u0241(.A(men_men_n130_), .B(men_men_n269_), .C(l), .Y(men_men_n270_));
  NAi31      u0242(.An(e), .B(d), .C(a), .Y(men_men_n271_));
  NA2        u0243(.A(men_men_n270_), .B(men_men_n128_), .Y(men_men_n272_));
  NA2        u0244(.A(men_men_n272_), .B(men_men_n268_), .Y(men_men_n273_));
  NA3        u0245(.A(men_men_n159_), .B(men_men_n158_), .C(men_men_n79_), .Y(men_men_n274_));
  NO2        u0246(.A(men_men_n274_), .B(men_men_n189_), .Y(men_men_n275_));
  INV        u0247(.A(men_men_n275_), .Y(men_men_n276_));
  NA3        u0248(.A(e), .B(c), .C(b), .Y(men_men_n277_));
  NO2        u0249(.A(men_men_n59_), .B(men_men_n277_), .Y(men_men_n278_));
  NAi32      u0250(.An(k), .Bn(i), .C(j), .Y(men_men_n279_));
  NAi31      u0251(.An(h), .B(l), .C(i), .Y(men_men_n280_));
  NA3        u0252(.A(men_men_n280_), .B(men_men_n279_), .C(men_men_n165_), .Y(men_men_n281_));
  NOi21      u0253(.An(men_men_n281_), .B(men_men_n49_), .Y(men_men_n282_));
  OAI210     u0254(.A0(men_men_n258_), .A1(men_men_n278_), .B0(men_men_n282_), .Y(men_men_n283_));
  NAi21      u0255(.An(l), .B(k), .Y(men_men_n284_));
  NO2        u0256(.A(men_men_n284_), .B(men_men_n49_), .Y(men_men_n285_));
  NOi21      u0257(.An(l), .B(j), .Y(men_men_n286_));
  NA2        u0258(.A(men_men_n162_), .B(men_men_n286_), .Y(men_men_n287_));
  NA3        u0259(.A(men_men_n115_), .B(men_men_n114_), .C(g), .Y(men_men_n288_));
  OR3        u0260(.A(men_men_n71_), .B(men_men_n73_), .C(e), .Y(men_men_n289_));
  AOI210     u0261(.A0(men_men_n288_), .A1(men_men_n287_), .B0(men_men_n289_), .Y(men_men_n290_));
  INV        u0262(.A(men_men_n290_), .Y(men_men_n291_));
  NAi32      u0263(.An(j), .Bn(h), .C(i), .Y(men_men_n292_));
  NAi21      u0264(.An(m), .B(l), .Y(men_men_n293_));
  NO3        u0265(.A(men_men_n293_), .B(men_men_n292_), .C(men_men_n79_), .Y(men_men_n294_));
  NA2        u0266(.A(h), .B(g), .Y(men_men_n295_));
  NA2        u0267(.A(men_men_n168_), .B(men_men_n45_), .Y(men_men_n296_));
  NO2        u0268(.A(men_men_n296_), .B(men_men_n295_), .Y(men_men_n297_));
  OAI210     u0269(.A0(men_men_n297_), .A1(men_men_n294_), .B0(men_men_n163_), .Y(men_men_n298_));
  NA4        u0270(.A(men_men_n298_), .B(men_men_n291_), .C(men_men_n283_), .D(men_men_n276_), .Y(men_men_n299_));
  NO2        u0271(.A(men_men_n144_), .B(d), .Y(men_men_n300_));
  NA2        u0272(.A(men_men_n300_), .B(men_men_n52_), .Y(men_men_n301_));
  NO2        u0273(.A(men_men_n102_), .B(men_men_n99_), .Y(men_men_n302_));
  NAi32      u0274(.An(n), .Bn(m), .C(l), .Y(men_men_n303_));
  NO2        u0275(.A(men_men_n303_), .B(men_men_n292_), .Y(men_men_n304_));
  NO2        u0276(.A(men_men_n119_), .B(men_men_n113_), .Y(men_men_n305_));
  NAi31      u0277(.An(k), .B(l), .C(j), .Y(men_men_n306_));
  OAI210     u0278(.A0(men_men_n284_), .A1(j), .B0(men_men_n306_), .Y(men_men_n307_));
  NOi21      u0279(.An(men_men_n307_), .B(men_men_n117_), .Y(men_men_n308_));
  NA2        u0280(.A(men_men_n308_), .B(men_men_n305_), .Y(men_men_n309_));
  NA2        u0281(.A(men_men_n309_), .B(men_men_n301_), .Y(men_men_n310_));
  NO4        u0282(.A(men_men_n310_), .B(men_men_n299_), .C(men_men_n273_), .D(men_men_n265_), .Y(men_men_n311_));
  NA2        u0283(.A(men_men_n250_), .B(men_men_n188_), .Y(men_men_n312_));
  NAi21      u0284(.An(m), .B(k), .Y(men_men_n313_));
  NO2        u0285(.A(men_men_n221_), .B(men_men_n313_), .Y(men_men_n314_));
  NAi41      u0286(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n315_));
  NO2        u0287(.A(men_men_n315_), .B(e), .Y(men_men_n316_));
  NA2        u0288(.A(men_men_n316_), .B(men_men_n314_), .Y(men_men_n317_));
  NAi31      u0289(.An(i), .B(l), .C(h), .Y(men_men_n318_));
  NO4        u0290(.A(men_men_n318_), .B(e), .C(men_men_n71_), .D(men_men_n73_), .Y(men_men_n319_));
  NA2        u0291(.A(e), .B(c), .Y(men_men_n320_));
  NO3        u0292(.A(men_men_n320_), .B(n), .C(d), .Y(men_men_n321_));
  NOi21      u0293(.An(f), .B(h), .Y(men_men_n322_));
  NA2        u0294(.A(men_men_n322_), .B(men_men_n115_), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n323_), .B(men_men_n211_), .Y(men_men_n324_));
  NAi31      u0296(.An(d), .B(e), .C(b), .Y(men_men_n325_));
  NO2        u0297(.A(men_men_n130_), .B(men_men_n325_), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n326_), .B(men_men_n324_), .Y(men_men_n327_));
  NAi41      u0299(.An(men_men_n319_), .B(men_men_n327_), .C(men_men_n317_), .D(men_men_n312_), .Y(men_men_n328_));
  NA2        u0300(.A(men_men_n245_), .B(men_men_n100_), .Y(men_men_n329_));
  NOi31      u0301(.An(l), .B(n), .C(m), .Y(men_men_n330_));
  NA2        u0302(.A(men_men_n330_), .B(men_men_n212_), .Y(men_men_n331_));
  NO2        u0303(.A(men_men_n331_), .B(men_men_n189_), .Y(men_men_n332_));
  NAi32      u0304(.An(m), .Bn(j), .C(k), .Y(men_men_n333_));
  NAi41      u0305(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n334_));
  NOi31      u0306(.An(j), .B(m), .C(k), .Y(men_men_n335_));
  AN3        u0307(.A(h), .B(g), .C(f), .Y(men_men_n336_));
  NOi32      u0308(.An(m), .Bn(j), .C(l), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n337_), .B(men_men_n93_), .Y(men_men_n338_));
  NAi32      u0310(.An(men_men_n338_), .Bn(men_men_n197_), .C(men_men_n300_), .Y(men_men_n339_));
  NO2        u0311(.A(men_men_n293_), .B(men_men_n292_), .Y(men_men_n340_));
  NO2        u0312(.A(men_men_n214_), .B(g), .Y(men_men_n341_));
  INV        u0313(.A(men_men_n155_), .Y(men_men_n342_));
  AOI220     u0314(.A0(men_men_n342_), .A1(men_men_n341_), .B0(men_men_n242_), .B1(men_men_n340_), .Y(men_men_n343_));
  INV        u0315(.A(men_men_n229_), .Y(men_men_n344_));
  NA3        u0316(.A(men_men_n344_), .B(men_men_n336_), .C(men_men_n209_), .Y(men_men_n345_));
  NA3        u0317(.A(men_men_n345_), .B(men_men_n343_), .C(men_men_n339_), .Y(men_men_n346_));
  NA3        u0318(.A(h), .B(g), .C(f), .Y(men_men_n347_));
  NA2        u0319(.A(men_men_n162_), .B(e), .Y(men_men_n348_));
  NO2        u0320(.A(men_men_n348_), .B(men_men_n41_), .Y(men_men_n349_));
  NA2        u0321(.A(men_men_n349_), .B(men_men_n305_), .Y(men_men_n350_));
  NOi32      u0322(.An(j), .Bn(g), .C(i), .Y(men_men_n351_));
  NA3        u0323(.A(men_men_n351_), .B(men_men_n284_), .C(men_men_n110_), .Y(men_men_n352_));
  OR2        u0324(.A(men_men_n108_), .B(men_men_n352_), .Y(men_men_n353_));
  NOi32      u0325(.An(e), .Bn(b), .C(a), .Y(men_men_n354_));
  AN2        u0326(.A(l), .B(j), .Y(men_men_n355_));
  NO2        u0327(.A(men_men_n313_), .B(men_men_n355_), .Y(men_men_n356_));
  NO3        u0328(.A(men_men_n315_), .B(e), .C(men_men_n211_), .Y(men_men_n357_));
  NA3        u0329(.A(men_men_n205_), .B(men_men_n203_), .C(men_men_n35_), .Y(men_men_n358_));
  AOI220     u0330(.A0(men_men_n358_), .A1(men_men_n354_), .B0(men_men_n357_), .B1(men_men_n356_), .Y(men_men_n359_));
  NO2        u0331(.A(men_men_n325_), .B(n), .Y(men_men_n360_));
  NA2        u0332(.A(men_men_n204_), .B(k), .Y(men_men_n361_));
  NA3        u0333(.A(m), .B(men_men_n109_), .C(men_men_n210_), .Y(men_men_n362_));
  NA4        u0334(.A(men_men_n199_), .B(men_men_n82_), .C(g), .D(men_men_n210_), .Y(men_men_n363_));
  OAI210     u0335(.A0(men_men_n362_), .A1(men_men_n361_), .B0(men_men_n363_), .Y(men_men_n364_));
  NAi41      u0336(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n365_));
  NA2        u0337(.A(men_men_n50_), .B(men_men_n110_), .Y(men_men_n366_));
  NA2        u0338(.A(men_men_n364_), .B(men_men_n360_), .Y(men_men_n367_));
  NA4        u0339(.A(men_men_n367_), .B(men_men_n359_), .C(men_men_n353_), .D(men_men_n350_), .Y(men_men_n368_));
  NO4        u0340(.A(men_men_n368_), .B(men_men_n346_), .C(men_men_n332_), .D(men_men_n328_), .Y(men_men_n369_));
  NA4        u0341(.A(men_men_n369_), .B(men_men_n311_), .C(men_men_n263_), .D(men_men_n195_), .Y(men10));
  NA3        u0342(.A(m), .B(k), .C(i), .Y(men_men_n371_));
  NO3        u0343(.A(men_men_n371_), .B(j), .C(men_men_n211_), .Y(men_men_n372_));
  NOi21      u0344(.An(e), .B(f), .Y(men_men_n373_));
  NO4        u0345(.A(men_men_n150_), .B(men_men_n373_), .C(n), .D(men_men_n107_), .Y(men_men_n374_));
  NAi31      u0346(.An(b), .B(f), .C(c), .Y(men_men_n375_));
  INV        u0347(.A(men_men_n375_), .Y(men_men_n376_));
  NOi32      u0348(.An(k), .Bn(h), .C(j), .Y(men_men_n377_));
  NA2        u0349(.A(men_men_n377_), .B(men_men_n216_), .Y(men_men_n378_));
  INV        u0350(.A(men_men_n378_), .Y(men_men_n379_));
  AOI220     u0351(.A0(men_men_n379_), .A1(men_men_n376_), .B0(men_men_n374_), .B1(men_men_n372_), .Y(men_men_n380_));
  AN2        u0352(.A(j), .B(h), .Y(men_men_n381_));
  NO3        u0353(.A(n), .B(m), .C(k), .Y(men_men_n382_));
  NA2        u0354(.A(men_men_n382_), .B(men_men_n381_), .Y(men_men_n383_));
  NO3        u0355(.A(men_men_n383_), .B(men_men_n150_), .C(men_men_n210_), .Y(men_men_n384_));
  OR2        u0356(.A(m), .B(k), .Y(men_men_n385_));
  NO2        u0357(.A(men_men_n175_), .B(men_men_n385_), .Y(men_men_n386_));
  NA4        u0358(.A(n), .B(f), .C(c), .D(men_men_n113_), .Y(men_men_n387_));
  NOi21      u0359(.An(men_men_n386_), .B(men_men_n387_), .Y(men_men_n388_));
  NOi32      u0360(.An(d), .Bn(a), .C(c), .Y(men_men_n389_));
  NA2        u0361(.A(men_men_n389_), .B(men_men_n182_), .Y(men_men_n390_));
  NAi21      u0362(.An(i), .B(g), .Y(men_men_n391_));
  NAi31      u0363(.An(k), .B(m), .C(j), .Y(men_men_n392_));
  NO3        u0364(.A(men_men_n392_), .B(men_men_n391_), .C(n), .Y(men_men_n393_));
  NOi21      u0365(.An(men_men_n393_), .B(men_men_n390_), .Y(men_men_n394_));
  NO3        u0366(.A(men_men_n394_), .B(men_men_n388_), .C(men_men_n384_), .Y(men_men_n395_));
  NO2        u0367(.A(men_men_n387_), .B(men_men_n293_), .Y(men_men_n396_));
  NOi32      u0368(.An(f), .Bn(d), .C(c), .Y(men_men_n397_));
  AOI220     u0369(.A0(men_men_n397_), .A1(men_men_n304_), .B0(men_men_n396_), .B1(men_men_n212_), .Y(men_men_n398_));
  NA3        u0370(.A(men_men_n398_), .B(men_men_n395_), .C(men_men_n380_), .Y(men_men_n399_));
  NO2        u0371(.A(men_men_n58_), .B(men_men_n113_), .Y(men_men_n400_));
  NA2        u0372(.A(men_men_n245_), .B(men_men_n400_), .Y(men_men_n401_));
  INV        u0373(.A(e), .Y(men_men_n402_));
  NA2        u0374(.A(men_men_n46_), .B(e), .Y(men_men_n403_));
  OAI220     u0375(.A0(men_men_n403_), .A1(men_men_n196_), .B0(men_men_n200_), .B1(men_men_n402_), .Y(men_men_n404_));
  AN2        u0376(.A(g), .B(e), .Y(men_men_n405_));
  NA3        u0377(.A(men_men_n405_), .B(men_men_n199_), .C(i), .Y(men_men_n406_));
  OAI210     u0378(.A0(men_men_n84_), .A1(men_men_n402_), .B0(men_men_n406_), .Y(men_men_n407_));
  NO2        u0379(.A(men_men_n96_), .B(men_men_n402_), .Y(men_men_n408_));
  NO2        u0380(.A(men_men_n408_), .B(men_men_n407_), .Y(men_men_n409_));
  NOi32      u0381(.An(h), .Bn(e), .C(g), .Y(men_men_n410_));
  NA3        u0382(.A(men_men_n410_), .B(men_men_n286_), .C(m), .Y(men_men_n411_));
  NOi21      u0383(.An(g), .B(h), .Y(men_men_n412_));
  AN3        u0384(.A(m), .B(l), .C(i), .Y(men_men_n413_));
  NA3        u0385(.A(men_men_n413_), .B(men_men_n412_), .C(e), .Y(men_men_n414_));
  AN3        u0386(.A(h), .B(g), .C(e), .Y(men_men_n415_));
  NA2        u0387(.A(men_men_n415_), .B(men_men_n93_), .Y(men_men_n416_));
  AN3        u0388(.A(men_men_n416_), .B(men_men_n414_), .C(men_men_n411_), .Y(men_men_n417_));
  AOI210     u0389(.A0(men_men_n417_), .A1(men_men_n409_), .B0(men_men_n401_), .Y(men_men_n418_));
  NA3        u0390(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n419_));
  NO2        u0391(.A(men_men_n419_), .B(men_men_n401_), .Y(men_men_n420_));
  NA2        u0392(.A(men_men_n389_), .B(men_men_n79_), .Y(men_men_n421_));
  NAi31      u0393(.An(b), .B(c), .C(a), .Y(men_men_n422_));
  NO2        u0394(.A(men_men_n422_), .B(n), .Y(men_men_n423_));
  NA2        u0395(.A(men_men_n50_), .B(m), .Y(men_men_n424_));
  NO2        u0396(.A(men_men_n424_), .B(men_men_n147_), .Y(men_men_n425_));
  NA2        u0397(.A(men_men_n425_), .B(men_men_n423_), .Y(men_men_n426_));
  INV        u0398(.A(men_men_n426_), .Y(men_men_n427_));
  NO4        u0399(.A(men_men_n427_), .B(men_men_n420_), .C(men_men_n418_), .D(men_men_n399_), .Y(men_men_n428_));
  NA2        u0400(.A(i), .B(g), .Y(men_men_n429_));
  NO3        u0401(.A(men_men_n271_), .B(men_men_n429_), .C(c), .Y(men_men_n430_));
  NOi21      u0402(.An(a), .B(n), .Y(men_men_n431_));
  NOi21      u0403(.An(d), .B(c), .Y(men_men_n432_));
  NA2        u0404(.A(men_men_n432_), .B(men_men_n431_), .Y(men_men_n433_));
  NA3        u0405(.A(i), .B(g), .C(f), .Y(men_men_n434_));
  OR2        u0406(.A(men_men_n434_), .B(men_men_n70_), .Y(men_men_n435_));
  NA2        u0407(.A(men_men_n413_), .B(men_men_n412_), .Y(men_men_n436_));
  AOI210     u0408(.A0(men_men_n436_), .A1(men_men_n435_), .B0(men_men_n433_), .Y(men_men_n437_));
  AOI210     u0409(.A0(men_men_n430_), .A1(men_men_n285_), .B0(men_men_n437_), .Y(men_men_n438_));
  OR2        u0410(.A(n), .B(m), .Y(men_men_n439_));
  NO2        u0411(.A(men_men_n439_), .B(men_men_n151_), .Y(men_men_n440_));
  NO2        u0412(.A(men_men_n183_), .B(men_men_n147_), .Y(men_men_n441_));
  OAI210     u0413(.A0(men_men_n440_), .A1(men_men_n177_), .B0(men_men_n441_), .Y(men_men_n442_));
  INV        u0414(.A(men_men_n366_), .Y(men_men_n443_));
  NA3        u0415(.A(men_men_n443_), .B(men_men_n354_), .C(d), .Y(men_men_n444_));
  NO2        u0416(.A(men_men_n422_), .B(men_men_n49_), .Y(men_men_n445_));
  NAi21      u0417(.An(k), .B(j), .Y(men_men_n446_));
  NAi21      u0418(.An(e), .B(d), .Y(men_men_n447_));
  INV        u0419(.A(men_men_n447_), .Y(men_men_n448_));
  NO2        u0420(.A(men_men_n249_), .B(men_men_n210_), .Y(men_men_n449_));
  NA3        u0421(.A(men_men_n449_), .B(men_men_n448_), .C(men_men_n222_), .Y(men_men_n450_));
  NA3        u0422(.A(men_men_n450_), .B(men_men_n444_), .C(men_men_n442_), .Y(men_men_n451_));
  NO2        u0423(.A(men_men_n331_), .B(men_men_n210_), .Y(men_men_n452_));
  NA2        u0424(.A(men_men_n452_), .B(men_men_n448_), .Y(men_men_n453_));
  NAi31      u0425(.An(g), .B(f), .C(c), .Y(men_men_n454_));
  INV        u0426(.A(men_men_n453_), .Y(men_men_n455_));
  NOi41      u0427(.An(men_men_n438_), .B(men_men_n455_), .C(men_men_n451_), .D(men_men_n261_), .Y(men_men_n456_));
  NOi32      u0428(.An(c), .Bn(a), .C(b), .Y(men_men_n457_));
  NA2        u0429(.A(men_men_n457_), .B(men_men_n110_), .Y(men_men_n458_));
  INV        u0430(.A(men_men_n269_), .Y(men_men_n459_));
  AN2        u0431(.A(e), .B(d), .Y(men_men_n460_));
  NA2        u0432(.A(men_men_n460_), .B(men_men_n459_), .Y(men_men_n461_));
  INV        u0433(.A(men_men_n147_), .Y(men_men_n462_));
  NO2        u0434(.A(men_men_n129_), .B(men_men_n41_), .Y(men_men_n463_));
  NO2        u0435(.A(men_men_n65_), .B(e), .Y(men_men_n464_));
  NOi31      u0436(.An(j), .B(k), .C(i), .Y(men_men_n465_));
  NOi21      u0437(.An(men_men_n165_), .B(men_men_n465_), .Y(men_men_n466_));
  AOI210     u0438(.A0(men_men_n463_), .A1(men_men_n462_), .B0(men_men_n464_), .Y(men_men_n467_));
  AOI210     u0439(.A0(men_men_n467_), .A1(men_men_n461_), .B0(men_men_n458_), .Y(men_men_n468_));
  NO2        u0440(.A(men_men_n206_), .B(men_men_n201_), .Y(men_men_n469_));
  NOi21      u0441(.An(a), .B(b), .Y(men_men_n470_));
  NA3        u0442(.A(e), .B(d), .C(c), .Y(men_men_n471_));
  NAi21      u0443(.An(men_men_n471_), .B(men_men_n470_), .Y(men_men_n472_));
  AOI210     u0444(.A0(men_men_n264_), .A1(men_men_n469_), .B0(men_men_n472_), .Y(men_men_n473_));
  NO4        u0445(.A(men_men_n185_), .B(men_men_n99_), .C(men_men_n55_), .D(b), .Y(men_men_n474_));
  NA2        u0446(.A(men_men_n376_), .B(men_men_n152_), .Y(men_men_n475_));
  OR2        u0447(.A(k), .B(j), .Y(men_men_n476_));
  NA2        u0448(.A(l), .B(k), .Y(men_men_n477_));
  NA3        u0449(.A(men_men_n477_), .B(men_men_n476_), .C(men_men_n216_), .Y(men_men_n478_));
  AOI210     u0450(.A0(men_men_n229_), .A1(men_men_n333_), .B0(men_men_n79_), .Y(men_men_n479_));
  NOi21      u0451(.An(men_men_n478_), .B(men_men_n479_), .Y(men_men_n480_));
  OR3        u0452(.A(men_men_n480_), .B(men_men_n143_), .C(men_men_n133_), .Y(men_men_n481_));
  NA2        u0453(.A(men_men_n126_), .B(men_men_n124_), .Y(men_men_n482_));
  NA2        u0454(.A(men_men_n389_), .B(men_men_n110_), .Y(men_men_n483_));
  NO4        u0455(.A(men_men_n483_), .B(men_men_n90_), .C(men_men_n109_), .D(e), .Y(men_men_n484_));
  NO3        u0456(.A(men_men_n421_), .B(men_men_n87_), .C(men_men_n129_), .Y(men_men_n485_));
  NO4        u0457(.A(men_men_n485_), .B(men_men_n484_), .C(men_men_n482_), .D(men_men_n319_), .Y(men_men_n486_));
  NA3        u0458(.A(men_men_n486_), .B(men_men_n481_), .C(men_men_n475_), .Y(men_men_n487_));
  NO3        u0459(.A(men_men_n487_), .B(men_men_n473_), .C(men_men_n468_), .Y(men_men_n488_));
  NA2        u0460(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n489_));
  NOi21      u0461(.An(d), .B(e), .Y(men_men_n490_));
  NO2        u0462(.A(men_men_n185_), .B(men_men_n55_), .Y(men_men_n491_));
  NAi31      u0463(.An(j), .B(l), .C(i), .Y(men_men_n492_));
  OAI210     u0464(.A0(men_men_n492_), .A1(men_men_n130_), .B0(men_men_n99_), .Y(men_men_n493_));
  NA3        u0465(.A(men_men_n493_), .B(men_men_n491_), .C(men_men_n490_), .Y(men_men_n494_));
  NO3        u0466(.A(men_men_n390_), .B(men_men_n338_), .C(men_men_n197_), .Y(men_men_n495_));
  NO2        u0467(.A(men_men_n390_), .B(men_men_n366_), .Y(men_men_n496_));
  NO3        u0468(.A(men_men_n496_), .B(men_men_n495_), .C(men_men_n302_), .Y(men_men_n497_));
  NA4        u0469(.A(men_men_n497_), .B(men_men_n494_), .C(men_men_n489_), .D(men_men_n239_), .Y(men_men_n498_));
  AN2        u0470(.A(men_men_n294_), .B(men_men_n188_), .Y(men_men_n499_));
  XO2        u0471(.A(i), .B(h), .Y(men_men_n500_));
  NA3        u0472(.A(men_men_n500_), .B(men_men_n159_), .C(n), .Y(men_men_n501_));
  NAi31      u0473(.An(men_men_n294_), .B(men_men_n501_), .C(men_men_n378_), .Y(men_men_n502_));
  NAi31      u0474(.An(c), .B(f), .C(d), .Y(men_men_n503_));
  AOI210     u0475(.A0(men_men_n274_), .A1(men_men_n191_), .B0(men_men_n503_), .Y(men_men_n504_));
  INV        u0476(.A(men_men_n504_), .Y(men_men_n505_));
  NA3        u0477(.A(men_men_n374_), .B(men_men_n93_), .C(men_men_n92_), .Y(men_men_n506_));
  NA2        u0478(.A(men_men_n223_), .B(men_men_n105_), .Y(men_men_n507_));
  AOI210     u0479(.A0(men_men_n352_), .A1(men_men_n35_), .B0(men_men_n472_), .Y(men_men_n508_));
  NOi21      u0480(.An(men_men_n506_), .B(men_men_n508_), .Y(men_men_n509_));
  AO220      u0481(.A0(men_men_n282_), .A1(men_men_n258_), .B0(men_men_n166_), .B1(men_men_n66_), .Y(men_men_n510_));
  NA3        u0482(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n511_));
  NO2        u0483(.A(men_men_n511_), .B(men_men_n433_), .Y(men_men_n512_));
  NO2        u0484(.A(men_men_n512_), .B(men_men_n290_), .Y(men_men_n513_));
  NAi41      u0485(.An(men_men_n510_), .B(men_men_n513_), .C(men_men_n509_), .D(men_men_n505_), .Y(men_men_n514_));
  NO3        u0486(.A(men_men_n514_), .B(men_men_n499_), .C(men_men_n498_), .Y(men_men_n515_));
  NA4        u0487(.A(men_men_n515_), .B(men_men_n488_), .C(men_men_n456_), .D(men_men_n428_), .Y(men11));
  NO2        u0488(.A(men_men_n71_), .B(f), .Y(men_men_n517_));
  NA2        u0489(.A(j), .B(g), .Y(men_men_n518_));
  NAi31      u0490(.An(i), .B(m), .C(l), .Y(men_men_n519_));
  NA3        u0491(.A(m), .B(k), .C(j), .Y(men_men_n520_));
  NA2        u0492(.A(men_men_n254_), .B(men_men_n110_), .Y(men_men_n521_));
  NA2        u0493(.A(men_men_n46_), .B(j), .Y(men_men_n522_));
  NO2        u0494(.A(men_men_n522_), .B(men_men_n296_), .Y(men_men_n523_));
  NAi31      u0495(.An(d), .B(e), .C(a), .Y(men_men_n524_));
  NO2        u0496(.A(men_men_n524_), .B(n), .Y(men_men_n525_));
  AOI220     u0497(.A0(men_men_n525_), .A1(men_men_n97_), .B0(men_men_n523_), .B1(e), .Y(men_men_n526_));
  NAi41      u0498(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n527_));
  AN2        u0499(.A(men_men_n527_), .B(men_men_n365_), .Y(men_men_n528_));
  AOI210     u0500(.A0(men_men_n528_), .A1(men_men_n390_), .B0(men_men_n267_), .Y(men_men_n529_));
  NA2        u0501(.A(j), .B(i), .Y(men_men_n530_));
  NAi31      u0502(.An(n), .B(m), .C(k), .Y(men_men_n531_));
  NO3        u0503(.A(men_men_n531_), .B(men_men_n530_), .C(men_men_n109_), .Y(men_men_n532_));
  NO4        u0504(.A(n), .B(d), .C(men_men_n113_), .D(a), .Y(men_men_n533_));
  OR2        u0505(.A(n), .B(c), .Y(men_men_n534_));
  NO2        u0506(.A(men_men_n534_), .B(men_men_n149_), .Y(men_men_n535_));
  NO2        u0507(.A(men_men_n535_), .B(men_men_n533_), .Y(men_men_n536_));
  NOi32      u0508(.An(g), .Bn(f), .C(i), .Y(men_men_n537_));
  NA2        u0509(.A(men_men_n537_), .B(men_men_n95_), .Y(men_men_n538_));
  NO2        u0510(.A(men_men_n269_), .B(men_men_n49_), .Y(men_men_n539_));
  NO2        u0511(.A(men_men_n538_), .B(men_men_n536_), .Y(men_men_n540_));
  AOI210     u0512(.A0(men_men_n532_), .A1(men_men_n529_), .B0(men_men_n540_), .Y(men_men_n541_));
  NA2        u0513(.A(men_men_n139_), .B(men_men_n34_), .Y(men_men_n542_));
  OAI220     u0514(.A0(men_men_n542_), .A1(m), .B0(men_men_n522_), .B1(men_men_n229_), .Y(men_men_n543_));
  NOi41      u0515(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n544_));
  NAi32      u0516(.An(e), .Bn(b), .C(c), .Y(men_men_n545_));
  AN2        u0517(.A(men_men_n544_), .B(men_men_n543_), .Y(men_men_n546_));
  OAI220     u0518(.A0(men_men_n392_), .A1(men_men_n391_), .B0(men_men_n519_), .B1(men_men_n518_), .Y(men_men_n547_));
  NAi31      u0519(.An(d), .B(c), .C(a), .Y(men_men_n548_));
  NO2        u0520(.A(men_men_n548_), .B(n), .Y(men_men_n549_));
  NA3        u0521(.A(men_men_n549_), .B(men_men_n547_), .C(e), .Y(men_men_n550_));
  NO3        u0522(.A(men_men_n61_), .B(men_men_n49_), .C(men_men_n211_), .Y(men_men_n551_));
  NO2        u0523(.A(men_men_n226_), .B(men_men_n107_), .Y(men_men_n552_));
  OAI210     u0524(.A0(men_men_n551_), .A1(men_men_n393_), .B0(men_men_n552_), .Y(men_men_n553_));
  NA2        u0525(.A(men_men_n553_), .B(men_men_n550_), .Y(men_men_n554_));
  NO2        u0526(.A(men_men_n271_), .B(n), .Y(men_men_n555_));
  NO2        u0527(.A(men_men_n423_), .B(men_men_n555_), .Y(men_men_n556_));
  NA2        u0528(.A(men_men_n547_), .B(f), .Y(men_men_n557_));
  NAi32      u0529(.An(d), .Bn(a), .C(b), .Y(men_men_n558_));
  NA2        u0530(.A(h), .B(f), .Y(men_men_n559_));
  NO2        u0531(.A(men_men_n559_), .B(men_men_n90_), .Y(men_men_n560_));
  NO2        u0532(.A(men_men_n557_), .B(men_men_n556_), .Y(men_men_n561_));
  NA3        u0533(.A(f), .B(d), .C(b), .Y(men_men_n562_));
  NO3        u0534(.A(men_men_n562_), .B(men_men_n178_), .C(men_men_n175_), .Y(men_men_n563_));
  NO4        u0535(.A(men_men_n563_), .B(men_men_n561_), .C(men_men_n554_), .D(men_men_n546_), .Y(men_men_n564_));
  AN3        u0536(.A(men_men_n564_), .B(men_men_n541_), .C(men_men_n526_), .Y(men_men_n565_));
  INV        u0537(.A(k), .Y(men_men_n566_));
  NA3        u0538(.A(l), .B(men_men_n566_), .C(i), .Y(men_men_n567_));
  INV        u0539(.A(men_men_n567_), .Y(men_men_n568_));
  NA3        u0540(.A(men_men_n389_), .B(men_men_n412_), .C(men_men_n110_), .Y(men_men_n569_));
  NAi32      u0541(.An(h), .Bn(f), .C(g), .Y(men_men_n570_));
  NAi41      u0542(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n571_));
  OAI210     u0543(.A0(men_men_n524_), .A1(n), .B0(men_men_n571_), .Y(men_men_n572_));
  NA2        u0544(.A(men_men_n572_), .B(m), .Y(men_men_n573_));
  NAi31      u0545(.An(h), .B(g), .C(f), .Y(men_men_n574_));
  OR3        u0546(.A(men_men_n574_), .B(men_men_n271_), .C(men_men_n49_), .Y(men_men_n575_));
  NA4        u0547(.A(men_men_n412_), .B(men_men_n118_), .C(men_men_n110_), .D(e), .Y(men_men_n576_));
  AN2        u0548(.A(men_men_n576_), .B(men_men_n575_), .Y(men_men_n577_));
  OA210      u0549(.A0(men_men_n573_), .A1(men_men_n570_), .B0(men_men_n577_), .Y(men_men_n578_));
  NO4        u0550(.A(men_men_n574_), .B(men_men_n534_), .C(men_men_n149_), .D(men_men_n73_), .Y(men_men_n579_));
  NAi31      u0551(.An(men_men_n579_), .B(men_men_n578_), .C(men_men_n569_), .Y(men_men_n580_));
  NAi31      u0552(.An(f), .B(h), .C(g), .Y(men_men_n581_));
  NO4        u0553(.A(men_men_n306_), .B(men_men_n581_), .C(men_men_n71_), .D(men_men_n73_), .Y(men_men_n582_));
  NOi32      u0554(.An(b), .Bn(a), .C(c), .Y(men_men_n583_));
  NOi41      u0555(.An(men_men_n583_), .B(men_men_n347_), .C(men_men_n68_), .D(men_men_n114_), .Y(men_men_n584_));
  OR2        u0556(.A(men_men_n584_), .B(men_men_n582_), .Y(men_men_n585_));
  NOi32      u0557(.An(d), .Bn(a), .C(e), .Y(men_men_n586_));
  NA2        u0558(.A(men_men_n586_), .B(men_men_n110_), .Y(men_men_n587_));
  NO2        u0559(.A(n), .B(c), .Y(men_men_n588_));
  NA3        u0560(.A(men_men_n588_), .B(men_men_n29_), .C(m), .Y(men_men_n589_));
  NAi32      u0561(.An(n), .Bn(f), .C(m), .Y(men_men_n590_));
  NA3        u0562(.A(men_men_n590_), .B(men_men_n589_), .C(men_men_n587_), .Y(men_men_n591_));
  NOi32      u0563(.An(e), .Bn(a), .C(d), .Y(men_men_n592_));
  AOI210     u0564(.A0(men_men_n29_), .A1(d), .B0(men_men_n592_), .Y(men_men_n593_));
  AOI210     u0565(.A0(men_men_n593_), .A1(men_men_n210_), .B0(men_men_n542_), .Y(men_men_n594_));
  AOI210     u0566(.A0(men_men_n594_), .A1(men_men_n591_), .B0(men_men_n585_), .Y(men_men_n595_));
  OAI210     u0567(.A0(men_men_n244_), .A1(men_men_n82_), .B0(men_men_n595_), .Y(men_men_n596_));
  AOI210     u0568(.A0(men_men_n580_), .A1(men_men_n568_), .B0(men_men_n596_), .Y(men_men_n597_));
  NO3        u0569(.A(men_men_n313_), .B(men_men_n60_), .C(n), .Y(men_men_n598_));
  NA3        u0570(.A(men_men_n503_), .B(men_men_n173_), .C(men_men_n172_), .Y(men_men_n599_));
  NA2        u0571(.A(men_men_n454_), .B(men_men_n226_), .Y(men_men_n600_));
  OR2        u0572(.A(men_men_n600_), .B(men_men_n599_), .Y(men_men_n601_));
  NA2        u0573(.A(men_men_n74_), .B(men_men_n110_), .Y(men_men_n602_));
  NO2        u0574(.A(men_men_n602_), .B(men_men_n45_), .Y(men_men_n603_));
  AOI220     u0575(.A0(men_men_n603_), .A1(men_men_n529_), .B0(men_men_n601_), .B1(men_men_n598_), .Y(men_men_n604_));
  NO2        u0576(.A(men_men_n604_), .B(men_men_n82_), .Y(men_men_n605_));
  NOi32      u0577(.An(e), .Bn(c), .C(f), .Y(men_men_n606_));
  NOi21      u0578(.An(f), .B(g), .Y(men_men_n607_));
  NO2        u0579(.A(men_men_n607_), .B(men_men_n208_), .Y(men_men_n608_));
  NA2        u0580(.A(men_men_n606_), .B(men_men_n177_), .Y(men_men_n609_));
  NA2        u0581(.A(men_men_n609_), .B(men_men_n180_), .Y(men_men_n610_));
  AOI210     u0582(.A0(men_men_n528_), .A1(men_men_n390_), .B0(men_men_n295_), .Y(men_men_n611_));
  NA2        u0583(.A(men_men_n611_), .B(men_men_n259_), .Y(men_men_n612_));
  NOi21      u0584(.An(j), .B(l), .Y(men_men_n613_));
  NO2        u0585(.A(k), .B(men_men_n257_), .Y(men_men_n614_));
  NA2        u0586(.A(men_men_n614_), .B(men_men_n613_), .Y(men_men_n615_));
  NOi31      u0587(.An(m), .B(n), .C(k), .Y(men_men_n616_));
  NA2        u0588(.A(men_men_n613_), .B(men_men_n616_), .Y(men_men_n617_));
  AOI210     u0589(.A0(men_men_n390_), .A1(men_men_n365_), .B0(men_men_n295_), .Y(men_men_n618_));
  NAi21      u0590(.An(men_men_n617_), .B(men_men_n618_), .Y(men_men_n619_));
  NO2        u0591(.A(men_men_n271_), .B(men_men_n49_), .Y(men_men_n620_));
  NO2        u0592(.A(men_men_n306_), .B(men_men_n581_), .Y(men_men_n621_));
  NO2        u0593(.A(men_men_n524_), .B(men_men_n49_), .Y(men_men_n622_));
  AOI220     u0594(.A0(men_men_n622_), .A1(men_men_n621_), .B0(men_men_n620_), .B1(men_men_n560_), .Y(men_men_n623_));
  NA3        u0595(.A(men_men_n623_), .B(men_men_n619_), .C(men_men_n612_), .Y(men_men_n624_));
  NA2        u0596(.A(men_men_n105_), .B(men_men_n36_), .Y(men_men_n625_));
  NO2        u0597(.A(k), .B(men_men_n211_), .Y(men_men_n626_));
  INV        u0598(.A(men_men_n354_), .Y(men_men_n627_));
  NO2        u0599(.A(men_men_n627_), .B(n), .Y(men_men_n628_));
  NAi31      u0600(.An(men_men_n625_), .B(men_men_n628_), .C(men_men_n626_), .Y(men_men_n629_));
  AN3        u0601(.A(f), .B(d), .C(b), .Y(men_men_n630_));
  NAi31      u0602(.An(m), .B(n), .C(k), .Y(men_men_n631_));
  OR2        u0603(.A(men_men_n133_), .B(men_men_n60_), .Y(men_men_n632_));
  OAI210     u0604(.A0(men_men_n632_), .A1(men_men_n631_), .B0(men_men_n246_), .Y(men_men_n633_));
  NA2        u0605(.A(men_men_n633_), .B(j), .Y(men_men_n634_));
  NA2        u0606(.A(men_men_n634_), .B(men_men_n629_), .Y(men_men_n635_));
  NO4        u0607(.A(men_men_n635_), .B(men_men_n624_), .C(men_men_n610_), .D(men_men_n605_), .Y(men_men_n636_));
  NA2        u0608(.A(men_men_n374_), .B(men_men_n162_), .Y(men_men_n637_));
  NAi31      u0609(.An(g), .B(h), .C(f), .Y(men_men_n638_));
  OR3        u0610(.A(men_men_n638_), .B(men_men_n271_), .C(n), .Y(men_men_n639_));
  OA210      u0611(.A0(men_men_n524_), .A1(n), .B0(men_men_n571_), .Y(men_men_n640_));
  NO2        u0612(.A(men_men_n640_), .B(men_men_n86_), .Y(men_men_n641_));
  NOi21      u0613(.An(men_men_n639_), .B(men_men_n641_), .Y(men_men_n642_));
  AOI210     u0614(.A0(men_men_n642_), .A1(men_men_n637_), .B0(men_men_n520_), .Y(men_men_n643_));
  NO3        u0615(.A(g), .B(men_men_n210_), .C(men_men_n55_), .Y(men_men_n644_));
  NAi21      u0616(.An(h), .B(j), .Y(men_men_n645_));
  NO2        u0617(.A(men_men_n507_), .B(men_men_n82_), .Y(men_men_n646_));
  OAI210     u0618(.A0(men_men_n646_), .A1(men_men_n386_), .B0(men_men_n644_), .Y(men_men_n647_));
  OR2        u0619(.A(men_men_n71_), .B(men_men_n73_), .Y(men_men_n648_));
  NA2        u0620(.A(men_men_n583_), .B(men_men_n336_), .Y(men_men_n649_));
  OA220      u0621(.A0(men_men_n617_), .A1(men_men_n649_), .B0(men_men_n615_), .B1(men_men_n648_), .Y(men_men_n650_));
  NA2        u0622(.A(h), .B(men_men_n37_), .Y(men_men_n651_));
  NA2        u0623(.A(men_men_n95_), .B(men_men_n46_), .Y(men_men_n652_));
  NO2        u0624(.A(men_men_n652_), .B(men_men_n329_), .Y(men_men_n653_));
  AOI210     u0625(.A0(men_men_n558_), .A1(men_men_n422_), .B0(men_men_n49_), .Y(men_men_n654_));
  OAI220     u0626(.A0(men_men_n574_), .A1(men_men_n567_), .B0(men_men_n323_), .B1(men_men_n518_), .Y(men_men_n655_));
  AOI210     u0627(.A0(men_men_n655_), .A1(men_men_n654_), .B0(men_men_n653_), .Y(men_men_n656_));
  NA3        u0628(.A(men_men_n656_), .B(men_men_n650_), .C(men_men_n647_), .Y(men_men_n657_));
  INV        u0629(.A(f), .Y(men_men_n658_));
  NA2        u0630(.A(men_men_n326_), .B(men_men_n139_), .Y(men_men_n659_));
  NA2        u0631(.A(men_men_n354_), .B(men_men_n110_), .Y(men_men_n660_));
  OA220      u0632(.A0(men_men_n660_), .A1(men_men_n542_), .B0(men_men_n352_), .B1(men_men_n108_), .Y(men_men_n661_));
  OAI210     u0633(.A0(men_men_n659_), .A1(men_men_n607_), .B0(men_men_n661_), .Y(men_men_n662_));
  NO3        u0634(.A(men_men_n397_), .B(men_men_n188_), .C(men_men_n187_), .Y(men_men_n663_));
  NA2        u0635(.A(men_men_n663_), .B(men_men_n226_), .Y(men_men_n664_));
  NA3        u0636(.A(men_men_n664_), .B(men_men_n250_), .C(j), .Y(men_men_n665_));
  NO3        u0637(.A(men_men_n454_), .B(men_men_n175_), .C(i), .Y(men_men_n666_));
  NA2        u0638(.A(men_men_n457_), .B(men_men_n79_), .Y(men_men_n667_));
  NO3        u0639(.A(men_men_n520_), .B(men_men_n667_), .C(men_men_n129_), .Y(men_men_n668_));
  INV        u0640(.A(men_men_n668_), .Y(men_men_n669_));
  NA4        u0641(.A(men_men_n669_), .B(men_men_n665_), .C(men_men_n506_), .D(men_men_n395_), .Y(men_men_n670_));
  NO4        u0642(.A(men_men_n670_), .B(men_men_n662_), .C(men_men_n657_), .D(men_men_n643_), .Y(men_men_n671_));
  NA4        u0643(.A(men_men_n671_), .B(men_men_n636_), .C(men_men_n597_), .D(men_men_n565_), .Y(men08));
  NO2        u0644(.A(k), .B(h), .Y(men_men_n673_));
  AO210      u0645(.A0(men_men_n248_), .A1(men_men_n446_), .B0(men_men_n673_), .Y(men_men_n674_));
  NO2        u0646(.A(men_men_n674_), .B(men_men_n293_), .Y(men_men_n675_));
  NA2        u0647(.A(men_men_n606_), .B(men_men_n79_), .Y(men_men_n676_));
  NA2        u0648(.A(men_men_n676_), .B(men_men_n454_), .Y(men_men_n677_));
  AOI210     u0649(.A0(men_men_n677_), .A1(men_men_n675_), .B0(men_men_n485_), .Y(men_men_n678_));
  NA2        u0650(.A(men_men_n79_), .B(men_men_n107_), .Y(men_men_n679_));
  NO2        u0651(.A(men_men_n679_), .B(men_men_n56_), .Y(men_men_n680_));
  NO4        u0652(.A(men_men_n371_), .B(men_men_n109_), .C(j), .D(men_men_n211_), .Y(men_men_n681_));
  NA2        u0653(.A(men_men_n562_), .B(men_men_n228_), .Y(men_men_n682_));
  AOI220     u0654(.A0(men_men_n682_), .A1(men_men_n341_), .B0(men_men_n681_), .B1(men_men_n680_), .Y(men_men_n683_));
  AOI210     u0655(.A0(men_men_n562_), .A1(men_men_n155_), .B0(men_men_n79_), .Y(men_men_n684_));
  NA4        u0656(.A(men_men_n213_), .B(men_men_n139_), .C(men_men_n45_), .D(h), .Y(men_men_n685_));
  AN2        u0657(.A(l), .B(k), .Y(men_men_n686_));
  NA4        u0658(.A(men_men_n686_), .B(men_men_n105_), .C(men_men_n73_), .D(men_men_n211_), .Y(men_men_n687_));
  NA3        u0659(.A(men_men_n683_), .B(men_men_n678_), .C(men_men_n343_), .Y(men_men_n688_));
  AN2        u0660(.A(men_men_n525_), .B(men_men_n91_), .Y(men_men_n689_));
  NO4        u0661(.A(men_men_n175_), .B(men_men_n385_), .C(men_men_n109_), .D(g), .Y(men_men_n690_));
  AOI210     u0662(.A0(men_men_n690_), .A1(men_men_n682_), .B0(men_men_n512_), .Y(men_men_n691_));
  NO2        u0663(.A(men_men_n38_), .B(men_men_n210_), .Y(men_men_n692_));
  NA2        u0664(.A(men_men_n692_), .B(men_men_n555_), .Y(men_men_n693_));
  NAi31      u0665(.An(men_men_n689_), .B(men_men_n693_), .C(men_men_n691_), .Y(men_men_n694_));
  NO2        u0666(.A(men_men_n528_), .B(men_men_n35_), .Y(men_men_n695_));
  OAI210     u0667(.A0(men_men_n545_), .A1(men_men_n47_), .B0(men_men_n632_), .Y(men_men_n696_));
  NO2        u0668(.A(men_men_n477_), .B(men_men_n130_), .Y(men_men_n697_));
  AOI210     u0669(.A0(men_men_n697_), .A1(men_men_n696_), .B0(men_men_n695_), .Y(men_men_n698_));
  NO3        u0670(.A(men_men_n313_), .B(men_men_n129_), .C(men_men_n41_), .Y(men_men_n699_));
  NAi21      u0671(.An(men_men_n699_), .B(men_men_n687_), .Y(men_men_n700_));
  NA2        u0672(.A(men_men_n674_), .B(men_men_n134_), .Y(men_men_n701_));
  AOI220     u0673(.A0(men_men_n701_), .A1(men_men_n396_), .B0(men_men_n700_), .B1(men_men_n75_), .Y(men_men_n702_));
  OAI210     u0674(.A0(men_men_n698_), .A1(men_men_n82_), .B0(men_men_n702_), .Y(men_men_n703_));
  NA2        u0675(.A(men_men_n354_), .B(men_men_n43_), .Y(men_men_n704_));
  NA3        u0676(.A(men_men_n664_), .B(men_men_n330_), .C(men_men_n377_), .Y(men_men_n705_));
  NA2        u0677(.A(men_men_n686_), .B(men_men_n216_), .Y(men_men_n706_));
  NO2        u0678(.A(men_men_n706_), .B(men_men_n325_), .Y(men_men_n707_));
  AOI210     u0679(.A0(men_men_n707_), .A1(men_men_n658_), .B0(men_men_n484_), .Y(men_men_n708_));
  NA3        u0680(.A(m), .B(l), .C(k), .Y(men_men_n709_));
  NO2        u0681(.A(men_men_n639_), .B(men_men_n709_), .Y(men_men_n710_));
  NO2        u0682(.A(men_men_n527_), .B(men_men_n267_), .Y(men_men_n711_));
  NOi21      u0683(.An(men_men_n711_), .B(men_men_n521_), .Y(men_men_n712_));
  NA4        u0684(.A(men_men_n110_), .B(l), .C(k), .D(men_men_n82_), .Y(men_men_n713_));
  NA3        u0685(.A(men_men_n118_), .B(men_men_n405_), .C(i), .Y(men_men_n714_));
  NO2        u0686(.A(men_men_n714_), .B(men_men_n713_), .Y(men_men_n715_));
  NO3        u0687(.A(men_men_n715_), .B(men_men_n712_), .C(men_men_n710_), .Y(men_men_n716_));
  NA4        u0688(.A(men_men_n716_), .B(men_men_n708_), .C(men_men_n705_), .D(men_men_n704_), .Y(men_men_n717_));
  NO4        u0689(.A(men_men_n717_), .B(men_men_n703_), .C(men_men_n694_), .D(men_men_n688_), .Y(men_men_n718_));
  NA2        u0690(.A(men_men_n608_), .B(men_men_n386_), .Y(men_men_n719_));
  NOi31      u0691(.An(g), .B(h), .C(f), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n622_), .B(men_men_n720_), .Y(men_men_n721_));
  AO210      u0693(.A0(men_men_n721_), .A1(men_men_n575_), .B0(men_men_n530_), .Y(men_men_n722_));
  NO3        u0694(.A(men_men_n390_), .B(men_men_n518_), .C(h), .Y(men_men_n723_));
  AOI210     u0695(.A0(men_men_n723_), .A1(men_men_n110_), .B0(men_men_n496_), .Y(men_men_n724_));
  NA4        u0696(.A(men_men_n724_), .B(men_men_n722_), .C(men_men_n719_), .D(men_men_n247_), .Y(men_men_n725_));
  NA2        u0697(.A(men_men_n686_), .B(men_men_n73_), .Y(men_men_n726_));
  NO4        u0698(.A(men_men_n663_), .B(men_men_n175_), .C(n), .D(i), .Y(men_men_n727_));
  NOi21      u0699(.An(h), .B(j), .Y(men_men_n728_));
  NA2        u0700(.A(men_men_n728_), .B(f), .Y(men_men_n729_));
  NO2        u0701(.A(men_men_n729_), .B(men_men_n241_), .Y(men_men_n730_));
  NO3        u0702(.A(men_men_n730_), .B(men_men_n727_), .C(men_men_n666_), .Y(men_men_n731_));
  OAI220     u0703(.A0(men_men_n731_), .A1(men_men_n726_), .B0(men_men_n577_), .B1(men_men_n61_), .Y(men_men_n732_));
  AOI210     u0704(.A0(men_men_n725_), .A1(l), .B0(men_men_n732_), .Y(men_men_n733_));
  NO2        u0705(.A(j), .B(i), .Y(men_men_n734_));
  NA3        u0706(.A(men_men_n734_), .B(men_men_n77_), .C(l), .Y(men_men_n735_));
  NA2        u0707(.A(men_men_n734_), .B(men_men_n33_), .Y(men_men_n736_));
  NA2        u0708(.A(men_men_n415_), .B(men_men_n118_), .Y(men_men_n737_));
  OA220      u0709(.A0(men_men_n737_), .A1(men_men_n736_), .B0(men_men_n735_), .B1(men_men_n573_), .Y(men_men_n738_));
  NO3        u0710(.A(men_men_n150_), .B(men_men_n49_), .C(men_men_n107_), .Y(men_men_n739_));
  NO3        u0711(.A(men_men_n534_), .B(men_men_n149_), .C(men_men_n73_), .Y(men_men_n740_));
  NO3        u0712(.A(men_men_n477_), .B(men_men_n434_), .C(j), .Y(men_men_n741_));
  OAI210     u0713(.A0(men_men_n740_), .A1(men_men_n739_), .B0(men_men_n741_), .Y(men_men_n742_));
  OAI210     u0714(.A0(men_men_n721_), .A1(men_men_n61_), .B0(men_men_n742_), .Y(men_men_n743_));
  NA2        u0715(.A(k), .B(j), .Y(men_men_n744_));
  NO3        u0716(.A(men_men_n293_), .B(men_men_n744_), .C(men_men_n40_), .Y(men_men_n745_));
  AN3        u0717(.A(men_men_n1451_), .B(men_men_n745_), .C(men_men_n94_), .Y(men_men_n746_));
  NO3        u0718(.A(men_men_n175_), .B(men_men_n385_), .C(men_men_n109_), .Y(men_men_n747_));
  AOI220     u0719(.A0(men_men_n747_), .A1(men_men_n242_), .B0(men_men_n600_), .B1(men_men_n304_), .Y(men_men_n748_));
  NAi31      u0720(.An(men_men_n593_), .B(men_men_n88_), .C(men_men_n79_), .Y(men_men_n749_));
  NA2        u0721(.A(men_men_n749_), .B(men_men_n748_), .Y(men_men_n750_));
  NO2        u0722(.A(men_men_n293_), .B(men_men_n134_), .Y(men_men_n751_));
  AOI220     u0723(.A0(men_men_n751_), .A1(men_men_n608_), .B0(men_men_n699_), .B1(men_men_n684_), .Y(men_men_n752_));
  NO2        u0724(.A(men_men_n709_), .B(men_men_n86_), .Y(men_men_n753_));
  NA2        u0725(.A(men_men_n753_), .B(men_men_n572_), .Y(men_men_n754_));
  NO2        u0726(.A(men_men_n574_), .B(men_men_n114_), .Y(men_men_n755_));
  OAI210     u0727(.A0(men_men_n755_), .A1(men_men_n741_), .B0(men_men_n654_), .Y(men_men_n756_));
  NA3        u0728(.A(men_men_n756_), .B(men_men_n754_), .C(men_men_n752_), .Y(men_men_n757_));
  OR4        u0729(.A(men_men_n757_), .B(men_men_n750_), .C(men_men_n746_), .D(men_men_n743_), .Y(men_men_n758_));
  NO4        u0730(.A(men_men_n477_), .B(men_men_n429_), .C(j), .D(f), .Y(men_men_n759_));
  OAI220     u0731(.A0(men_men_n685_), .A1(men_men_n676_), .B0(men_men_n329_), .B1(men_men_n38_), .Y(men_men_n760_));
  AOI210     u0732(.A0(men_men_n759_), .A1(men_men_n253_), .B0(men_men_n760_), .Y(men_men_n761_));
  NA3        u0733(.A(men_men_n537_), .B(men_men_n286_), .C(h), .Y(men_men_n762_));
  NOi21      u0734(.An(men_men_n654_), .B(men_men_n762_), .Y(men_men_n763_));
  NO2        u0735(.A(men_men_n87_), .B(men_men_n47_), .Y(men_men_n764_));
  OAI220     u0736(.A0(men_men_n762_), .A1(men_men_n589_), .B0(men_men_n735_), .B1(men_men_n648_), .Y(men_men_n765_));
  AOI210     u0737(.A0(men_men_n764_), .A1(men_men_n628_), .B0(men_men_n765_), .Y(men_men_n766_));
  NAi31      u0738(.An(men_men_n763_), .B(men_men_n766_), .C(men_men_n761_), .Y(men_men_n767_));
  BUFFER     u0739(.A(men_men_n91_), .Y(men_men_n768_));
  AOI220     u0740(.A0(men_men_n768_), .A1(men_men_n234_), .B0(men_men_n741_), .B1(men_men_n620_), .Y(men_men_n769_));
  NO2        u0741(.A(men_men_n640_), .B(men_men_n73_), .Y(men_men_n770_));
  AOI210     u0742(.A0(men_men_n759_), .A1(men_men_n770_), .B0(men_men_n332_), .Y(men_men_n771_));
  AOI220     u0743(.A0(men_men_n588_), .A1(men_men_n29_), .B0(men_men_n457_), .B1(men_men_n79_), .Y(men_men_n772_));
  NO2        u0744(.A(men_men_n762_), .B(men_men_n483_), .Y(men_men_n773_));
  INV        u0745(.A(men_men_n773_), .Y(men_men_n774_));
  NA3        u0746(.A(men_men_n774_), .B(men_men_n771_), .C(men_men_n769_), .Y(men_men_n775_));
  NOi41      u0747(.An(men_men_n738_), .B(men_men_n775_), .C(men_men_n767_), .D(men_men_n758_), .Y(men_men_n776_));
  OR3        u0748(.A(men_men_n685_), .B(men_men_n228_), .C(g), .Y(men_men_n777_));
  NA2        u0749(.A(men_men_n46_), .B(men_men_n55_), .Y(men_men_n778_));
  NO3        u0750(.A(men_men_n778_), .B(men_men_n736_), .C(men_men_n271_), .Y(men_men_n779_));
  NO3        u0751(.A(men_men_n518_), .B(men_men_n89_), .C(h), .Y(men_men_n780_));
  AOI210     u0752(.A0(men_men_n780_), .A1(men_men_n680_), .B0(men_men_n779_), .Y(men_men_n781_));
  NA3        u0753(.A(men_men_n781_), .B(men_men_n777_), .C(men_men_n398_), .Y(men_men_n782_));
  OR2        u0754(.A(men_men_n638_), .B(men_men_n87_), .Y(men_men_n783_));
  NOi31      u0755(.An(b), .B(d), .C(a), .Y(men_men_n784_));
  NO2        u0756(.A(men_men_n784_), .B(men_men_n586_), .Y(men_men_n785_));
  NO2        u0757(.A(men_men_n785_), .B(n), .Y(men_men_n786_));
  NOi21      u0758(.An(men_men_n772_), .B(men_men_n786_), .Y(men_men_n787_));
  OAI220     u0759(.A0(men_men_n787_), .A1(men_men_n783_), .B0(men_men_n762_), .B1(men_men_n587_), .Y(men_men_n788_));
  NO3        u0760(.A(men_men_n607_), .B(men_men_n325_), .C(men_men_n114_), .Y(men_men_n789_));
  NOi21      u0761(.An(men_men_n789_), .B(men_men_n160_), .Y(men_men_n790_));
  NO2        u0762(.A(men_men_n663_), .B(n), .Y(men_men_n791_));
  AOI220     u0763(.A0(men_men_n751_), .A1(men_men_n644_), .B0(men_men_n791_), .B1(men_men_n675_), .Y(men_men_n792_));
  NO2        u0764(.A(men_men_n320_), .B(men_men_n233_), .Y(men_men_n793_));
  OAI210     u0765(.A0(men_men_n91_), .A1(men_men_n88_), .B0(men_men_n793_), .Y(men_men_n794_));
  NA2        u0766(.A(men_men_n118_), .B(men_men_n79_), .Y(men_men_n795_));
  AOI210     u0767(.A0(men_men_n419_), .A1(men_men_n411_), .B0(men_men_n795_), .Y(men_men_n796_));
  NAi21      u0768(.An(men_men_n796_), .B(men_men_n794_), .Y(men_men_n797_));
  NA2        u0769(.A(men_men_n707_), .B(men_men_n34_), .Y(men_men_n798_));
  NAi21      u0770(.An(men_men_n713_), .B(men_men_n430_), .Y(men_men_n799_));
  NO2        u0771(.A(men_men_n267_), .B(i), .Y(men_men_n800_));
  NA2        u0772(.A(men_men_n690_), .B(men_men_n342_), .Y(men_men_n801_));
  NA2        u0773(.A(men_men_n579_), .B(men_men_n355_), .Y(men_men_n802_));
  AN3        u0774(.A(men_men_n802_), .B(men_men_n801_), .C(men_men_n799_), .Y(men_men_n803_));
  NAi41      u0775(.An(men_men_n797_), .B(men_men_n803_), .C(men_men_n798_), .D(men_men_n792_), .Y(men_men_n804_));
  NO4        u0776(.A(men_men_n804_), .B(men_men_n790_), .C(men_men_n788_), .D(men_men_n782_), .Y(men_men_n805_));
  NA4        u0777(.A(men_men_n805_), .B(men_men_n776_), .C(men_men_n733_), .D(men_men_n718_), .Y(men09));
  INV        u0778(.A(men_men_n119_), .Y(men_men_n807_));
  NA2        u0779(.A(f), .B(e), .Y(men_men_n808_));
  NO2        u0780(.A(men_men_n221_), .B(men_men_n109_), .Y(men_men_n809_));
  NA2        u0781(.A(men_men_n809_), .B(g), .Y(men_men_n810_));
  NA4        u0782(.A(men_men_n306_), .B(men_men_n466_), .C(men_men_n255_), .D(men_men_n116_), .Y(men_men_n811_));
  AOI210     u0783(.A0(men_men_n811_), .A1(g), .B0(men_men_n463_), .Y(men_men_n812_));
  AOI210     u0784(.A0(men_men_n812_), .A1(men_men_n810_), .B0(men_men_n808_), .Y(men_men_n813_));
  NA2        u0785(.A(men_men_n440_), .B(e), .Y(men_men_n814_));
  NO2        u0786(.A(men_men_n814_), .B(men_men_n503_), .Y(men_men_n815_));
  AOI210     u0787(.A0(men_men_n813_), .A1(men_men_n807_), .B0(men_men_n815_), .Y(men_men_n816_));
  NO2        u0788(.A(men_men_n200_), .B(men_men_n210_), .Y(men_men_n817_));
  NA3        u0789(.A(m), .B(l), .C(i), .Y(men_men_n818_));
  OAI220     u0790(.A0(men_men_n574_), .A1(men_men_n818_), .B0(men_men_n347_), .B1(men_men_n519_), .Y(men_men_n819_));
  NA4        u0791(.A(men_men_n83_), .B(men_men_n82_), .C(g), .D(f), .Y(men_men_n820_));
  NAi31      u0792(.An(men_men_n819_), .B(men_men_n820_), .C(men_men_n435_), .Y(men_men_n821_));
  OR2        u0793(.A(men_men_n821_), .B(men_men_n817_), .Y(men_men_n822_));
  NA3        u0794(.A(men_men_n783_), .B(men_men_n557_), .C(men_men_n511_), .Y(men_men_n823_));
  OA210      u0795(.A0(men_men_n823_), .A1(men_men_n822_), .B0(men_men_n786_), .Y(men_men_n824_));
  INV        u0796(.A(men_men_n334_), .Y(men_men_n825_));
  NO2        u0797(.A(men_men_n125_), .B(men_men_n123_), .Y(men_men_n826_));
  INV        u0798(.A(men_men_n329_), .Y(men_men_n827_));
  NA2        u0799(.A(men_men_n336_), .B(men_men_n337_), .Y(men_men_n828_));
  NA3        u0800(.A(men_men_n111_), .B(men_men_n186_), .C(men_men_n31_), .Y(men_men_n829_));
  NA2        u0801(.A(men_men_n829_), .B(men_men_n609_), .Y(men_men_n830_));
  NO2        u0802(.A(men_men_n570_), .B(men_men_n492_), .Y(men_men_n831_));
  NOi21      u0803(.An(f), .B(d), .Y(men_men_n832_));
  NA2        u0804(.A(men_men_n832_), .B(m), .Y(men_men_n833_));
  NO2        u0805(.A(men_men_n833_), .B(men_men_n51_), .Y(men_men_n834_));
  NOi32      u0806(.An(g), .Bn(f), .C(d), .Y(men_men_n835_));
  NA4        u0807(.A(men_men_n835_), .B(men_men_n588_), .C(men_men_n29_), .D(m), .Y(men_men_n836_));
  NOi21      u0808(.An(men_men_n307_), .B(men_men_n836_), .Y(men_men_n837_));
  AOI210     u0809(.A0(men_men_n834_), .A1(men_men_n535_), .B0(men_men_n837_), .Y(men_men_n838_));
  NA3        u0810(.A(men_men_n306_), .B(men_men_n255_), .C(men_men_n116_), .Y(men_men_n839_));
  AN2        u0811(.A(f), .B(d), .Y(men_men_n840_));
  NA3        u0812(.A(men_men_n470_), .B(men_men_n840_), .C(men_men_n79_), .Y(men_men_n841_));
  NO3        u0813(.A(men_men_n841_), .B(men_men_n73_), .C(men_men_n211_), .Y(men_men_n842_));
  NA2        u0814(.A(men_men_n839_), .B(men_men_n842_), .Y(men_men_n843_));
  NAi31      u0815(.An(men_men_n482_), .B(men_men_n843_), .C(men_men_n838_), .Y(men_men_n844_));
  NO2        u0816(.A(men_men_n631_), .B(men_men_n325_), .Y(men_men_n845_));
  INV        u0817(.A(men_men_n230_), .Y(men_men_n846_));
  NA2        u0818(.A(men_men_n586_), .B(men_men_n79_), .Y(men_men_n847_));
  NO2        u0819(.A(men_men_n828_), .B(men_men_n847_), .Y(men_men_n848_));
  NA3        u0820(.A(men_men_n159_), .B(men_men_n105_), .C(men_men_n104_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n334_), .B(men_men_n849_), .Y(men_men_n850_));
  NOi41      u0822(.An(men_men_n219_), .B(men_men_n850_), .C(men_men_n848_), .D(men_men_n302_), .Y(men_men_n851_));
  NA2        u0823(.A(c), .B(men_men_n113_), .Y(men_men_n852_));
  NO2        u0824(.A(men_men_n852_), .B(men_men_n402_), .Y(men_men_n853_));
  NA3        u0825(.A(men_men_n853_), .B(men_men_n502_), .C(f), .Y(men_men_n854_));
  OR2        u0826(.A(men_men_n638_), .B(men_men_n531_), .Y(men_men_n855_));
  INV        u0827(.A(men_men_n855_), .Y(men_men_n856_));
  NA2        u0828(.A(men_men_n785_), .B(men_men_n108_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n857_), .B(men_men_n856_), .Y(men_men_n858_));
  NA4        u0830(.A(men_men_n858_), .B(men_men_n854_), .C(men_men_n851_), .D(men_men_n846_), .Y(men_men_n859_));
  NO4        u0831(.A(men_men_n859_), .B(men_men_n844_), .C(men_men_n830_), .D(men_men_n824_), .Y(men_men_n860_));
  OR2        u0832(.A(men_men_n841_), .B(men_men_n73_), .Y(men_men_n861_));
  NA2        u0833(.A(men_men_n809_), .B(g), .Y(men_men_n862_));
  AOI210     u0834(.A0(men_men_n862_), .A1(men_men_n287_), .B0(men_men_n861_), .Y(men_men_n863_));
  NO2        u0835(.A(men_men_n329_), .B(men_men_n820_), .Y(men_men_n864_));
  NO2        u0836(.A(men_men_n134_), .B(men_men_n130_), .Y(men_men_n865_));
  NO2        u0837(.A(men_men_n226_), .B(men_men_n220_), .Y(men_men_n866_));
  AOI220     u0838(.A0(men_men_n866_), .A1(men_men_n223_), .B0(men_men_n300_), .B1(men_men_n865_), .Y(men_men_n867_));
  NA2        u0839(.A(e), .B(d), .Y(men_men_n868_));
  OAI220     u0840(.A0(men_men_n868_), .A1(c), .B0(men_men_n320_), .B1(d), .Y(men_men_n869_));
  NA3        u0841(.A(men_men_n869_), .B(men_men_n449_), .C(men_men_n500_), .Y(men_men_n870_));
  NO2        u0842(.A(men_men_n507_), .B(men_men_n226_), .Y(men_men_n871_));
  INV        u0843(.A(men_men_n871_), .Y(men_men_n872_));
  NA2        u0844(.A(men_men_n279_), .B(men_men_n165_), .Y(men_men_n873_));
  NA2        u0845(.A(men_men_n842_), .B(men_men_n873_), .Y(men_men_n874_));
  NA3        u0846(.A(men_men_n168_), .B(men_men_n80_), .C(men_men_n34_), .Y(men_men_n875_));
  NA4        u0847(.A(men_men_n875_), .B(men_men_n874_), .C(men_men_n872_), .D(men_men_n870_), .Y(men_men_n876_));
  NO4        u0848(.A(men_men_n876_), .B(men_men_n1450_), .C(men_men_n864_), .D(men_men_n863_), .Y(men_men_n877_));
  NA2        u0849(.A(men_men_n825_), .B(men_men_n31_), .Y(men_men_n878_));
  AO210      u0850(.A0(men_men_n878_), .A1(men_men_n676_), .B0(men_men_n214_), .Y(men_men_n879_));
  OAI220     u0851(.A0(men_men_n607_), .A1(men_men_n60_), .B0(men_men_n295_), .B1(j), .Y(men_men_n880_));
  AOI220     u0852(.A0(men_men_n880_), .A1(men_men_n845_), .B0(men_men_n598_), .B1(men_men_n606_), .Y(men_men_n881_));
  OAI210     u0853(.A0(men_men_n814_), .A1(men_men_n172_), .B0(men_men_n881_), .Y(men_men_n882_));
  OAI210     u0854(.A0(men_men_n809_), .A1(men_men_n873_), .B0(men_men_n835_), .Y(men_men_n883_));
  NO2        u0855(.A(men_men_n883_), .B(men_men_n589_), .Y(men_men_n884_));
  AOI210     u0856(.A0(men_men_n115_), .A1(men_men_n114_), .B0(men_men_n254_), .Y(men_men_n885_));
  NO2        u0857(.A(men_men_n885_), .B(men_men_n836_), .Y(men_men_n886_));
  AO210      u0858(.A0(men_men_n827_), .A1(men_men_n819_), .B0(men_men_n886_), .Y(men_men_n887_));
  NOi31      u0859(.An(men_men_n535_), .B(men_men_n833_), .C(men_men_n287_), .Y(men_men_n888_));
  NO4        u0860(.A(men_men_n888_), .B(men_men_n887_), .C(men_men_n884_), .D(men_men_n882_), .Y(men_men_n889_));
  AO220      u0861(.A0(men_men_n449_), .A1(men_men_n728_), .B0(men_men_n177_), .B1(f), .Y(men_men_n890_));
  OAI210     u0862(.A0(men_men_n890_), .A1(men_men_n452_), .B0(men_men_n869_), .Y(men_men_n891_));
  NO2        u0863(.A(men_men_n434_), .B(men_men_n70_), .Y(men_men_n892_));
  OAI210     u0864(.A0(men_men_n823_), .A1(men_men_n892_), .B0(men_men_n680_), .Y(men_men_n893_));
  AN4        u0865(.A(men_men_n893_), .B(men_men_n891_), .C(men_men_n889_), .D(men_men_n879_), .Y(men_men_n894_));
  NA4        u0866(.A(men_men_n894_), .B(men_men_n877_), .C(men_men_n860_), .D(men_men_n816_), .Y(men12));
  NO2        u0867(.A(men_men_n447_), .B(c), .Y(men_men_n896_));
  NO4        u0868(.A(men_men_n439_), .B(men_men_n248_), .C(men_men_n566_), .D(men_men_n211_), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n897_), .B(men_men_n896_), .Y(men_men_n898_));
  NA2        u0870(.A(men_men_n535_), .B(men_men_n892_), .Y(men_men_n899_));
  NO2        u0871(.A(men_men_n447_), .B(men_men_n113_), .Y(men_men_n900_));
  NO2        u0872(.A(men_men_n826_), .B(men_men_n347_), .Y(men_men_n901_));
  NO2        u0873(.A(men_men_n638_), .B(men_men_n371_), .Y(men_men_n902_));
  AOI220     u0874(.A0(men_men_n902_), .A1(men_men_n533_), .B0(men_men_n901_), .B1(men_men_n900_), .Y(men_men_n903_));
  NA4        u0875(.A(men_men_n903_), .B(men_men_n899_), .C(men_men_n898_), .D(men_men_n438_), .Y(men_men_n904_));
  AOI210     u0876(.A0(men_men_n229_), .A1(men_men_n333_), .B0(men_men_n197_), .Y(men_men_n905_));
  BUFFER     u0877(.A(men_men_n905_), .Y(men_men_n906_));
  AOI210     u0878(.A0(men_men_n331_), .A1(men_men_n383_), .B0(men_men_n211_), .Y(men_men_n907_));
  OAI210     u0879(.A0(men_men_n907_), .A1(men_men_n906_), .B0(men_men_n397_), .Y(men_men_n908_));
  NO2        u0880(.A(men_men_n625_), .B(men_men_n257_), .Y(men_men_n909_));
  NO2        u0881(.A(men_men_n574_), .B(men_men_n818_), .Y(men_men_n910_));
  AOI220     u0882(.A0(men_men_n910_), .A1(men_men_n555_), .B0(men_men_n793_), .B1(men_men_n909_), .Y(men_men_n911_));
  NO2        u0883(.A(men_men_n150_), .B(men_men_n233_), .Y(men_men_n912_));
  NA3        u0884(.A(men_men_n912_), .B(men_men_n236_), .C(i), .Y(men_men_n913_));
  NA3        u0885(.A(men_men_n913_), .B(men_men_n911_), .C(men_men_n908_), .Y(men_men_n914_));
  NA4        u0886(.A(men_men_n440_), .B(men_men_n432_), .C(men_men_n182_), .D(g), .Y(men_men_n915_));
  INV        u0887(.A(men_men_n915_), .Y(men_men_n916_));
  NO3        u0888(.A(men_men_n642_), .B(men_men_n87_), .C(men_men_n45_), .Y(men_men_n917_));
  NO4        u0889(.A(men_men_n917_), .B(men_men_n916_), .C(men_men_n914_), .D(men_men_n904_), .Y(men_men_n918_));
  NO2        u0890(.A(men_men_n362_), .B(men_men_n361_), .Y(men_men_n919_));
  NA2        u0891(.A(men_men_n571_), .B(men_men_n71_), .Y(men_men_n920_));
  NA2        u0892(.A(men_men_n920_), .B(men_men_n919_), .Y(men_men_n921_));
  OAI210     u0893(.A0(men_men_n246_), .A1(men_men_n45_), .B0(men_men_n921_), .Y(men_men_n922_));
  NA2        u0894(.A(men_men_n430_), .B(men_men_n259_), .Y(men_men_n923_));
  NO3        u0895(.A(men_men_n795_), .B(men_men_n84_), .C(men_men_n402_), .Y(men_men_n924_));
  NAi31      u0896(.An(men_men_n924_), .B(men_men_n923_), .C(men_men_n317_), .Y(men_men_n925_));
  NO2        u0897(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n926_));
  NA2        u0898(.A(men_men_n616_), .B(men_men_n355_), .Y(men_men_n927_));
  OAI210     u0899(.A0(men_men_n714_), .A1(men_men_n927_), .B0(men_men_n359_), .Y(men_men_n928_));
  NO3        u0900(.A(men_men_n928_), .B(men_men_n925_), .C(men_men_n922_), .Y(men_men_n929_));
  NA2        u0901(.A(men_men_n162_), .B(i), .Y(men_men_n930_));
  NO2        u0902(.A(men_men_n930_), .B(men_men_n87_), .Y(men_men_n931_));
  AOI210     u0903(.A0(men_men_n413_), .A1(men_men_n37_), .B0(men_men_n931_), .Y(men_men_n932_));
  NO2        u0904(.A(men_men_n932_), .B(men_men_n329_), .Y(men_men_n933_));
  NO2        u0905(.A(men_men_n638_), .B(men_men_n492_), .Y(men_men_n934_));
  NA3        u0906(.A(men_men_n336_), .B(men_men_n613_), .C(i), .Y(men_men_n935_));
  OAI210     u0907(.A0(men_men_n434_), .A1(men_men_n306_), .B0(men_men_n935_), .Y(men_men_n936_));
  OAI220     u0908(.A0(men_men_n936_), .A1(men_men_n934_), .B0(men_men_n654_), .B1(men_men_n740_), .Y(men_men_n937_));
  NA2        u0909(.A(men_men_n592_), .B(men_men_n110_), .Y(men_men_n938_));
  OR3        u0910(.A(men_men_n306_), .B(men_men_n429_), .C(f), .Y(men_men_n939_));
  NA3        u0911(.A(men_men_n613_), .B(men_men_n77_), .C(i), .Y(men_men_n940_));
  OA220      u0912(.A0(men_men_n940_), .A1(men_men_n938_), .B0(men_men_n939_), .B1(men_men_n573_), .Y(men_men_n941_));
  NA3        u0913(.A(men_men_n322_), .B(men_men_n115_), .C(g), .Y(men_men_n942_));
  AOI210     u0914(.A0(men_men_n651_), .A1(men_men_n942_), .B0(m), .Y(men_men_n943_));
  OAI210     u0915(.A0(men_men_n943_), .A1(men_men_n901_), .B0(men_men_n321_), .Y(men_men_n944_));
  NA2        u0916(.A(men_men_n667_), .B(men_men_n847_), .Y(men_men_n945_));
  NA2        u0917(.A(men_men_n820_), .B(men_men_n435_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n217_), .B(men_men_n76_), .Y(men_men_n947_));
  NA3        u0919(.A(men_men_n947_), .B(men_men_n940_), .C(men_men_n939_), .Y(men_men_n948_));
  AOI220     u0920(.A0(men_men_n948_), .A1(men_men_n253_), .B0(men_men_n946_), .B1(men_men_n945_), .Y(men_men_n949_));
  NA4        u0921(.A(men_men_n949_), .B(men_men_n944_), .C(men_men_n941_), .D(men_men_n937_), .Y(men_men_n950_));
  NA2        u0922(.A(men_men_n641_), .B(men_men_n83_), .Y(men_men_n951_));
  NA2        u0923(.A(men_men_n572_), .B(men_men_n85_), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n952_), .B(men_men_n951_), .Y(men_men_n953_));
  OAI210     u0925(.A0(men_men_n946_), .A1(men_men_n910_), .B0(men_men_n533_), .Y(men_men_n954_));
  AOI210     u0926(.A0(men_men_n414_), .A1(men_men_n406_), .B0(men_men_n795_), .Y(men_men_n955_));
  OAI210     u0927(.A0(men_men_n362_), .A1(men_men_n361_), .B0(men_men_n106_), .Y(men_men_n956_));
  AOI210     u0928(.A0(men_men_n956_), .A1(men_men_n525_), .B0(men_men_n955_), .Y(men_men_n957_));
  NA2        u0929(.A(men_men_n943_), .B(men_men_n900_), .Y(men_men_n958_));
  NO3        u0930(.A(l), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n959_));
  NA2        u0931(.A(men_men_n959_), .B(men_men_n611_), .Y(men_men_n960_));
  NA4        u0932(.A(men_men_n960_), .B(men_men_n958_), .C(men_men_n957_), .D(men_men_n954_), .Y(men_men_n961_));
  NO4        u0933(.A(men_men_n961_), .B(men_men_n953_), .C(men_men_n950_), .D(men_men_n933_), .Y(men_men_n962_));
  NAi31      u0934(.An(men_men_n140_), .B(men_men_n415_), .C(n), .Y(men_men_n963_));
  NA2        u0935(.A(men_men_n226_), .B(men_men_n173_), .Y(men_men_n964_));
  NO3        u0936(.A(men_men_n304_), .B(men_men_n440_), .C(men_men_n177_), .Y(men_men_n965_));
  NOi31      u0937(.An(men_men_n964_), .B(men_men_n965_), .C(men_men_n211_), .Y(men_men_n966_));
  NA2        u0938(.A(men_men_n433_), .B(men_men_n847_), .Y(men_men_n967_));
  NO2        u0939(.A(men_men_n434_), .B(men_men_n306_), .Y(men_men_n968_));
  AOI220     u0940(.A0(men_men_n968_), .A1(men_men_n967_), .B0(men_men_n474_), .B1(g), .Y(men_men_n969_));
  INV        u0941(.A(men_men_n969_), .Y(men_men_n970_));
  OAI220     u0942(.A0(men_men_n963_), .A1(men_men_n229_), .B0(men_men_n935_), .B1(men_men_n587_), .Y(men_men_n971_));
  NO2        u0943(.A(men_men_n639_), .B(men_men_n371_), .Y(men_men_n972_));
  NA2        u0944(.A(men_men_n905_), .B(men_men_n896_), .Y(men_men_n973_));
  NO3        u0945(.A(men_men_n534_), .B(men_men_n149_), .C(men_men_n210_), .Y(men_men_n974_));
  OAI210     u0946(.A0(men_men_n974_), .A1(men_men_n517_), .B0(men_men_n372_), .Y(men_men_n975_));
  OAI220     u0947(.A0(men_men_n902_), .A1(men_men_n910_), .B0(men_men_n535_), .B1(men_men_n423_), .Y(men_men_n976_));
  NA3        u0948(.A(men_men_n976_), .B(men_men_n975_), .C(men_men_n973_), .Y(men_men_n977_));
  OAI210     u0949(.A0(men_men_n905_), .A1(men_men_n897_), .B0(men_men_n964_), .Y(men_men_n978_));
  NA3        u0950(.A(c), .B(men_men_n479_), .C(men_men_n46_), .Y(men_men_n979_));
  NA2        u0951(.A(men_men_n374_), .B(men_men_n372_), .Y(men_men_n980_));
  NA4        u0952(.A(men_men_n980_), .B(men_men_n979_), .C(men_men_n978_), .D(men_men_n268_), .Y(men_men_n981_));
  OR4        u0953(.A(men_men_n981_), .B(men_men_n977_), .C(men_men_n972_), .D(men_men_n971_), .Y(men_men_n982_));
  NO4        u0954(.A(men_men_n982_), .B(men_men_n970_), .C(men_men_n966_), .D(men_men_n485_), .Y(men_men_n983_));
  NA4        u0955(.A(men_men_n983_), .B(men_men_n962_), .C(men_men_n929_), .D(men_men_n918_), .Y(men13));
  NA2        u0956(.A(men_men_n46_), .B(men_men_n82_), .Y(men_men_n985_));
  AN2        u0957(.A(c), .B(b), .Y(men_men_n986_));
  NA3        u0958(.A(men_men_n245_), .B(men_men_n986_), .C(m), .Y(men_men_n987_));
  NO3        u0959(.A(men_men_n987_), .B(men_men_n985_), .C(men_men_n567_), .Y(men_men_n988_));
  NA2        u0960(.A(men_men_n259_), .B(men_men_n986_), .Y(men_men_n989_));
  NO4        u0961(.A(men_men_n989_), .B(e), .C(men_men_n930_), .D(a), .Y(men_men_n990_));
  NAi32      u0962(.An(d), .Bn(c), .C(e), .Y(men_men_n991_));
  NA2        u0963(.A(men_men_n139_), .B(men_men_n45_), .Y(men_men_n992_));
  NO4        u0964(.A(men_men_n992_), .B(men_men_n991_), .C(men_men_n574_), .D(men_men_n303_), .Y(men_men_n993_));
  NA2        u0965(.A(men_men_n645_), .B(men_men_n220_), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n405_), .B(men_men_n210_), .Y(men_men_n995_));
  AN2        u0967(.A(d), .B(c), .Y(men_men_n996_));
  NA2        u0968(.A(men_men_n996_), .B(men_men_n113_), .Y(men_men_n997_));
  NO3        u0969(.A(men_men_n997_), .B(men_men_n995_), .C(men_men_n178_), .Y(men_men_n998_));
  NA2        u0970(.A(men_men_n490_), .B(c), .Y(men_men_n999_));
  NO4        u0971(.A(men_men_n992_), .B(men_men_n570_), .C(men_men_n999_), .D(men_men_n303_), .Y(men_men_n1000_));
  AO210      u0972(.A0(men_men_n998_), .A1(men_men_n994_), .B0(men_men_n1000_), .Y(men_men_n1001_));
  OR4        u0973(.A(men_men_n1001_), .B(men_men_n993_), .C(men_men_n990_), .D(men_men_n988_), .Y(men_men_n1002_));
  NAi32      u0974(.An(f), .Bn(e), .C(c), .Y(men_men_n1003_));
  NO2        u0975(.A(men_men_n1003_), .B(men_men_n146_), .Y(men_men_n1004_));
  NA2        u0976(.A(men_men_n1004_), .B(g), .Y(men_men_n1005_));
  OR3        u0977(.A(men_men_n220_), .B(men_men_n178_), .C(men_men_n169_), .Y(men_men_n1006_));
  NO2        u0978(.A(men_men_n1006_), .B(men_men_n1005_), .Y(men_men_n1007_));
  NO2        u0979(.A(men_men_n999_), .B(men_men_n303_), .Y(men_men_n1008_));
  NA2        u0980(.A(men_men_n614_), .B(i), .Y(men_men_n1009_));
  NOi21      u0981(.An(men_men_n1008_), .B(men_men_n1009_), .Y(men_men_n1010_));
  NOi41      u0982(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n1011_), .B(j), .Y(men_men_n1012_));
  NO2        u0984(.A(men_men_n1012_), .B(men_men_n1005_), .Y(men_men_n1013_));
  OR3        u0985(.A(e), .B(d), .C(c), .Y(men_men_n1014_));
  NA3        u0986(.A(k), .B(j), .C(i), .Y(men_men_n1015_));
  NO3        u0987(.A(men_men_n1015_), .B(men_men_n303_), .C(men_men_n86_), .Y(men_men_n1016_));
  NOi21      u0988(.An(men_men_n1016_), .B(men_men_n1014_), .Y(men_men_n1017_));
  OR4        u0989(.A(men_men_n1017_), .B(men_men_n1013_), .C(men_men_n1010_), .D(men_men_n1007_), .Y(men_men_n1018_));
  NA3        u0990(.A(men_men_n460_), .B(men_men_n330_), .C(men_men_n55_), .Y(men_men_n1019_));
  NO2        u0991(.A(men_men_n1019_), .B(men_men_n1009_), .Y(men_men_n1020_));
  NO2        u0992(.A(f), .B(c), .Y(men_men_n1021_));
  NOi21      u0993(.An(men_men_n1021_), .B(men_men_n439_), .Y(men_men_n1022_));
  NA2        u0994(.A(men_men_n1022_), .B(men_men_n58_), .Y(men_men_n1023_));
  NO3        u0995(.A(i), .B(men_men_n240_), .C(l), .Y(men_men_n1024_));
  NOi21      u0996(.An(men_men_n1024_), .B(men_men_n1023_), .Y(men_men_n1025_));
  OR2        u0997(.A(men_men_n1025_), .B(men_men_n1020_), .Y(men_men_n1026_));
  OR3        u0998(.A(men_men_n1026_), .B(men_men_n1018_), .C(men_men_n1002_), .Y(men02));
  OR3        u0999(.A(h), .B(g), .C(f), .Y(men_men_n1028_));
  OR3        u1000(.A(n), .B(m), .C(i), .Y(men_men_n1029_));
  NO4        u1001(.A(men_men_n1029_), .B(men_men_n1028_), .C(l), .D(men_men_n1014_), .Y(men_men_n1030_));
  NOi31      u1002(.An(e), .B(d), .C(c), .Y(men_men_n1031_));
  AOI210     u1003(.A0(men_men_n1016_), .A1(men_men_n1031_), .B0(men_men_n993_), .Y(men_men_n1032_));
  AN3        u1004(.A(g), .B(f), .C(c), .Y(men_men_n1033_));
  NA3        u1005(.A(men_men_n1033_), .B(men_men_n460_), .C(h), .Y(men_men_n1034_));
  OR2        u1006(.A(men_men_n1015_), .B(men_men_n303_), .Y(men_men_n1035_));
  OR2        u1007(.A(men_men_n1035_), .B(men_men_n1034_), .Y(men_men_n1036_));
  NO3        u1008(.A(men_men_n1019_), .B(men_men_n992_), .C(men_men_n570_), .Y(men_men_n1037_));
  NO2        u1009(.A(men_men_n1037_), .B(men_men_n1007_), .Y(men_men_n1038_));
  NA2        u1010(.A(i), .B(h), .Y(men_men_n1039_));
  NO2        u1011(.A(men_men_n1039_), .B(men_men_n130_), .Y(men_men_n1040_));
  NO3        u1012(.A(men_men_n141_), .B(men_men_n277_), .C(men_men_n211_), .Y(men_men_n1041_));
  AOI210     u1013(.A0(men_men_n1041_), .A1(men_men_n1040_), .B0(men_men_n1010_), .Y(men_men_n1042_));
  NA3        u1014(.A(c), .B(b), .C(a), .Y(men_men_n1043_));
  NO3        u1015(.A(men_men_n1043_), .B(men_men_n868_), .C(men_men_n210_), .Y(men_men_n1044_));
  NO3        u1016(.A(men_men_n1015_), .B(men_men_n295_), .C(men_men_n109_), .Y(men_men_n1045_));
  AOI210     u1017(.A0(men_men_n1045_), .A1(men_men_n1044_), .B0(men_men_n1020_), .Y(men_men_n1046_));
  AN4        u1018(.A(men_men_n1046_), .B(men_men_n1042_), .C(men_men_n1038_), .D(men_men_n1036_), .Y(men_men_n1047_));
  NO2        u1019(.A(men_men_n997_), .B(men_men_n995_), .Y(men_men_n1048_));
  NA2        u1020(.A(men_men_n1012_), .B(men_men_n1006_), .Y(men_men_n1049_));
  AOI210     u1021(.A0(men_men_n1049_), .A1(men_men_n1048_), .B0(men_men_n988_), .Y(men_men_n1050_));
  NAi41      u1022(.An(men_men_n1030_), .B(men_men_n1050_), .C(men_men_n1047_), .D(men_men_n1032_), .Y(men03));
  NO2        u1023(.A(men_men_n519_), .B(men_men_n581_), .Y(men_men_n1052_));
  NA4        u1024(.A(men_men_n83_), .B(men_men_n82_), .C(g), .D(men_men_n210_), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n363_), .B(men_men_n1053_), .Y(men_men_n1054_));
  NO3        u1026(.A(men_men_n1054_), .B(men_men_n1052_), .C(men_men_n956_), .Y(men_men_n1055_));
  NOi31      u1027(.An(men_men_n783_), .B(men_men_n821_), .C(men_men_n692_), .Y(men_men_n1056_));
  OAI220     u1028(.A0(men_men_n1056_), .A1(men_men_n667_), .B0(men_men_n1055_), .B1(men_men_n571_), .Y(men_men_n1057_));
  NA4        u1029(.A(i), .B(men_men_n1031_), .C(men_men_n336_), .D(men_men_n330_), .Y(men_men_n1058_));
  OAI210     u1030(.A0(men_men_n795_), .A1(men_men_n416_), .B0(men_men_n1058_), .Y(men_men_n1059_));
  NOi31      u1031(.An(m), .B(n), .C(f), .Y(men_men_n1060_));
  NA2        u1032(.A(men_men_n1060_), .B(men_men_n50_), .Y(men_men_n1061_));
  AN2        u1033(.A(e), .B(c), .Y(men_men_n1062_));
  NA2        u1034(.A(men_men_n1062_), .B(a), .Y(men_men_n1063_));
  OAI220     u1035(.A0(men_men_n1063_), .A1(men_men_n1061_), .B0(men_men_n855_), .B1(men_men_n422_), .Y(men_men_n1064_));
  NA2        u1036(.A(men_men_n500_), .B(l), .Y(men_men_n1065_));
  NOi31      u1037(.An(men_men_n835_), .B(men_men_n987_), .C(men_men_n1065_), .Y(men_men_n1066_));
  NO4        u1038(.A(men_men_n1066_), .B(men_men_n1064_), .C(men_men_n1059_), .D(men_men_n955_), .Y(men_men_n1067_));
  NO2        u1039(.A(men_men_n277_), .B(a), .Y(men_men_n1068_));
  INV        u1040(.A(men_men_n993_), .Y(men_men_n1069_));
  NO2        u1041(.A(men_men_n1039_), .B(men_men_n477_), .Y(men_men_n1070_));
  NO2        u1042(.A(men_men_n82_), .B(g), .Y(men_men_n1071_));
  NO2        u1043(.A(men_men_n1070_), .B(men_men_n1024_), .Y(men_men_n1072_));
  OR2        u1044(.A(men_men_n1072_), .B(men_men_n1023_), .Y(men_men_n1073_));
  NA3        u1045(.A(men_men_n1073_), .B(men_men_n1069_), .C(men_men_n1067_), .Y(men_men_n1074_));
  NO4        u1046(.A(men_men_n1074_), .B(men_men_n1057_), .C(men_men_n797_), .D(men_men_n554_), .Y(men_men_n1075_));
  NA2        u1047(.A(c), .B(b), .Y(men_men_n1076_));
  NO2        u1048(.A(men_men_n679_), .B(men_men_n1076_), .Y(men_men_n1077_));
  OAI210     u1049(.A0(men_men_n833_), .A1(men_men_n812_), .B0(men_men_n409_), .Y(men_men_n1078_));
  OAI210     u1050(.A0(men_men_n1078_), .A1(men_men_n834_), .B0(men_men_n1077_), .Y(men_men_n1079_));
  NAi21      u1051(.An(men_men_n417_), .B(men_men_n1077_), .Y(men_men_n1080_));
  NA3        u1052(.A(men_men_n423_), .B(men_men_n547_), .C(f), .Y(men_men_n1081_));
  OAI210     u1053(.A0(men_men_n539_), .A1(men_men_n39_), .B0(men_men_n1068_), .Y(men_men_n1082_));
  NA3        u1054(.A(men_men_n1082_), .B(men_men_n1081_), .C(men_men_n1080_), .Y(men_men_n1083_));
  NA2        u1055(.A(men_men_n255_), .B(men_men_n116_), .Y(men_men_n1084_));
  OAI210     u1056(.A0(men_men_n1084_), .A1(men_men_n281_), .B0(g), .Y(men_men_n1085_));
  NAi21      u1057(.An(f), .B(d), .Y(men_men_n1086_));
  NO2        u1058(.A(men_men_n1086_), .B(men_men_n1043_), .Y(men_men_n1087_));
  INV        u1059(.A(men_men_n1087_), .Y(men_men_n1088_));
  AOI210     u1060(.A0(men_men_n1085_), .A1(men_men_n287_), .B0(men_men_n1088_), .Y(men_men_n1089_));
  AOI210     u1061(.A0(men_men_n1089_), .A1(men_men_n110_), .B0(men_men_n1083_), .Y(men_men_n1090_));
  NA2        u1062(.A(men_men_n463_), .B(men_men_n462_), .Y(men_men_n1091_));
  NO2        u1063(.A(men_men_n183_), .B(men_men_n233_), .Y(men_men_n1092_));
  NA2        u1064(.A(men_men_n1092_), .B(m), .Y(men_men_n1093_));
  NA3        u1065(.A(men_men_n885_), .B(men_men_n1065_), .C(men_men_n466_), .Y(men_men_n1094_));
  OAI210     u1066(.A0(men_men_n1094_), .A1(men_men_n307_), .B0(men_men_n464_), .Y(men_men_n1095_));
  AOI210     u1067(.A0(men_men_n1095_), .A1(men_men_n1091_), .B0(men_men_n1093_), .Y(men_men_n1096_));
  NA2        u1068(.A(men_men_n549_), .B(men_men_n404_), .Y(men_men_n1097_));
  NA2        u1069(.A(men_men_n158_), .B(men_men_n33_), .Y(men_men_n1098_));
  AOI210     u1070(.A0(men_men_n927_), .A1(men_men_n1098_), .B0(men_men_n211_), .Y(men_men_n1099_));
  NA2        u1071(.A(men_men_n1099_), .B(men_men_n1087_), .Y(men_men_n1100_));
  AOI210     u1072(.A0(men_men_n1092_), .A1(men_men_n425_), .B0(men_men_n924_), .Y(men_men_n1101_));
  NA3        u1073(.A(men_men_n1101_), .B(men_men_n1100_), .C(men_men_n1097_), .Y(men_men_n1102_));
  NO2        u1074(.A(men_men_n1102_), .B(men_men_n1096_), .Y(men_men_n1103_));
  NA4        u1075(.A(men_men_n1103_), .B(men_men_n1090_), .C(men_men_n1079_), .D(men_men_n1075_), .Y(men00));
  AOI210     u1076(.A0(men_men_n294_), .A1(men_men_n211_), .B0(men_men_n270_), .Y(men_men_n1105_));
  NO2        u1077(.A(men_men_n1105_), .B(men_men_n562_), .Y(men_men_n1106_));
  INV        u1078(.A(men_men_n1059_), .Y(men_men_n1107_));
  NO3        u1079(.A(men_men_n1037_), .B(men_men_n924_), .C(men_men_n689_), .Y(men_men_n1108_));
  NA3        u1080(.A(men_men_n1108_), .B(men_men_n1107_), .C(men_men_n957_), .Y(men_men_n1109_));
  NA2        u1081(.A(men_men_n502_), .B(f), .Y(men_men_n1110_));
  NO2        u1082(.A(men_men_n1110_), .B(men_men_n997_), .Y(men_men_n1111_));
  NO4        u1083(.A(men_men_n1111_), .B(men_men_n1109_), .C(men_men_n1106_), .D(men_men_n1018_), .Y(men_men_n1112_));
  NA2        u1084(.A(men_men_n168_), .B(men_men_n46_), .Y(men_men_n1113_));
  NA3        u1085(.A(d), .B(men_men_n55_), .C(b), .Y(men_men_n1114_));
  NOi31      u1086(.An(n), .B(m), .C(i), .Y(men_men_n1115_));
  NA3        u1087(.A(men_men_n1115_), .B(men_men_n630_), .C(men_men_n50_), .Y(men_men_n1116_));
  OAI210     u1088(.A0(men_men_n1114_), .A1(men_men_n1113_), .B0(men_men_n1116_), .Y(men_men_n1117_));
  NO2        u1089(.A(men_men_n1117_), .B(men_men_n888_), .Y(men_men_n1118_));
  NO4        u1090(.A(men_men_n480_), .B(men_men_n348_), .C(men_men_n1076_), .D(men_men_n58_), .Y(men_men_n1119_));
  OR2        u1091(.A(men_men_n378_), .B(men_men_n133_), .Y(men_men_n1120_));
  NO2        u1092(.A(h), .B(g), .Y(men_men_n1121_));
  NA4        u1093(.A(men_men_n493_), .B(men_men_n460_), .C(men_men_n1121_), .D(men_men_n986_), .Y(men_men_n1122_));
  OAI220     u1094(.A0(men_men_n519_), .A1(men_men_n581_), .B0(men_men_n87_), .B1(men_men_n86_), .Y(men_men_n1123_));
  NA2        u1095(.A(men_men_n1123_), .B(men_men_n525_), .Y(men_men_n1124_));
  NA2        u1096(.A(men_men_n314_), .B(men_men_n242_), .Y(men_men_n1125_));
  NA4        u1097(.A(men_men_n1125_), .B(men_men_n1124_), .C(men_men_n1122_), .D(men_men_n1120_), .Y(men_men_n1126_));
  NO3        u1098(.A(men_men_n1126_), .B(men_men_n1119_), .C(men_men_n261_), .Y(men_men_n1127_));
  INV        u1099(.A(men_men_n319_), .Y(men_men_n1128_));
  AOI210     u1100(.A0(men_men_n242_), .A1(men_men_n340_), .B0(men_men_n563_), .Y(men_men_n1129_));
  NA3        u1101(.A(men_men_n1129_), .B(men_men_n1128_), .C(men_men_n153_), .Y(men_men_n1130_));
  NA3        u1102(.A(men_men_n181_), .B(men_men_n109_), .C(g), .Y(men_men_n1131_));
  NA3        u1103(.A(men_men_n460_), .B(men_men_n40_), .C(f), .Y(men_men_n1132_));
  NOi31      u1104(.An(j), .B(men_men_n1132_), .C(men_men_n1131_), .Y(men_men_n1133_));
  NAi31      u1105(.An(men_men_n184_), .B(men_men_n831_), .C(men_men_n460_), .Y(men_men_n1134_));
  NAi21      u1106(.An(men_men_n1133_), .B(men_men_n1134_), .Y(men_men_n1135_));
  NO2        u1107(.A(men_men_n269_), .B(men_men_n73_), .Y(men_men_n1136_));
  NO3        u1108(.A(men_men_n422_), .B(men_men_n808_), .C(n), .Y(men_men_n1137_));
  AOI210     u1109(.A0(men_men_n1137_), .A1(men_men_n1136_), .B0(men_men_n1030_), .Y(men_men_n1138_));
  NAi31      u1110(.An(men_men_n1000_), .B(men_men_n1138_), .C(men_men_n72_), .Y(men_men_n1139_));
  NO4        u1111(.A(men_men_n1139_), .B(men_men_n1135_), .C(men_men_n1130_), .D(men_men_n510_), .Y(men_men_n1140_));
  AN3        u1112(.A(men_men_n1140_), .B(men_men_n1127_), .C(men_men_n1118_), .Y(men_men_n1141_));
  NA2        u1113(.A(men_men_n525_), .B(men_men_n97_), .Y(men_men_n1142_));
  NA3        u1114(.A(men_men_n1060_), .B(men_men_n592_), .C(men_men_n459_), .Y(men_men_n1143_));
  NA4        u1115(.A(men_men_n1143_), .B(men_men_n550_), .C(men_men_n1142_), .D(men_men_n238_), .Y(men_men_n1144_));
  NA2        u1116(.A(men_men_n1054_), .B(men_men_n525_), .Y(men_men_n1145_));
  NA4        u1117(.A(men_men_n630_), .B(men_men_n202_), .C(men_men_n216_), .D(men_men_n162_), .Y(men_men_n1146_));
  NA3        u1118(.A(men_men_n1146_), .B(men_men_n1145_), .C(men_men_n291_), .Y(men_men_n1147_));
  OAI210     u1119(.A0(men_men_n458_), .A1(men_men_n117_), .B0(men_men_n836_), .Y(men_men_n1148_));
  AOI220     u1120(.A0(men_men_n1148_), .A1(men_men_n1094_), .B0(men_men_n549_), .B1(men_men_n404_), .Y(men_men_n1149_));
  OR4        u1121(.A(men_men_n997_), .B(men_men_n267_), .C(men_men_n218_), .D(e), .Y(men_men_n1150_));
  OAI210     u1122(.A0(men_men_n349_), .A1(men_men_n308_), .B0(men_men_n445_), .Y(men_men_n1151_));
  NA3        u1123(.A(men_men_n1151_), .B(men_men_n1150_), .C(men_men_n1149_), .Y(men_men_n1152_));
  INV        u1124(.A(men_men_n796_), .Y(men_men_n1153_));
  NO2        u1125(.A(men_men_n67_), .B(h), .Y(men_men_n1154_));
  NO3        u1126(.A(men_men_n997_), .B(men_men_n995_), .C(men_men_n706_), .Y(men_men_n1155_));
  OAI210     u1127(.A0(men_men_n1041_), .A1(men_men_n1155_), .B0(men_men_n1154_), .Y(men_men_n1156_));
  NA3        u1128(.A(men_men_n1156_), .B(men_men_n1153_), .C(men_men_n838_), .Y(men_men_n1157_));
  NO4        u1129(.A(men_men_n1157_), .B(men_men_n1152_), .C(men_men_n1147_), .D(men_men_n1144_), .Y(men_men_n1158_));
  NA2        u1130(.A(men_men_n813_), .B(men_men_n739_), .Y(men_men_n1159_));
  NA4        u1131(.A(men_men_n1159_), .B(men_men_n1158_), .C(men_men_n1141_), .D(men_men_n1112_), .Y(men01));
  AN2        u1132(.A(men_men_n975_), .B(men_men_n973_), .Y(men_men_n1161_));
  NO3        u1133(.A(men_men_n779_), .B(men_men_n773_), .C(men_men_n275_), .Y(men_men_n1162_));
  INV        u1134(.A(men_men_n388_), .Y(men_men_n1163_));
  NA3        u1135(.A(men_men_n1163_), .B(men_men_n1162_), .C(men_men_n1161_), .Y(men_men_n1164_));
  NA2        u1136(.A(men_men_n572_), .B(men_men_n85_), .Y(men_men_n1165_));
  NA2        u1137(.A(men_men_n1165_), .B(men_men_n881_), .Y(men_men_n1166_));
  NA2        u1138(.A(men_men_n45_), .B(f), .Y(men_men_n1167_));
  NA2        u1139(.A(men_men_n686_), .B(men_men_n92_), .Y(men_men_n1168_));
  NO2        u1140(.A(men_men_n1168_), .B(men_men_n1167_), .Y(men_men_n1169_));
  OAI210     u1141(.A0(men_men_n762_), .A1(men_men_n587_), .B0(men_men_n1146_), .Y(men_men_n1170_));
  AOI210     u1142(.A0(men_men_n1169_), .A1(men_men_n620_), .B0(men_men_n1170_), .Y(men_men_n1171_));
  INV        u1143(.A(men_men_n115_), .Y(men_men_n1172_));
  OA220      u1144(.A0(men_men_n1172_), .A1(men_men_n569_), .B0(men_men_n640_), .B1(men_men_n363_), .Y(men_men_n1173_));
  NAi41      u1145(.An(men_men_n161_), .B(men_men_n1173_), .C(men_men_n1171_), .D(men_men_n867_), .Y(men_men_n1174_));
  NO3        u1146(.A(men_men_n763_), .B(men_men_n653_), .C(men_men_n504_), .Y(men_men_n1175_));
  NA4        u1147(.A(men_men_n686_), .B(men_men_n92_), .C(men_men_n45_), .D(men_men_n210_), .Y(men_men_n1176_));
  OA220      u1148(.A0(men_men_n1176_), .A1(men_men_n648_), .B0(men_men_n191_), .B1(men_men_n189_), .Y(men_men_n1177_));
  NA3        u1149(.A(men_men_n1177_), .B(men_men_n1175_), .C(men_men_n136_), .Y(men_men_n1178_));
  NO4        u1150(.A(men_men_n1178_), .B(men_men_n1174_), .C(men_men_n1166_), .D(men_men_n1164_), .Y(men_men_n1179_));
  NA2        u1151(.A(men_men_n297_), .B(e), .Y(men_men_n1180_));
  NA2        u1152(.A(men_men_n528_), .B(men_men_n390_), .Y(men_men_n1181_));
  NOi21      u1153(.An(men_men_n551_), .B(men_men_n566_), .Y(men_men_n1182_));
  NA2        u1154(.A(men_men_n1182_), .B(men_men_n1181_), .Y(men_men_n1183_));
  AOI210     u1155(.A0(men_men_n200_), .A1(men_men_n84_), .B0(men_men_n210_), .Y(men_men_n1184_));
  OAI210     u1156(.A0(men_men_n786_), .A1(men_men_n423_), .B0(men_men_n1184_), .Y(men_men_n1185_));
  AN3        u1157(.A(m), .B(l), .C(k), .Y(men_men_n1186_));
  OAI210     u1158(.A0(men_men_n351_), .A1(men_men_n34_), .B0(men_men_n1186_), .Y(men_men_n1187_));
  NA2        u1159(.A(men_men_n199_), .B(men_men_n34_), .Y(men_men_n1188_));
  AO210      u1160(.A0(men_men_n1188_), .A1(men_men_n1187_), .B0(men_men_n329_), .Y(men_men_n1189_));
  NA4        u1161(.A(men_men_n1189_), .B(men_men_n1185_), .C(men_men_n1183_), .D(men_men_n1180_), .Y(men_men_n1190_));
  AOI210     u1162(.A0(men_men_n579_), .A1(men_men_n115_), .B0(men_men_n585_), .Y(men_men_n1191_));
  OAI210     u1163(.A0(men_men_n1172_), .A1(men_men_n578_), .B0(men_men_n1191_), .Y(men_men_n1192_));
  NA2        u1164(.A(men_men_n274_), .B(men_men_n191_), .Y(men_men_n1193_));
  NA2        u1165(.A(men_men_n1193_), .B(men_men_n644_), .Y(men_men_n1194_));
  NO3        u1166(.A(men_men_n795_), .B(men_men_n200_), .C(men_men_n402_), .Y(men_men_n1195_));
  NO2        u1167(.A(men_men_n1195_), .B(men_men_n924_), .Y(men_men_n1196_));
  OAI210     u1168(.A0(men_men_n1169_), .A1(men_men_n324_), .B0(men_men_n654_), .Y(men_men_n1197_));
  NA4        u1169(.A(men_men_n1197_), .B(men_men_n1196_), .C(men_men_n1194_), .D(men_men_n766_), .Y(men_men_n1198_));
  NO3        u1170(.A(men_men_n1198_), .B(men_men_n1192_), .C(men_men_n1190_), .Y(men_men_n1199_));
  NA3        u1171(.A(men_men_n588_), .B(men_men_n29_), .C(f), .Y(men_men_n1200_));
  NO2        u1172(.A(men_men_n1200_), .B(men_men_n200_), .Y(men_men_n1201_));
  INV        u1173(.A(men_men_n1201_), .Y(men_men_n1202_));
  OR3        u1174(.A(men_men_n1168_), .B(men_men_n589_), .C(men_men_n1167_), .Y(men_men_n1203_));
  NO2        u1175(.A(men_men_n1176_), .B(men_men_n938_), .Y(men_men_n1204_));
  NO2        u1176(.A(men_men_n203_), .B(men_men_n108_), .Y(men_men_n1205_));
  NO3        u1177(.A(men_men_n1205_), .B(men_men_n1204_), .C(men_men_n1117_), .Y(men_men_n1206_));
  NA4        u1178(.A(men_men_n1206_), .B(men_men_n1203_), .C(men_men_n1202_), .D(men_men_n738_), .Y(men_men_n1207_));
  INV        u1179(.A(men_men_n650_), .Y(men_men_n1208_));
  NO2        u1180(.A(men_men_n363_), .B(men_men_n71_), .Y(men_men_n1209_));
  INV        u1181(.A(men_men_n1209_), .Y(men_men_n1210_));
  NA2        u1182(.A(men_men_n1210_), .B(men_men_n380_), .Y(men_men_n1211_));
  NO3        u1183(.A(men_men_n1211_), .B(men_men_n1208_), .C(men_men_n1207_), .Y(men_men_n1212_));
  NO2        u1184(.A(men_men_n129_), .B(men_men_n45_), .Y(men_men_n1213_));
  NO2        u1185(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1214_));
  AO220      u1186(.A0(men_men_n1214_), .A1(men_men_n608_), .B0(men_men_n1213_), .B1(men_men_n684_), .Y(men_men_n1215_));
  NA2        u1187(.A(men_men_n1215_), .B(men_men_n335_), .Y(men_men_n1216_));
  INV        u1188(.A(men_men_n133_), .Y(men_men_n1217_));
  NO3        u1189(.A(men_men_n1039_), .B(men_men_n178_), .C(men_men_n82_), .Y(men_men_n1218_));
  NA2        u1190(.A(men_men_n1218_), .B(men_men_n1217_), .Y(men_men_n1219_));
  NA2        u1191(.A(men_men_n1219_), .B(men_men_n1216_), .Y(men_men_n1220_));
  NO2        u1192(.A(men_men_n600_), .B(men_men_n599_), .Y(men_men_n1221_));
  NO4        u1193(.A(men_men_n1039_), .B(men_men_n1221_), .C(men_men_n176_), .D(men_men_n82_), .Y(men_men_n1222_));
  NO3        u1194(.A(men_men_n1222_), .B(men_men_n1220_), .C(men_men_n624_), .Y(men_men_n1223_));
  NA4        u1195(.A(men_men_n1223_), .B(men_men_n1212_), .C(men_men_n1199_), .D(men_men_n1179_), .Y(men06));
  NO2        u1196(.A(men_men_n403_), .B(men_men_n548_), .Y(men_men_n1225_));
  INV        u1197(.A(men_men_n713_), .Y(men_men_n1226_));
  OAI210     u1198(.A0(men_men_n1226_), .A1(men_men_n262_), .B0(men_men_n1225_), .Y(men_men_n1227_));
  NO2        u1199(.A(men_men_n220_), .B(men_men_n99_), .Y(men_men_n1228_));
  OAI210     u1200(.A0(men_men_n1228_), .A1(men_men_n1218_), .B0(men_men_n376_), .Y(men_men_n1229_));
  NO3        u1201(.A(men_men_n583_), .B(men_men_n784_), .C(men_men_n586_), .Y(men_men_n1230_));
  OR2        u1202(.A(men_men_n1230_), .B(men_men_n855_), .Y(men_men_n1231_));
  NA3        u1203(.A(men_men_n1231_), .B(men_men_n1229_), .C(men_men_n1227_), .Y(men_men_n1232_));
  NO3        u1204(.A(men_men_n1232_), .B(men_men_n1208_), .C(men_men_n252_), .Y(men_men_n1233_));
  INV        u1205(.A(men_men_n1215_), .Y(men_men_n1234_));
  NO2        u1206(.A(men_men_n1234_), .B(men_men_n333_), .Y(men_men_n1235_));
  OAI210     u1207(.A0(men_men_n84_), .A1(men_men_n40_), .B0(men_men_n652_), .Y(men_men_n1236_));
  NA2        u1208(.A(men_men_n1236_), .B(men_men_n628_), .Y(men_men_n1237_));
  NO2        u1209(.A(men_men_n507_), .B(men_men_n173_), .Y(men_men_n1238_));
  NOi21      u1210(.An(men_men_n135_), .B(men_men_n45_), .Y(men_men_n1239_));
  NO2        u1211(.A(men_men_n593_), .B(men_men_n1061_), .Y(men_men_n1240_));
  OAI210     u1212(.A0(men_men_n454_), .A1(men_men_n243_), .B0(men_men_n875_), .Y(men_men_n1241_));
  NO4        u1213(.A(men_men_n1241_), .B(men_men_n1240_), .C(men_men_n1239_), .D(men_men_n1238_), .Y(men_men_n1242_));
  OR2        u1214(.A(men_men_n584_), .B(men_men_n582_), .Y(men_men_n1243_));
  INV        u1215(.A(men_men_n1243_), .Y(men_men_n1244_));
  NA3        u1216(.A(men_men_n1244_), .B(men_men_n1242_), .C(men_men_n1237_), .Y(men_men_n1245_));
  NO2        u1217(.A(men_men_n729_), .B(men_men_n361_), .Y(men_men_n1246_));
  NO3        u1218(.A(men_men_n654_), .B(men_men_n740_), .C(men_men_n620_), .Y(men_men_n1247_));
  NOi21      u1219(.An(men_men_n1246_), .B(men_men_n1247_), .Y(men_men_n1248_));
  NO3        u1220(.A(men_men_n1248_), .B(men_men_n1245_), .C(men_men_n1235_), .Y(men_men_n1249_));
  NO2        u1221(.A(men_men_n778_), .B(men_men_n271_), .Y(men_men_n1250_));
  OAI220     u1222(.A0(men_men_n713_), .A1(men_men_n47_), .B0(men_men_n220_), .B1(men_men_n602_), .Y(men_men_n1251_));
  OAI210     u1223(.A0(men_men_n271_), .A1(c), .B0(men_men_n627_), .Y(men_men_n1252_));
  AOI220     u1224(.A0(men_men_n1252_), .A1(men_men_n1251_), .B0(men_men_n1250_), .B1(men_men_n262_), .Y(men_men_n1253_));
  NO3        u1225(.A(men_men_n240_), .B(men_men_n99_), .C(men_men_n277_), .Y(men_men_n1254_));
  NO2        u1226(.A(men_men_n676_), .B(men_men_n243_), .Y(men_men_n1255_));
  NO2        u1227(.A(men_men_n581_), .B(j), .Y(men_men_n1256_));
  NOi21      u1228(.An(men_men_n1256_), .B(men_men_n648_), .Y(men_men_n1257_));
  NO4        u1229(.A(men_men_n1257_), .B(men_men_n1255_), .C(men_men_n1254_), .D(men_men_n1064_), .Y(men_men_n1258_));
  NA3        u1230(.A(men_men_n772_), .B(men_men_n433_), .C(men_men_n847_), .Y(men_men_n1259_));
  NAi31      u1231(.An(men_men_n729_), .B(men_men_n1259_), .C(men_men_n199_), .Y(men_men_n1260_));
  NA3        u1232(.A(men_men_n1260_), .B(men_men_n1258_), .C(men_men_n1253_), .Y(men_men_n1261_));
  NOi31      u1233(.An(men_men_n1230_), .B(men_men_n457_), .C(men_men_n389_), .Y(men_men_n1262_));
  OR3        u1234(.A(men_men_n1262_), .B(men_men_n762_), .C(men_men_n531_), .Y(men_men_n1263_));
  OR3        u1235(.A(men_men_n365_), .B(men_men_n220_), .C(men_men_n602_), .Y(men_men_n1264_));
  NA2        u1236(.A(men_men_n1256_), .B(men_men_n770_), .Y(men_men_n1265_));
  NA3        u1237(.A(men_men_n1265_), .B(men_men_n1264_), .C(men_men_n1263_), .Y(men_men_n1266_));
  NA2        u1238(.A(men_men_n1246_), .B(men_men_n739_), .Y(men_men_n1267_));
  AN2        u1239(.A(men_men_n897_), .B(men_men_n896_), .Y(men_men_n1268_));
  NO3        u1240(.A(men_men_n1268_), .B(men_men_n496_), .C(men_men_n474_), .Y(men_men_n1269_));
  NA2        u1241(.A(men_men_n1269_), .B(men_men_n1267_), .Y(men_men_n1270_));
  NAi21      u1242(.An(j), .B(i), .Y(men_men_n1271_));
  NO4        u1243(.A(men_men_n1221_), .B(men_men_n1271_), .C(men_men_n439_), .D(men_men_n231_), .Y(men_men_n1272_));
  NO4        u1244(.A(men_men_n1272_), .B(men_men_n1270_), .C(men_men_n1266_), .D(men_men_n1261_), .Y(men_men_n1273_));
  NA4        u1245(.A(men_men_n1273_), .B(men_men_n1249_), .C(men_men_n1233_), .D(men_men_n1223_), .Y(men07));
  NOi21      u1246(.An(j), .B(k), .Y(men_men_n1275_));
  NAi32      u1247(.An(m), .Bn(b), .C(n), .Y(men_men_n1276_));
  NAi21      u1248(.An(f), .B(c), .Y(men_men_n1277_));
  OR2        u1249(.A(e), .B(d), .Y(men_men_n1278_));
  NOi31      u1250(.An(n), .B(m), .C(b), .Y(men_men_n1279_));
  NOi41      u1251(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1280_));
  NA3        u1252(.A(men_men_n1280_), .B(men_men_n840_), .C(men_men_n405_), .Y(men_men_n1281_));
  INV        u1253(.A(men_men_n1281_), .Y(men_men_n1282_));
  NA2        u1254(.A(men_men_n1041_), .B(men_men_n216_), .Y(men_men_n1283_));
  NO2        u1255(.A(men_men_n1283_), .B(men_men_n60_), .Y(men_men_n1284_));
  NO2        u1256(.A(k), .B(i), .Y(men_men_n1285_));
  NO2        u1257(.A(men_men_n1015_), .B(men_men_n303_), .Y(men_men_n1286_));
  NA2        u1258(.A(men_men_n1154_), .B(men_men_n285_), .Y(men_men_n1287_));
  INV        u1259(.A(men_men_n1287_), .Y(men_men_n1288_));
  NO3        u1260(.A(men_men_n1288_), .B(men_men_n1284_), .C(men_men_n1282_), .Y(men_men_n1289_));
  NO3        u1261(.A(e), .B(d), .C(c), .Y(men_men_n1290_));
  OAI210     u1262(.A0(men_men_n130_), .A1(men_men_n211_), .B0(men_men_n590_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n1291_), .B(men_men_n1290_), .Y(men_men_n1292_));
  INV        u1264(.A(men_men_n1292_), .Y(men_men_n1293_));
  OR2        u1265(.A(h), .B(f), .Y(men_men_n1294_));
  NO3        u1266(.A(n), .B(m), .C(i), .Y(men_men_n1295_));
  OAI210     u1267(.A0(men_men_n1062_), .A1(men_men_n156_), .B0(men_men_n1295_), .Y(men_men_n1296_));
  NO2        u1268(.A(i), .B(g), .Y(men_men_n1297_));
  OR3        u1269(.A(men_men_n1297_), .B(men_men_n1276_), .C(e), .Y(men_men_n1298_));
  OAI220     u1270(.A0(men_men_n1298_), .A1(men_men_n476_), .B0(men_men_n1296_), .B1(men_men_n1294_), .Y(men_men_n1299_));
  NA3        u1271(.A(men_men_n673_), .B(men_men_n1452_), .C(men_men_n109_), .Y(men_men_n1300_));
  NA3        u1272(.A(men_men_n1279_), .B(j), .C(h), .Y(men_men_n1301_));
  AOI210     u1273(.A0(men_men_n1301_), .A1(men_men_n1300_), .B0(men_men_n45_), .Y(men_men_n1302_));
  NA2        u1274(.A(men_men_n1295_), .B(men_men_n626_), .Y(men_men_n1303_));
  NO3        u1275(.A(men_men_n439_), .B(d), .C(c), .Y(men_men_n1304_));
  NO3        u1276(.A(men_men_n1302_), .B(men_men_n1299_), .C(men_men_n1293_), .Y(men_men_n1305_));
  NO2        u1277(.A(men_men_n147_), .B(h), .Y(men_men_n1306_));
  NO2        u1278(.A(g), .B(c), .Y(men_men_n1307_));
  NO2        u1279(.A(men_men_n447_), .B(a), .Y(men_men_n1308_));
  NA3        u1280(.A(men_men_n1308_), .B(k), .C(men_men_n110_), .Y(men_men_n1309_));
  NO2        u1281(.A(i), .B(h), .Y(men_men_n1310_));
  NA2        u1282(.A(men_men_n1086_), .B(h), .Y(men_men_n1311_));
  NA2        u1283(.A(men_men_n137_), .B(men_men_n216_), .Y(men_men_n1312_));
  NO2        u1284(.A(men_men_n1312_), .B(men_men_n1311_), .Y(men_men_n1313_));
  NO2        u1285(.A(men_men_n736_), .B(men_men_n185_), .Y(men_men_n1314_));
  NOi31      u1286(.An(m), .B(n), .C(b), .Y(men_men_n1315_));
  NOi31      u1287(.An(f), .B(d), .C(c), .Y(men_men_n1316_));
  NA2        u1288(.A(men_men_n1316_), .B(men_men_n1315_), .Y(men_men_n1317_));
  INV        u1289(.A(men_men_n1317_), .Y(men_men_n1318_));
  NO3        u1290(.A(men_men_n1318_), .B(men_men_n1314_), .C(men_men_n1313_), .Y(men_men_n1319_));
  OAI210     u1291(.A0(men_men_n183_), .A1(men_men_n518_), .B0(men_men_n1011_), .Y(men_men_n1320_));
  NO3        u1292(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1321_));
  AN3        u1293(.A(men_men_n1320_), .B(men_men_n1319_), .C(men_men_n1309_), .Y(men_men_n1322_));
  NA2        u1294(.A(men_men_n1279_), .B(men_men_n373_), .Y(men_men_n1323_));
  NO2        u1295(.A(men_men_n1323_), .B(men_men_n994_), .Y(men_men_n1324_));
  NA2        u1296(.A(men_men_n1304_), .B(men_men_n212_), .Y(men_men_n1325_));
  NO2        u1297(.A(men_men_n185_), .B(b), .Y(men_men_n1326_));
  NA2        u1298(.A(men_men_n1115_), .B(men_men_n1326_), .Y(men_men_n1327_));
  NO2        u1299(.A(i), .B(men_men_n210_), .Y(men_men_n1328_));
  NA4        u1300(.A(men_men_n1092_), .B(men_men_n1328_), .C(men_men_n100_), .D(m), .Y(men_men_n1329_));
  NAi41      u1301(.An(men_men_n1324_), .B(men_men_n1329_), .C(men_men_n1327_), .D(men_men_n1325_), .Y(men_men_n1330_));
  NO4        u1302(.A(men_men_n130_), .B(g), .C(f), .D(e), .Y(men_men_n1331_));
  NA2        u1303(.A(men_men_n1285_), .B(h), .Y(men_men_n1332_));
  NA2        u1304(.A(men_men_n190_), .B(men_men_n94_), .Y(men_men_n1333_));
  NA2        u1305(.A(men_men_n30_), .B(h), .Y(men_men_n1334_));
  NO2        u1306(.A(men_men_n1334_), .B(men_men_n1029_), .Y(men_men_n1335_));
  NOi41      u1307(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1336_));
  NA2        u1308(.A(men_men_n1336_), .B(men_men_n110_), .Y(men_men_n1337_));
  INV        u1309(.A(men_men_n1337_), .Y(men_men_n1338_));
  OR3        u1310(.A(men_men_n531_), .B(men_men_n530_), .C(men_men_n109_), .Y(men_men_n1339_));
  NA2        u1311(.A(men_men_n1060_), .B(men_men_n402_), .Y(men_men_n1340_));
  OAI220     u1312(.A0(men_men_n1340_), .A1(men_men_n432_), .B0(men_men_n1339_), .B1(men_men_n295_), .Y(men_men_n1341_));
  AO210      u1313(.A0(men_men_n1341_), .A1(men_men_n113_), .B0(men_men_n1338_), .Y(men_men_n1342_));
  NO3        u1314(.A(men_men_n1342_), .B(men_men_n1335_), .C(men_men_n1330_), .Y(men_men_n1343_));
  NA4        u1315(.A(men_men_n1343_), .B(men_men_n1322_), .C(men_men_n1305_), .D(men_men_n1289_), .Y(men_men_n1344_));
  NO2        u1316(.A(men_men_n1076_), .B(men_men_n107_), .Y(men_men_n1345_));
  NA2        u1317(.A(men_men_n373_), .B(men_men_n55_), .Y(men_men_n1346_));
  AOI210     u1318(.A0(men_men_n1346_), .A1(men_men_n1003_), .B0(men_men_n1303_), .Y(men_men_n1347_));
  NA2        u1319(.A(men_men_n212_), .B(men_men_n181_), .Y(men_men_n1348_));
  AOI210     u1320(.A0(men_men_n1348_), .A1(men_men_n1131_), .B0(men_men_n1346_), .Y(men_men_n1349_));
  NO2        u1321(.A(men_men_n1034_), .B(men_men_n1029_), .Y(men_men_n1350_));
  NO3        u1322(.A(men_men_n1350_), .B(men_men_n1349_), .C(men_men_n1347_), .Y(men_men_n1351_));
  NO2        u1323(.A(men_men_n385_), .B(j), .Y(men_men_n1352_));
  NA3        u1324(.A(men_men_n1321_), .B(men_men_n1278_), .C(men_men_n1060_), .Y(men_men_n1353_));
  INV        u1325(.A(men_men_n1353_), .Y(men_men_n1354_));
  NA3        u1326(.A(g), .B(men_men_n1352_), .C(men_men_n158_), .Y(men_men_n1355_));
  INV        u1327(.A(men_men_n1355_), .Y(men_men_n1356_));
  NO3        u1328(.A(men_men_n729_), .B(men_men_n176_), .C(men_men_n405_), .Y(men_men_n1357_));
  NO3        u1329(.A(men_men_n1357_), .B(men_men_n1356_), .C(men_men_n1354_), .Y(men_men_n1358_));
  NO3        u1330(.A(men_men_n1029_), .B(men_men_n566_), .C(g), .Y(men_men_n1359_));
  NOi21      u1331(.An(men_men_n1348_), .B(men_men_n1359_), .Y(men_men_n1360_));
  AOI210     u1332(.A0(men_men_n1360_), .A1(men_men_n1333_), .B0(men_men_n1003_), .Y(men_men_n1361_));
  OR2        u1333(.A(n), .B(i), .Y(men_men_n1362_));
  OAI210     u1334(.A0(men_men_n1362_), .A1(men_men_n1021_), .B0(men_men_n49_), .Y(men_men_n1363_));
  AOI220     u1335(.A0(men_men_n1363_), .A1(men_men_n1121_), .B0(men_men_n800_), .B1(men_men_n190_), .Y(men_men_n1364_));
  INV        u1336(.A(men_men_n1364_), .Y(men_men_n1365_));
  NA2        u1337(.A(men_men_n1326_), .B(men_men_n41_), .Y(men_men_n1366_));
  NO2        u1338(.A(men_men_n130_), .B(l), .Y(men_men_n1367_));
  NO2        u1339(.A(men_men_n220_), .B(k), .Y(men_men_n1368_));
  OAI210     u1340(.A0(men_men_n1368_), .A1(men_men_n1310_), .B0(men_men_n1367_), .Y(men_men_n1369_));
  OAI220     u1341(.A0(men_men_n1369_), .A1(men_men_n31_), .B0(men_men_n1366_), .B1(men_men_n178_), .Y(men_men_n1370_));
  NO3        u1342(.A(men_men_n1370_), .B(men_men_n1365_), .C(men_men_n1361_), .Y(men_men_n1371_));
  INV        u1343(.A(men_men_n49_), .Y(men_men_n1372_));
  NO3        u1344(.A(men_men_n1043_), .B(men_men_n1278_), .C(men_men_n49_), .Y(men_men_n1373_));
  NA2        u1345(.A(men_men_n1044_), .B(men_men_n1372_), .Y(men_men_n1374_));
  NO2        u1346(.A(men_men_n1374_), .B(j), .Y(men_men_n1375_));
  NA3        u1347(.A(men_men_n1345_), .B(men_men_n460_), .C(f), .Y(men_men_n1376_));
  NA2        u1348(.A(men_men_n181_), .B(men_men_n109_), .Y(men_men_n1377_));
  NO2        u1349(.A(men_men_n1275_), .B(men_men_n42_), .Y(men_men_n1378_));
  AOI210     u1350(.A0(men_men_n110_), .A1(men_men_n40_), .B0(men_men_n1378_), .Y(men_men_n1379_));
  NO2        u1351(.A(men_men_n1379_), .B(men_men_n1376_), .Y(men_men_n1380_));
  AOI210     u1352(.A0(men_men_n518_), .A1(h), .B0(men_men_n68_), .Y(men_men_n1381_));
  NA2        u1353(.A(men_men_n1381_), .B(men_men_n1308_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n1271_), .B(men_men_n176_), .Y(men_men_n1383_));
  NOi21      u1355(.An(d), .B(f), .Y(men_men_n1384_));
  NO3        u1356(.A(men_men_n1316_), .B(men_men_n1384_), .C(men_men_n40_), .Y(men_men_n1385_));
  NA2        u1357(.A(men_men_n1385_), .B(men_men_n1383_), .Y(men_men_n1386_));
  NA2        u1358(.A(men_men_n1308_), .B(men_men_n1378_), .Y(men_men_n1387_));
  NO2        u1359(.A(men_men_n295_), .B(c), .Y(men_men_n1388_));
  NA2        u1360(.A(men_men_n1388_), .B(men_men_n532_), .Y(men_men_n1389_));
  NA4        u1361(.A(men_men_n1389_), .B(men_men_n1387_), .C(men_men_n1386_), .D(men_men_n1382_), .Y(men_men_n1390_));
  NO3        u1362(.A(men_men_n1390_), .B(men_men_n1380_), .C(men_men_n1375_), .Y(men_men_n1391_));
  NA4        u1363(.A(men_men_n1391_), .B(men_men_n1371_), .C(men_men_n1358_), .D(men_men_n1351_), .Y(men_men_n1392_));
  NO3        u1364(.A(men_men_n1033_), .B(men_men_n1021_), .C(men_men_n40_), .Y(men_men_n1393_));
  NO2        u1365(.A(men_men_n460_), .B(men_men_n295_), .Y(men_men_n1394_));
  OAI210     u1366(.A0(men_men_n1394_), .A1(men_men_n1393_), .B0(men_men_n1286_), .Y(men_men_n1395_));
  OAI210     u1367(.A0(men_men_n1331_), .A1(men_men_n1279_), .B0(men_men_n852_), .Y(men_men_n1396_));
  OAI220     u1368(.A0(men_men_n991_), .A1(men_men_n130_), .B0(men_men_n645_), .B1(men_men_n176_), .Y(men_men_n1397_));
  NA2        u1369(.A(men_men_n1397_), .B(men_men_n607_), .Y(men_men_n1398_));
  NA3        u1370(.A(men_men_n1398_), .B(men_men_n1396_), .C(men_men_n1395_), .Y(men_men_n1399_));
  NA2        u1371(.A(men_men_n1307_), .B(men_men_n1384_), .Y(men_men_n1400_));
  NO2        u1372(.A(men_men_n1400_), .B(m), .Y(men_men_n1401_));
  NA3        u1373(.A(men_men_n1041_), .B(men_men_n105_), .C(men_men_n216_), .Y(men_men_n1402_));
  NA2        u1374(.A(men_men_n107_), .B(men_men_n1315_), .Y(men_men_n1403_));
  NA2        u1375(.A(men_men_n1403_), .B(men_men_n1402_), .Y(men_men_n1404_));
  NO3        u1376(.A(men_men_n1404_), .B(men_men_n1401_), .C(men_men_n1399_), .Y(men_men_n1405_));
  NO2        u1377(.A(men_men_n1277_), .B(e), .Y(men_men_n1406_));
  INV        u1378(.A(men_men_n1406_), .Y(men_men_n1407_));
  NA2        u1379(.A(men_men_n1071_), .B(men_men_n616_), .Y(men_men_n1408_));
  OR3        u1380(.A(men_men_n1368_), .B(men_men_n1154_), .C(men_men_n130_), .Y(men_men_n1409_));
  OAI220     u1381(.A0(men_men_n1409_), .A1(men_men_n1407_), .B0(men_men_n1408_), .B1(men_men_n441_), .Y(men_men_n1410_));
  NO3        u1382(.A(men_men_n1339_), .B(men_men_n347_), .C(a), .Y(men_men_n1411_));
  NO2        u1383(.A(men_men_n1411_), .B(men_men_n1410_), .Y(men_men_n1412_));
  AOI210     u1384(.A0(men_men_n868_), .A1(men_men_n412_), .B0(men_men_n101_), .Y(men_men_n1413_));
  OR2        u1385(.A(men_men_n1413_), .B(men_men_n530_), .Y(men_men_n1414_));
  NO2        u1386(.A(men_men_n1414_), .B(men_men_n176_), .Y(men_men_n1415_));
  NO2        u1387(.A(men_men_n49_), .B(l), .Y(men_men_n1416_));
  INV        u1388(.A(men_men_n476_), .Y(men_men_n1417_));
  OAI210     u1389(.A0(men_men_n1417_), .A1(men_men_n1044_), .B0(men_men_n1416_), .Y(men_men_n1418_));
  NO2        u1390(.A(men_men_n248_), .B(g), .Y(men_men_n1419_));
  NO2        u1391(.A(m), .B(i), .Y(men_men_n1420_));
  BUFFER     u1392(.A(men_men_n1420_), .Y(men_men_n1421_));
  AOI220     u1393(.A0(men_men_n1421_), .A1(men_men_n1306_), .B0(men_men_n1022_), .B1(men_men_n1419_), .Y(men_men_n1422_));
  NA2        u1394(.A(men_men_n1422_), .B(men_men_n1418_), .Y(men_men_n1423_));
  NO3        u1395(.A(men_men_n1423_), .B(men_men_n1415_), .C(men_men_n1373_), .Y(men_men_n1424_));
  NA3        u1396(.A(men_men_n1424_), .B(men_men_n1412_), .C(men_men_n1405_), .Y(men_men_n1425_));
  NA3        u1397(.A(men_men_n926_), .B(men_men_n137_), .C(men_men_n46_), .Y(men_men_n1426_));
  NO2        u1398(.A(e), .B(c), .Y(men_men_n1427_));
  NO3        u1399(.A(men_men_n184_), .B(men_men_n446_), .C(men_men_n45_), .Y(men_men_n1428_));
  AOI210     u1400(.A0(men_men_n1383_), .A1(men_men_n1427_), .B0(men_men_n1428_), .Y(men_men_n1429_));
  AOI210     u1401(.A0(men_men_n156_), .A1(men_men_n55_), .B0(men_men_n1406_), .Y(men_men_n1430_));
  NO2        u1402(.A(men_men_n1430_), .B(men_men_n1377_), .Y(men_men_n1431_));
  NO2        u1403(.A(men_men_n1426_), .B(men_men_n107_), .Y(men_men_n1432_));
  NO2        u1404(.A(men_men_n1432_), .B(men_men_n1431_), .Y(men_men_n1433_));
  NO2        u1405(.A(men_men_n1376_), .B(men_men_n68_), .Y(men_men_n1434_));
  NO2        u1406(.A(men_men_n1285_), .B(men_men_n115_), .Y(men_men_n1435_));
  NO2        u1407(.A(men_men_n1435_), .B(men_men_n1323_), .Y(men_men_n1436_));
  NO2        u1408(.A(men_men_n1436_), .B(men_men_n1434_), .Y(men_men_n1437_));
  NA3        u1409(.A(men_men_n1437_), .B(men_men_n1433_), .C(men_men_n1429_), .Y(men_men_n1438_));
  OR4        u1410(.A(men_men_n1438_), .B(men_men_n1425_), .C(men_men_n1392_), .D(men_men_n1344_), .Y(men04));
  NOi31      u1411(.An(men_men_n1331_), .B(men_men_n1332_), .C(men_men_n997_), .Y(men_men_n1440_));
  NO4        u1412(.A(men_men_n267_), .B(men_men_n987_), .C(men_men_n477_), .D(j), .Y(men_men_n1441_));
  OR3        u1413(.A(men_men_n1441_), .B(men_men_n1440_), .C(men_men_n1013_), .Y(men_men_n1442_));
  NO2        u1414(.A(men_men_n86_), .B(k), .Y(men_men_n1443_));
  AOI210     u1415(.A0(men_men_n1443_), .A1(men_men_n1008_), .B0(men_men_n1133_), .Y(men_men_n1444_));
  NA2        u1416(.A(men_men_n1444_), .B(men_men_n1156_), .Y(men_men_n1445_));
  NO3        u1417(.A(men_men_n1445_), .B(men_men_n1442_), .C(men_men_n1002_), .Y(men_men_n1446_));
  NA4        u1418(.A(men_men_n1446_), .B(men_men_n1073_), .C(men_men_n1058_), .D(men_men_n1047_), .Y(men05));
  INV        u1419(.A(men_men_n867_), .Y(men_men_n1450_));
  INV        u1420(.A(f), .Y(men_men_n1451_));
  INV        u1421(.A(n), .Y(men_men_n1452_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule