//Benchmark atmr_max1024_476_0.0313

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  INV        o005(.A(ori_ori_n19_), .Y(ori_ori_n22_));
  NA2        o006(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n23_));
  INV        o007(.A(x5), .Y(ori_ori_n24_));
  NA2        o008(.A(x7), .B(x6), .Y(ori_ori_n25_));
  NA2        o009(.A(x8), .B(x3), .Y(ori_ori_n26_));
  NA2        o010(.A(x4), .B(x2), .Y(ori_ori_n27_));
  NO4        o011(.A(ori_ori_n27_), .B(ori_ori_n26_), .C(ori_ori_n25_), .D(ori_ori_n24_), .Y(ori_ori_n28_));
  NO2        o012(.A(ori_ori_n28_), .B(ori_ori_n23_), .Y(ori_ori_n29_));
  NO2        o013(.A(x4), .B(x3), .Y(ori_ori_n30_));
  INV        o014(.A(ori_ori_n30_), .Y(ori_ori_n31_));
  NOi21      o015(.An(ori_ori_n22_), .B(ori_ori_n29_), .Y(ori00));
  NO2        o016(.A(x1), .B(x0), .Y(ori_ori_n33_));
  INV        o017(.A(x6), .Y(ori_ori_n34_));
  NO2        o018(.A(ori_ori_n34_), .B(ori_ori_n24_), .Y(ori_ori_n35_));
  AN2        o019(.A(x8), .B(x7), .Y(ori_ori_n36_));
  NA3        o020(.A(ori_ori_n36_), .B(ori_ori_n35_), .C(ori_ori_n33_), .Y(ori_ori_n37_));
  NA2        o021(.A(x4), .B(x3), .Y(ori_ori_n38_));
  AOI210     o022(.A0(ori_ori_n37_), .A1(ori_ori_n22_), .B0(ori_ori_n38_), .Y(ori_ori_n39_));
  NO2        o023(.A(x2), .B(x0), .Y(ori_ori_n40_));
  INV        o024(.A(x3), .Y(ori_ori_n41_));
  NO2        o025(.A(ori_ori_n41_), .B(ori_ori_n18_), .Y(ori_ori_n42_));
  INV        o026(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n35_), .B(x4), .Y(ori_ori_n44_));
  OAI210     o028(.A0(ori_ori_n44_), .A1(ori_ori_n43_), .B0(ori_ori_n40_), .Y(ori_ori_n45_));
  INV        o029(.A(x4), .Y(ori_ori_n46_));
  NO2        o030(.A(ori_ori_n46_), .B(ori_ori_n17_), .Y(ori_ori_n47_));
  NA2        o031(.A(ori_ori_n47_), .B(x2), .Y(ori_ori_n48_));
  OAI210     o032(.A0(ori_ori_n48_), .A1(ori_ori_n20_), .B0(ori_ori_n45_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n50_));
  NA2        o034(.A(ori_ori_n50_), .B(ori_ori_n33_), .Y(ori_ori_n51_));
  INV        o035(.A(x2), .Y(ori_ori_n52_));
  NO2        o036(.A(ori_ori_n52_), .B(ori_ori_n17_), .Y(ori_ori_n53_));
  NA2        o037(.A(ori_ori_n41_), .B(ori_ori_n18_), .Y(ori_ori_n54_));
  NA2        o038(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  OAI210     o039(.A0(ori_ori_n51_), .A1(ori_ori_n31_), .B0(ori_ori_n55_), .Y(ori_ori_n56_));
  NO3        o040(.A(ori_ori_n56_), .B(ori_ori_n49_), .C(ori_ori_n39_), .Y(ori01));
  NA2        o041(.A(x8), .B(x7), .Y(ori_ori_n58_));
  NA2        o042(.A(ori_ori_n41_), .B(x1), .Y(ori_ori_n59_));
  INV        o043(.A(x9), .Y(ori_ori_n60_));
  NO2        o044(.A(ori_ori_n60_), .B(ori_ori_n34_), .Y(ori_ori_n61_));
  INV        o045(.A(ori_ori_n61_), .Y(ori_ori_n62_));
  NO3        o046(.A(ori_ori_n62_), .B(ori_ori_n59_), .C(ori_ori_n58_), .Y(ori_ori_n63_));
  NO2        o047(.A(x7), .B(x6), .Y(ori_ori_n64_));
  NO2        o048(.A(ori_ori_n59_), .B(x5), .Y(ori_ori_n65_));
  NO2        o049(.A(x8), .B(x2), .Y(ori_ori_n66_));
  INV        o050(.A(ori_ori_n66_), .Y(ori_ori_n67_));
  AN2        o051(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n68_));
  OAI210     o052(.A0(ori_ori_n42_), .A1(ori_ori_n24_), .B0(ori_ori_n52_), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n54_), .A1(ori_ori_n20_), .B0(ori_ori_n69_), .Y(ori_ori_n70_));
  NO2        o054(.A(ori_ori_n70_), .B(ori_ori_n68_), .Y(ori_ori_n71_));
  OAI210     o055(.A0(ori_ori_n71_), .A1(ori_ori_n63_), .B0(x4), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n46_), .B(x2), .Y(ori_ori_n73_));
  OAI210     o057(.A0(ori_ori_n73_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n74_));
  NA2        o058(.A(x5), .B(x3), .Y(ori_ori_n75_));
  NO2        o059(.A(x8), .B(x6), .Y(ori_ori_n76_));
  NO4        o060(.A(ori_ori_n76_), .B(ori_ori_n75_), .C(ori_ori_n64_), .D(ori_ori_n52_), .Y(ori_ori_n77_));
  NAi21      o061(.An(x4), .B(x3), .Y(ori_ori_n78_));
  INV        o062(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NO2        o063(.A(x4), .B(x2), .Y(ori_ori_n80_));
  NO2        o064(.A(ori_ori_n78_), .B(ori_ori_n18_), .Y(ori_ori_n81_));
  NO3        o065(.A(ori_ori_n81_), .B(ori_ori_n77_), .C(ori_ori_n74_), .Y(ori_ori_n82_));
  NA2        o066(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n83_));
  NO2        o067(.A(ori_ori_n83_), .B(ori_ori_n24_), .Y(ori_ori_n84_));
  INV        o068(.A(x8), .Y(ori_ori_n85_));
  NA2        o069(.A(x2), .B(x1), .Y(ori_ori_n86_));
  NO2        o070(.A(ori_ori_n86_), .B(ori_ori_n85_), .Y(ori_ori_n87_));
  NO2        o071(.A(ori_ori_n87_), .B(ori_ori_n84_), .Y(ori_ori_n88_));
  NO2        o072(.A(ori_ori_n88_), .B(ori_ori_n25_), .Y(ori_ori_n89_));
  AOI210     o073(.A0(ori_ori_n54_), .A1(ori_ori_n24_), .B0(ori_ori_n52_), .Y(ori_ori_n90_));
  OAI210     o074(.A0(ori_ori_n43_), .A1(ori_ori_n35_), .B0(ori_ori_n46_), .Y(ori_ori_n91_));
  NO3        o075(.A(ori_ori_n91_), .B(ori_ori_n90_), .C(ori_ori_n89_), .Y(ori_ori_n92_));
  NA2        o076(.A(x4), .B(ori_ori_n41_), .Y(ori_ori_n93_));
  NO2        o077(.A(ori_ori_n46_), .B(ori_ori_n52_), .Y(ori_ori_n94_));
  OAI210     o078(.A0(ori_ori_n94_), .A1(ori_ori_n41_), .B0(ori_ori_n18_), .Y(ori_ori_n95_));
  AOI210     o079(.A0(ori_ori_n93_), .A1(ori_ori_n50_), .B0(ori_ori_n95_), .Y(ori_ori_n96_));
  NO2        o080(.A(x3), .B(x2), .Y(ori_ori_n97_));
  NA3        o081(.A(ori_ori_n97_), .B(ori_ori_n25_), .C(ori_ori_n24_), .Y(ori_ori_n98_));
  AOI210     o082(.A0(x8), .A1(x6), .B0(ori_ori_n98_), .Y(ori_ori_n99_));
  NA2        o083(.A(ori_ori_n52_), .B(x1), .Y(ori_ori_n100_));
  OAI210     o084(.A0(ori_ori_n100_), .A1(ori_ori_n38_), .B0(ori_ori_n17_), .Y(ori_ori_n101_));
  NO4        o085(.A(ori_ori_n101_), .B(ori_ori_n99_), .C(ori_ori_n96_), .D(ori_ori_n92_), .Y(ori_ori_n102_));
  AO210      o086(.A0(ori_ori_n82_), .A1(ori_ori_n72_), .B0(ori_ori_n102_), .Y(ori02));
  NO2        o087(.A(x3), .B(ori_ori_n52_), .Y(ori_ori_n104_));
  NO2        o088(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n105_));
  NA2        o089(.A(ori_ori_n52_), .B(ori_ori_n17_), .Y(ori_ori_n106_));
  NA2        o090(.A(ori_ori_n41_), .B(x0), .Y(ori_ori_n107_));
  NA2        o091(.A(ori_ori_n104_), .B(x4), .Y(ori_ori_n108_));
  NO3        o092(.A(ori_ori_n108_), .B(x7), .C(x5), .Y(ori_ori_n109_));
  NA2        o093(.A(x9), .B(x2), .Y(ori_ori_n110_));
  OR2        o094(.A(x8), .B(x0), .Y(ori_ori_n111_));
  INV        o095(.A(ori_ori_n111_), .Y(ori_ori_n112_));
  NAi21      o096(.An(x2), .B(x8), .Y(ori_ori_n113_));
  NO2        o097(.A(x4), .B(x1), .Y(ori_ori_n114_));
  NA3        o098(.A(ori_ori_n114_), .B(x2), .C(ori_ori_n58_), .Y(ori_ori_n115_));
  NOi21      o099(.An(x0), .B(x1), .Y(ori_ori_n116_));
  NO3        o100(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n117_));
  NOi21      o101(.An(x0), .B(x4), .Y(ori_ori_n118_));
  NAi21      o102(.An(x8), .B(x7), .Y(ori_ori_n119_));
  NO2        o103(.A(ori_ori_n119_), .B(ori_ori_n60_), .Y(ori_ori_n120_));
  AOI220     o104(.A0(ori_ori_n120_), .A1(ori_ori_n118_), .B0(ori_ori_n117_), .B1(ori_ori_n116_), .Y(ori_ori_n121_));
  AOI210     o105(.A0(ori_ori_n121_), .A1(ori_ori_n115_), .B0(ori_ori_n75_), .Y(ori_ori_n122_));
  NO2        o106(.A(x5), .B(ori_ori_n46_), .Y(ori_ori_n123_));
  NA2        o107(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n124_));
  AOI210     o108(.A0(ori_ori_n124_), .A1(ori_ori_n100_), .B0(ori_ori_n107_), .Y(ori_ori_n125_));
  OAI210     o109(.A0(ori_ori_n125_), .A1(ori_ori_n33_), .B0(ori_ori_n123_), .Y(ori_ori_n126_));
  NAi21      o110(.An(x0), .B(x4), .Y(ori_ori_n127_));
  NO2        o111(.A(ori_ori_n127_), .B(x1), .Y(ori_ori_n128_));
  NO2        o112(.A(x7), .B(x0), .Y(ori_ori_n129_));
  NO2        o113(.A(ori_ori_n80_), .B(ori_ori_n94_), .Y(ori_ori_n130_));
  NO2        o114(.A(ori_ori_n130_), .B(x3), .Y(ori_ori_n131_));
  OAI210     o115(.A0(ori_ori_n129_), .A1(ori_ori_n128_), .B0(ori_ori_n131_), .Y(ori_ori_n132_));
  NA2        o116(.A(x5), .B(x0), .Y(ori_ori_n133_));
  NO2        o117(.A(ori_ori_n46_), .B(x2), .Y(ori_ori_n134_));
  NA3        o118(.A(ori_ori_n132_), .B(ori_ori_n126_), .C(ori_ori_n34_), .Y(ori_ori_n135_));
  NO3        o119(.A(ori_ori_n135_), .B(ori_ori_n122_), .C(ori_ori_n109_), .Y(ori_ori_n136_));
  NO3        o120(.A(ori_ori_n75_), .B(ori_ori_n73_), .C(ori_ori_n23_), .Y(ori_ori_n137_));
  NO2        o121(.A(ori_ori_n27_), .B(ori_ori_n24_), .Y(ori_ori_n138_));
  AOI220     o122(.A0(ori_ori_n116_), .A1(ori_ori_n138_), .B0(ori_ori_n65_), .B1(ori_ori_n17_), .Y(ori_ori_n139_));
  NO3        o123(.A(ori_ori_n139_), .B(ori_ori_n58_), .C(ori_ori_n60_), .Y(ori_ori_n140_));
  NA2        o124(.A(x7), .B(x3), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n93_), .B(x5), .Y(ori_ori_n142_));
  NO2        o126(.A(x9), .B(x7), .Y(ori_ori_n143_));
  NOi21      o127(.An(x8), .B(x0), .Y(ori_ori_n144_));
  OA210      o128(.A0(ori_ori_n143_), .A1(x1), .B0(ori_ori_n144_), .Y(ori_ori_n145_));
  NO2        o129(.A(ori_ori_n41_), .B(x2), .Y(ori_ori_n146_));
  INV        o130(.A(x7), .Y(ori_ori_n147_));
  NA2        o131(.A(ori_ori_n147_), .B(ori_ori_n18_), .Y(ori_ori_n148_));
  AOI220     o132(.A0(ori_ori_n148_), .A1(ori_ori_n146_), .B0(ori_ori_n104_), .B1(ori_ori_n36_), .Y(ori_ori_n149_));
  NO2        o133(.A(ori_ori_n24_), .B(x4), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n150_), .B(ori_ori_n118_), .Y(ori_ori_n151_));
  NO2        o135(.A(ori_ori_n151_), .B(ori_ori_n149_), .Y(ori_ori_n152_));
  AOI210     o136(.A0(ori_ori_n145_), .A1(ori_ori_n142_), .B0(ori_ori_n152_), .Y(ori_ori_n153_));
  OAI210     o137(.A0(ori_ori_n141_), .A1(ori_ori_n48_), .B0(ori_ori_n153_), .Y(ori_ori_n154_));
  NA2        o138(.A(x5), .B(x1), .Y(ori_ori_n155_));
  INV        o139(.A(ori_ori_n155_), .Y(ori_ori_n156_));
  AOI210     o140(.A0(ori_ori_n156_), .A1(ori_ori_n118_), .B0(ori_ori_n34_), .Y(ori_ori_n157_));
  NO2        o141(.A(ori_ori_n60_), .B(ori_ori_n85_), .Y(ori_ori_n158_));
  NAi21      o142(.An(x2), .B(x7), .Y(ori_ori_n159_));
  NO3        o143(.A(ori_ori_n159_), .B(ori_ori_n158_), .C(ori_ori_n46_), .Y(ori_ori_n160_));
  NA2        o144(.A(ori_ori_n160_), .B(ori_ori_n65_), .Y(ori_ori_n161_));
  NAi31      o145(.An(ori_ori_n75_), .B(ori_ori_n36_), .C(ori_ori_n33_), .Y(ori_ori_n162_));
  NA3        o146(.A(ori_ori_n162_), .B(ori_ori_n161_), .C(ori_ori_n157_), .Y(ori_ori_n163_));
  NO4        o147(.A(ori_ori_n163_), .B(ori_ori_n154_), .C(ori_ori_n140_), .D(ori_ori_n137_), .Y(ori_ori_n164_));
  NO2        o148(.A(ori_ori_n164_), .B(ori_ori_n136_), .Y(ori_ori_n165_));
  NO2        o149(.A(ori_ori_n133_), .B(ori_ori_n130_), .Y(ori_ori_n166_));
  NA2        o150(.A(ori_ori_n24_), .B(ori_ori_n18_), .Y(ori_ori_n167_));
  NA2        o151(.A(ori_ori_n24_), .B(ori_ori_n17_), .Y(ori_ori_n168_));
  NA3        o152(.A(ori_ori_n168_), .B(ori_ori_n167_), .C(ori_ori_n23_), .Y(ori_ori_n169_));
  AN2        o153(.A(ori_ori_n169_), .B(ori_ori_n134_), .Y(ori_ori_n170_));
  NA2        o154(.A(x8), .B(x0), .Y(ori_ori_n171_));
  NO2        o155(.A(ori_ori_n147_), .B(ori_ori_n24_), .Y(ori_ori_n172_));
  NO2        o156(.A(ori_ori_n116_), .B(x4), .Y(ori_ori_n173_));
  NA2        o157(.A(ori_ori_n173_), .B(ori_ori_n172_), .Y(ori_ori_n174_));
  AOI210     o158(.A0(ori_ori_n171_), .A1(ori_ori_n124_), .B0(ori_ori_n174_), .Y(ori_ori_n175_));
  NA2        o159(.A(x2), .B(x0), .Y(ori_ori_n176_));
  NA2        o160(.A(x4), .B(x1), .Y(ori_ori_n177_));
  NAi21      o161(.An(ori_ori_n114_), .B(ori_ori_n177_), .Y(ori_ori_n178_));
  NOi31      o162(.An(ori_ori_n178_), .B(ori_ori_n150_), .C(ori_ori_n176_), .Y(ori_ori_n179_));
  NO4        o163(.A(ori_ori_n179_), .B(ori_ori_n175_), .C(ori_ori_n170_), .D(ori_ori_n166_), .Y(ori_ori_n180_));
  NO2        o164(.A(ori_ori_n180_), .B(ori_ori_n41_), .Y(ori_ori_n181_));
  NO2        o165(.A(ori_ori_n169_), .B(ori_ori_n73_), .Y(ori_ori_n182_));
  INV        o166(.A(ori_ori_n123_), .Y(ori_ori_n183_));
  NO2        o167(.A(ori_ori_n100_), .B(ori_ori_n17_), .Y(ori_ori_n184_));
  AOI210     o168(.A0(ori_ori_n33_), .A1(ori_ori_n85_), .B0(ori_ori_n184_), .Y(ori_ori_n185_));
  NO3        o169(.A(ori_ori_n185_), .B(ori_ori_n183_), .C(x7), .Y(ori_ori_n186_));
  NA3        o170(.A(ori_ori_n178_), .B(ori_ori_n183_), .C(ori_ori_n40_), .Y(ori_ori_n187_));
  OAI210     o171(.A0(ori_ori_n168_), .A1(ori_ori_n130_), .B0(ori_ori_n187_), .Y(ori_ori_n188_));
  NO3        o172(.A(ori_ori_n188_), .B(ori_ori_n186_), .C(ori_ori_n182_), .Y(ori_ori_n189_));
  NO2        o173(.A(ori_ori_n189_), .B(x3), .Y(ori_ori_n190_));
  NO3        o174(.A(ori_ori_n190_), .B(ori_ori_n181_), .C(ori_ori_n165_), .Y(ori03));
  NO2        o175(.A(ori_ori_n46_), .B(x3), .Y(ori_ori_n192_));
  NO2        o176(.A(x6), .B(ori_ori_n24_), .Y(ori_ori_n193_));
  INV        o177(.A(ori_ori_n193_), .Y(ori_ori_n194_));
  NO2        o178(.A(ori_ori_n52_), .B(x1), .Y(ori_ori_n195_));
  OAI210     o179(.A0(ori_ori_n195_), .A1(ori_ori_n24_), .B0(ori_ori_n61_), .Y(ori_ori_n196_));
  OAI220     o180(.A0(ori_ori_n196_), .A1(ori_ori_n17_), .B0(ori_ori_n194_), .B1(ori_ori_n100_), .Y(ori_ori_n197_));
  NA2        o181(.A(ori_ori_n197_), .B(ori_ori_n192_), .Y(ori_ori_n198_));
  NA2        o182(.A(x6), .B(ori_ori_n24_), .Y(ori_ori_n199_));
  NO2        o183(.A(ori_ori_n199_), .B(x4), .Y(ori_ori_n200_));
  NO2        o184(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n201_));
  NA2        o185(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n202_));
  NO2        o186(.A(ori_ori_n202_), .B(ori_ori_n199_), .Y(ori_ori_n203_));
  NA2        o187(.A(x9), .B(ori_ori_n52_), .Y(ori_ori_n204_));
  NA2        o188(.A(ori_ori_n204_), .B(x4), .Y(ori_ori_n205_));
  NA2        o189(.A(ori_ori_n199_), .B(ori_ori_n78_), .Y(ori_ori_n206_));
  AOI210     o190(.A0(ori_ori_n24_), .A1(x3), .B0(ori_ori_n176_), .Y(ori_ori_n207_));
  AOI220     o191(.A0(ori_ori_n207_), .A1(ori_ori_n206_), .B0(ori_ori_n205_), .B1(ori_ori_n203_), .Y(ori_ori_n208_));
  NO3        o192(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n209_));
  NO2        o193(.A(x5), .B(x1), .Y(ori_ori_n210_));
  NO2        o194(.A(ori_ori_n202_), .B(ori_ori_n167_), .Y(ori_ori_n211_));
  NO3        o195(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n212_));
  NO2        o196(.A(ori_ori_n212_), .B(ori_ori_n211_), .Y(ori_ori_n213_));
  INV        o197(.A(ori_ori_n213_), .Y(ori_ori_n214_));
  AOI220     o198(.A0(ori_ori_n214_), .A1(ori_ori_n46_), .B0(ori_ori_n209_), .B1(ori_ori_n123_), .Y(ori_ori_n215_));
  NA3        o199(.A(ori_ori_n215_), .B(ori_ori_n208_), .C(ori_ori_n198_), .Y(ori_ori_n216_));
  NO2        o200(.A(ori_ori_n46_), .B(ori_ori_n41_), .Y(ori_ori_n217_));
  NA2        o201(.A(ori_ori_n217_), .B(ori_ori_n19_), .Y(ori_ori_n218_));
  NO2        o202(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n219_));
  NO2        o203(.A(ori_ori_n219_), .B(x6), .Y(ori_ori_n220_));
  NOi21      o204(.An(ori_ori_n80_), .B(ori_ori_n220_), .Y(ori_ori_n221_));
  NA2        o205(.A(ori_ori_n60_), .B(ori_ori_n85_), .Y(ori_ori_n222_));
  NA3        o206(.A(ori_ori_n222_), .B(ori_ori_n219_), .C(x6), .Y(ori_ori_n223_));
  AOI210     o207(.A0(ori_ori_n223_), .A1(ori_ori_n221_), .B0(ori_ori_n147_), .Y(ori_ori_n224_));
  OR2        o208(.A(ori_ori_n224_), .B(ori_ori_n172_), .Y(ori_ori_n225_));
  NA2        o209(.A(ori_ori_n41_), .B(ori_ori_n52_), .Y(ori_ori_n226_));
  OAI210     o210(.A0(ori_ori_n226_), .A1(ori_ori_n24_), .B0(ori_ori_n168_), .Y(ori_ori_n227_));
  NO3        o211(.A(ori_ori_n177_), .B(ori_ori_n60_), .C(x6), .Y(ori_ori_n228_));
  AOI220     o212(.A0(ori_ori_n228_), .A1(ori_ori_n227_), .B0(ori_ori_n134_), .B1(ori_ori_n84_), .Y(ori_ori_n229_));
  NA2        o213(.A(x6), .B(ori_ori_n46_), .Y(ori_ori_n230_));
  OAI210     o214(.A0(ori_ori_n112_), .A1(ori_ori_n76_), .B0(x4), .Y(ori_ori_n231_));
  AOI210     o215(.A0(ori_ori_n231_), .A1(ori_ori_n230_), .B0(ori_ori_n75_), .Y(ori_ori_n232_));
  NO2        o216(.A(ori_ori_n60_), .B(x6), .Y(ori_ori_n233_));
  NO2        o217(.A(ori_ori_n155_), .B(ori_ori_n41_), .Y(ori_ori_n234_));
  OAI210     o218(.A0(ori_ori_n234_), .A1(ori_ori_n211_), .B0(ori_ori_n233_), .Y(ori_ori_n235_));
  NA2        o219(.A(ori_ori_n193_), .B(ori_ori_n128_), .Y(ori_ori_n236_));
  NA3        o220(.A(ori_ori_n202_), .B(ori_ori_n123_), .C(x6), .Y(ori_ori_n237_));
  OAI210     o221(.A0(ori_ori_n85_), .A1(ori_ori_n34_), .B0(ori_ori_n65_), .Y(ori_ori_n238_));
  NA4        o222(.A(ori_ori_n238_), .B(ori_ori_n237_), .C(ori_ori_n236_), .D(ori_ori_n235_), .Y(ori_ori_n239_));
  OAI210     o223(.A0(ori_ori_n239_), .A1(ori_ori_n232_), .B0(x2), .Y(ori_ori_n240_));
  NA3        o224(.A(ori_ori_n240_), .B(ori_ori_n229_), .C(ori_ori_n225_), .Y(ori_ori_n241_));
  AOI210     o225(.A0(ori_ori_n216_), .A1(x8), .B0(ori_ori_n241_), .Y(ori_ori_n242_));
  NO2        o226(.A(ori_ori_n85_), .B(x3), .Y(ori_ori_n243_));
  NA2        o227(.A(ori_ori_n243_), .B(ori_ori_n200_), .Y(ori_ori_n244_));
  NO2        o228(.A(ori_ori_n83_), .B(ori_ori_n24_), .Y(ori_ori_n245_));
  AOI210     o229(.A0(ori_ori_n220_), .A1(ori_ori_n150_), .B0(ori_ori_n245_), .Y(ori_ori_n246_));
  AOI210     o230(.A0(ori_ori_n246_), .A1(ori_ori_n244_), .B0(x2), .Y(ori_ori_n247_));
  NO2        o231(.A(x4), .B(ori_ori_n52_), .Y(ori_ori_n248_));
  AOI220     o232(.A0(ori_ori_n200_), .A1(ori_ori_n184_), .B0(ori_ori_n248_), .B1(ori_ori_n65_), .Y(ori_ori_n249_));
  NA2        o233(.A(ori_ori_n60_), .B(x6), .Y(ori_ori_n250_));
  NA3        o234(.A(ori_ori_n24_), .B(x3), .C(x2), .Y(ori_ori_n251_));
  AOI210     o235(.A0(ori_ori_n251_), .A1(ori_ori_n133_), .B0(ori_ori_n250_), .Y(ori_ori_n252_));
  NA2        o236(.A(ori_ori_n41_), .B(ori_ori_n17_), .Y(ori_ori_n253_));
  NO2        o237(.A(ori_ori_n253_), .B(ori_ori_n24_), .Y(ori_ori_n254_));
  OAI210     o238(.A0(ori_ori_n254_), .A1(ori_ori_n252_), .B0(ori_ori_n114_), .Y(ori_ori_n255_));
  NA2        o239(.A(ori_ori_n202_), .B(x6), .Y(ori_ori_n256_));
  NO2        o240(.A(ori_ori_n202_), .B(x6), .Y(ori_ori_n257_));
  NAi21      o241(.An(ori_ori_n158_), .B(ori_ori_n257_), .Y(ori_ori_n258_));
  NA3        o242(.A(ori_ori_n258_), .B(ori_ori_n256_), .C(ori_ori_n138_), .Y(ori_ori_n259_));
  NA4        o243(.A(ori_ori_n259_), .B(ori_ori_n255_), .C(ori_ori_n249_), .D(ori_ori_n147_), .Y(ori_ori_n260_));
  NA2        o244(.A(ori_ori_n193_), .B(ori_ori_n219_), .Y(ori_ori_n261_));
  NO2        o245(.A(x9), .B(x6), .Y(ori_ori_n262_));
  NO2        o246(.A(ori_ori_n133_), .B(ori_ori_n18_), .Y(ori_ori_n263_));
  NAi21      o247(.An(ori_ori_n263_), .B(ori_ori_n251_), .Y(ori_ori_n264_));
  NAi21      o248(.An(x1), .B(x4), .Y(ori_ori_n265_));
  AOI210     o249(.A0(x3), .A1(x2), .B0(ori_ori_n46_), .Y(ori_ori_n266_));
  OAI210     o250(.A0(ori_ori_n133_), .A1(x3), .B0(ori_ori_n266_), .Y(ori_ori_n267_));
  AOI220     o251(.A0(ori_ori_n267_), .A1(ori_ori_n265_), .B0(ori_ori_n264_), .B1(ori_ori_n262_), .Y(ori_ori_n268_));
  NA2        o252(.A(ori_ori_n268_), .B(ori_ori_n261_), .Y(ori_ori_n269_));
  NA2        o253(.A(ori_ori_n60_), .B(x2), .Y(ori_ori_n270_));
  NO2        o254(.A(ori_ori_n270_), .B(ori_ori_n261_), .Y(ori_ori_n271_));
  NA2        o255(.A(x6), .B(x2), .Y(ori_ori_n272_));
  NO2        o256(.A(ori_ori_n173_), .B(ori_ori_n44_), .Y(ori_ori_n273_));
  OAI210     o257(.A0(ori_ori_n273_), .A1(ori_ori_n271_), .B0(ori_ori_n269_), .Y(ori_ori_n274_));
  NO2        o258(.A(x3), .B(ori_ori_n199_), .Y(ori_ori_n275_));
  NA2        o259(.A(x4), .B(x0), .Y(ori_ori_n276_));
  NA2        o260(.A(ori_ori_n275_), .B(ori_ori_n40_), .Y(ori_ori_n277_));
  AOI210     o261(.A0(ori_ori_n277_), .A1(ori_ori_n274_), .B0(x8), .Y(ori_ori_n278_));
  INV        o262(.A(ori_ori_n250_), .Y(ori_ori_n279_));
  OAI210     o263(.A0(ori_ori_n263_), .A1(ori_ori_n210_), .B0(ori_ori_n279_), .Y(ori_ori_n280_));
  OAI210     o264(.A0(x0), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n281_));
  AOI210     o265(.A0(ori_ori_n281_), .A1(ori_ori_n280_), .B0(ori_ori_n226_), .Y(ori_ori_n282_));
  NO4        o266(.A(ori_ori_n282_), .B(ori_ori_n278_), .C(ori_ori_n260_), .D(ori_ori_n247_), .Y(ori_ori_n283_));
  NO2        o267(.A(ori_ori_n158_), .B(x1), .Y(ori_ori_n284_));
  NO3        o268(.A(ori_ori_n284_), .B(x3), .C(ori_ori_n34_), .Y(ori_ori_n285_));
  OAI210     o269(.A0(ori_ori_n285_), .A1(ori_ori_n257_), .B0(x2), .Y(ori_ori_n286_));
  OAI210     o270(.A0(x0), .A1(x6), .B0(ori_ori_n42_), .Y(ori_ori_n287_));
  AOI210     o271(.A0(ori_ori_n287_), .A1(ori_ori_n286_), .B0(ori_ori_n183_), .Y(ori_ori_n288_));
  NOi21      o272(.An(ori_ori_n272_), .B(ori_ori_n17_), .Y(ori_ori_n289_));
  NA3        o273(.A(ori_ori_n289_), .B(ori_ori_n210_), .C(ori_ori_n38_), .Y(ori_ori_n290_));
  AOI210     o274(.A0(ori_ori_n34_), .A1(ori_ori_n52_), .B0(x0), .Y(ori_ori_n291_));
  NA3        o275(.A(ori_ori_n291_), .B(ori_ori_n156_), .C(ori_ori_n31_), .Y(ori_ori_n292_));
  NA2        o276(.A(x3), .B(x2), .Y(ori_ori_n293_));
  AOI220     o277(.A0(ori_ori_n293_), .A1(ori_ori_n226_), .B0(ori_ori_n292_), .B1(ori_ori_n290_), .Y(ori_ori_n294_));
  NAi21      o278(.An(x4), .B(x0), .Y(ori_ori_n295_));
  NO3        o279(.A(ori_ori_n295_), .B(ori_ori_n42_), .C(x2), .Y(ori_ori_n296_));
  OAI210     o280(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n296_), .Y(ori_ori_n297_));
  OAI220     o281(.A0(ori_ori_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n298_));
  NO2        o282(.A(x9), .B(x8), .Y(ori_ori_n299_));
  NA3        o283(.A(ori_ori_n299_), .B(ori_ori_n34_), .C(ori_ori_n52_), .Y(ori_ori_n300_));
  OAI210     o284(.A0(ori_ori_n291_), .A1(ori_ori_n289_), .B0(ori_ori_n300_), .Y(ori_ori_n301_));
  AOI220     o285(.A0(ori_ori_n301_), .A1(ori_ori_n79_), .B0(ori_ori_n298_), .B1(ori_ori_n30_), .Y(ori_ori_n302_));
  AOI210     o286(.A0(ori_ori_n302_), .A1(ori_ori_n297_), .B0(ori_ori_n24_), .Y(ori_ori_n303_));
  NA3        o287(.A(ori_ori_n34_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n304_));
  OAI210     o288(.A0(ori_ori_n291_), .A1(ori_ori_n289_), .B0(ori_ori_n304_), .Y(ori_ori_n305_));
  INV        o289(.A(ori_ori_n211_), .Y(ori_ori_n306_));
  NA2        o290(.A(ori_ori_n34_), .B(ori_ori_n41_), .Y(ori_ori_n307_));
  OR2        o291(.A(ori_ori_n307_), .B(ori_ori_n276_), .Y(ori_ori_n308_));
  OAI220     o292(.A0(ori_ori_n308_), .A1(ori_ori_n155_), .B0(ori_ori_n230_), .B1(ori_ori_n306_), .Y(ori_ori_n309_));
  AO210      o293(.A0(ori_ori_n305_), .A1(ori_ori_n142_), .B0(ori_ori_n309_), .Y(ori_ori_n310_));
  NO4        o294(.A(ori_ori_n310_), .B(ori_ori_n303_), .C(ori_ori_n294_), .D(ori_ori_n288_), .Y(ori_ori_n311_));
  OAI210     o295(.A0(ori_ori_n283_), .A1(ori_ori_n242_), .B0(ori_ori_n311_), .Y(ori04));
  NO2        o296(.A(x2), .B(x1), .Y(ori_ori_n313_));
  OAI210     o297(.A0(ori_ori_n253_), .A1(ori_ori_n313_), .B0(ori_ori_n34_), .Y(ori_ori_n314_));
  NO2        o298(.A(ori_ori_n313_), .B(ori_ori_n295_), .Y(ori_ori_n315_));
  AOI210     o299(.A0(ori_ori_n60_), .A1(x4), .B0(ori_ori_n106_), .Y(ori_ori_n316_));
  OAI210     o300(.A0(ori_ori_n316_), .A1(ori_ori_n315_), .B0(ori_ori_n243_), .Y(ori_ori_n317_));
  NO2        o301(.A(ori_ori_n270_), .B(ori_ori_n83_), .Y(ori_ori_n318_));
  NO2        o302(.A(ori_ori_n318_), .B(ori_ori_n34_), .Y(ori_ori_n319_));
  NO2        o303(.A(ori_ori_n293_), .B(ori_ori_n201_), .Y(ori_ori_n320_));
  NA2        o304(.A(x9), .B(x0), .Y(ori_ori_n321_));
  AOI210     o305(.A0(ori_ori_n83_), .A1(ori_ori_n73_), .B0(ori_ori_n321_), .Y(ori_ori_n322_));
  OAI210     o306(.A0(ori_ori_n322_), .A1(ori_ori_n320_), .B0(ori_ori_n85_), .Y(ori_ori_n323_));
  NA3        o307(.A(ori_ori_n323_), .B(ori_ori_n319_), .C(ori_ori_n317_), .Y(ori_ori_n324_));
  NA2        o308(.A(ori_ori_n324_), .B(ori_ori_n314_), .Y(ori_ori_n325_));
  NO2        o309(.A(ori_ori_n204_), .B(ori_ori_n107_), .Y(ori_ori_n326_));
  NO3        o310(.A(ori_ori_n250_), .B(ori_ori_n113_), .C(ori_ori_n18_), .Y(ori_ori_n327_));
  NO2        o311(.A(ori_ori_n327_), .B(ori_ori_n326_), .Y(ori_ori_n328_));
  OAI210     o312(.A0(ori_ori_n111_), .A1(ori_ori_n100_), .B0(ori_ori_n171_), .Y(ori_ori_n329_));
  NA3        o313(.A(ori_ori_n329_), .B(x6), .C(x3), .Y(ori_ori_n330_));
  AOI210     o314(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n331_));
  OAI220     o315(.A0(ori_ori_n331_), .A1(ori_ori_n307_), .B0(ori_ori_n270_), .B1(ori_ori_n304_), .Y(ori_ori_n332_));
  INV        o316(.A(ori_ori_n332_), .Y(ori_ori_n333_));
  NA2        o317(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n334_));
  NA2        o318(.A(ori_ori_n318_), .B(ori_ori_n85_), .Y(ori_ori_n335_));
  NA4        o319(.A(ori_ori_n335_), .B(ori_ori_n333_), .C(ori_ori_n330_), .D(ori_ori_n328_), .Y(ori_ori_n336_));
  OAI210     o320(.A0(ori_ori_n105_), .A1(x3), .B0(ori_ori_n296_), .Y(ori_ori_n337_));
  NA2        o321(.A(ori_ori_n209_), .B(ori_ori_n80_), .Y(ori_ori_n338_));
  NA3        o322(.A(ori_ori_n338_), .B(ori_ori_n337_), .C(ori_ori_n147_), .Y(ori_ori_n339_));
  AOI210     o323(.A0(ori_ori_n336_), .A1(x4), .B0(ori_ori_n339_), .Y(ori_ori_n340_));
  NA3        o324(.A(ori_ori_n315_), .B(ori_ori_n204_), .C(ori_ori_n85_), .Y(ori_ori_n341_));
  NOi21      o325(.An(x4), .B(x0), .Y(ori_ori_n342_));
  XO2        o326(.A(x4), .B(x0), .Y(ori_ori_n343_));
  OAI210     o327(.A0(ori_ori_n343_), .A1(ori_ori_n110_), .B0(ori_ori_n265_), .Y(ori_ori_n344_));
  AOI220     o328(.A0(ori_ori_n344_), .A1(x8), .B0(ori_ori_n342_), .B1(ori_ori_n86_), .Y(ori_ori_n345_));
  AOI210     o329(.A0(ori_ori_n345_), .A1(ori_ori_n341_), .B0(x3), .Y(ori_ori_n346_));
  INV        o330(.A(ori_ori_n86_), .Y(ori_ori_n347_));
  NO2        o331(.A(ori_ori_n85_), .B(x4), .Y(ori_ori_n348_));
  AOI220     o332(.A0(ori_ori_n348_), .A1(ori_ori_n42_), .B0(ori_ori_n118_), .B1(ori_ori_n347_), .Y(ori_ori_n349_));
  NO3        o333(.A(ori_ori_n343_), .B(ori_ori_n158_), .C(x2), .Y(ori_ori_n350_));
  NO3        o334(.A(ori_ori_n222_), .B(ori_ori_n27_), .C(ori_ori_n23_), .Y(ori_ori_n351_));
  NO2        o335(.A(ori_ori_n351_), .B(ori_ori_n350_), .Y(ori_ori_n352_));
  NA4        o336(.A(ori_ori_n352_), .B(ori_ori_n349_), .C(ori_ori_n218_), .D(x6), .Y(ori_ori_n353_));
  OAI220     o337(.A0(ori_ori_n295_), .A1(ori_ori_n83_), .B0(ori_ori_n176_), .B1(ori_ori_n85_), .Y(ori_ori_n354_));
  NO2        o338(.A(ori_ori_n41_), .B(x0), .Y(ori_ori_n355_));
  OR2        o339(.A(ori_ori_n348_), .B(ori_ori_n355_), .Y(ori_ori_n356_));
  NO2        o340(.A(ori_ori_n144_), .B(ori_ori_n100_), .Y(ori_ori_n357_));
  AOI220     o341(.A0(ori_ori_n357_), .A1(ori_ori_n356_), .B0(ori_ori_n354_), .B1(ori_ori_n59_), .Y(ori_ori_n358_));
  NO2        o342(.A(ori_ori_n144_), .B(ori_ori_n78_), .Y(ori_ori_n359_));
  NO2        o343(.A(ori_ori_n33_), .B(x2), .Y(ori_ori_n360_));
  NOi21      o344(.An(ori_ori_n114_), .B(ori_ori_n26_), .Y(ori_ori_n361_));
  AOI210     o345(.A0(ori_ori_n360_), .A1(ori_ori_n359_), .B0(ori_ori_n361_), .Y(ori_ori_n362_));
  OAI210     o346(.A0(ori_ori_n358_), .A1(ori_ori_n60_), .B0(ori_ori_n362_), .Y(ori_ori_n363_));
  OAI220     o347(.A0(ori_ori_n363_), .A1(x6), .B0(ori_ori_n353_), .B1(ori_ori_n346_), .Y(ori_ori_n364_));
  OAI210     o348(.A0(ori_ori_n61_), .A1(ori_ori_n46_), .B0(ori_ori_n40_), .Y(ori_ori_n365_));
  OAI210     o349(.A0(ori_ori_n365_), .A1(ori_ori_n85_), .B0(ori_ori_n308_), .Y(ori_ori_n366_));
  AOI210     o350(.A0(ori_ori_n366_), .A1(ori_ori_n18_), .B0(ori_ori_n147_), .Y(ori_ori_n367_));
  AO220      o351(.A0(ori_ori_n367_), .A1(ori_ori_n364_), .B0(ori_ori_n340_), .B1(ori_ori_n325_), .Y(ori_ori_n368_));
  NA2        o352(.A(ori_ori_n360_), .B(x6), .Y(ori_ori_n369_));
  AOI210     o353(.A0(x6), .A1(x1), .B0(ori_ori_n146_), .Y(ori_ori_n370_));
  NA2        o354(.A(ori_ori_n348_), .B(x0), .Y(ori_ori_n371_));
  NA2        o355(.A(ori_ori_n80_), .B(x6), .Y(ori_ori_n372_));
  OAI210     o356(.A0(ori_ori_n371_), .A1(ori_ori_n370_), .B0(ori_ori_n372_), .Y(ori_ori_n373_));
  AOI220     o357(.A0(ori_ori_n373_), .A1(ori_ori_n369_), .B0(ori_ori_n212_), .B1(ori_ori_n47_), .Y(ori_ori_n374_));
  NA2        o358(.A(ori_ori_n374_), .B(ori_ori_n368_), .Y(ori_ori_n375_));
  AOI210     o359(.A0(ori_ori_n195_), .A1(x8), .B0(ori_ori_n105_), .Y(ori_ori_n376_));
  NA2        o360(.A(ori_ori_n376_), .B(ori_ori_n334_), .Y(ori_ori_n377_));
  NA3        o361(.A(ori_ori_n377_), .B(ori_ori_n192_), .C(ori_ori_n147_), .Y(ori_ori_n378_));
  NA3        o362(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n379_));
  NA2        o363(.A(ori_ori_n217_), .B(x0), .Y(ori_ori_n380_));
  OAI220     o364(.A0(ori_ori_n380_), .A1(ori_ori_n204_), .B0(ori_ori_n379_), .B1(ori_ori_n347_), .Y(ori_ori_n381_));
  INV        o365(.A(ori_ori_n381_), .Y(ori_ori_n382_));
  AOI210     o366(.A0(ori_ori_n382_), .A1(ori_ori_n378_), .B0(ori_ori_n24_), .Y(ori_ori_n383_));
  OAI210     o367(.A0(ori_ori_n192_), .A1(ori_ori_n66_), .B0(ori_ori_n201_), .Y(ori_ori_n384_));
  NA3        o368(.A(ori_ori_n195_), .B(ori_ori_n219_), .C(x8), .Y(ori_ori_n385_));
  AOI210     o369(.A0(ori_ori_n385_), .A1(ori_ori_n384_), .B0(ori_ori_n24_), .Y(ori_ori_n386_));
  AOI210     o370(.A0(ori_ori_n113_), .A1(ori_ori_n111_), .B0(ori_ori_n40_), .Y(ori_ori_n387_));
  NOi31      o371(.An(ori_ori_n387_), .B(ori_ori_n355_), .C(ori_ori_n177_), .Y(ori_ori_n388_));
  OAI210     o372(.A0(ori_ori_n388_), .A1(ori_ori_n386_), .B0(ori_ori_n143_), .Y(ori_ori_n389_));
  NAi31      o373(.An(ori_ori_n48_), .B(ori_ori_n284_), .C(ori_ori_n172_), .Y(ori_ori_n390_));
  NA2        o374(.A(ori_ori_n390_), .B(ori_ori_n389_), .Y(ori_ori_n391_));
  OAI210     o375(.A0(ori_ori_n391_), .A1(ori_ori_n383_), .B0(x6), .Y(ori_ori_n392_));
  OAI210     o376(.A0(ori_ori_n158_), .A1(ori_ori_n46_), .B0(ori_ori_n129_), .Y(ori_ori_n393_));
  NA3        o377(.A(ori_ori_n53_), .B(ori_ori_n36_), .C(ori_ori_n30_), .Y(ori_ori_n394_));
  AOI220     o378(.A0(ori_ori_n394_), .A1(ori_ori_n393_), .B0(ori_ori_n38_), .B1(ori_ori_n31_), .Y(ori_ori_n395_));
  NO2        o379(.A(ori_ori_n147_), .B(x0), .Y(ori_ori_n396_));
  AOI220     o380(.A0(ori_ori_n396_), .A1(ori_ori_n217_), .B0(ori_ori_n192_), .B1(ori_ori_n147_), .Y(ori_ori_n397_));
  AOI210     o381(.A0(ori_ori_n120_), .A1(ori_ori_n248_), .B0(x1), .Y(ori_ori_n398_));
  OAI210     o382(.A0(ori_ori_n397_), .A1(x8), .B0(ori_ori_n398_), .Y(ori_ori_n399_));
  NAi31      o383(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n400_));
  OAI210     o384(.A0(ori_ori_n400_), .A1(x4), .B0(ori_ori_n159_), .Y(ori_ori_n401_));
  NA3        o385(.A(ori_ori_n401_), .B(ori_ori_n141_), .C(x9), .Y(ori_ori_n402_));
  NO4        o386(.A(ori_ori_n119_), .B(ori_ori_n295_), .C(x9), .D(x2), .Y(ori_ori_n403_));
  NOi21      o387(.An(ori_ori_n117_), .B(ori_ori_n176_), .Y(ori_ori_n404_));
  NO3        o388(.A(ori_ori_n404_), .B(ori_ori_n403_), .C(ori_ori_n18_), .Y(ori_ori_n405_));
  NO3        o389(.A(x9), .B(ori_ori_n147_), .C(x0), .Y(ori_ori_n406_));
  AOI220     o390(.A0(ori_ori_n406_), .A1(ori_ori_n243_), .B0(ori_ori_n359_), .B1(ori_ori_n147_), .Y(ori_ori_n407_));
  NA4        o391(.A(ori_ori_n407_), .B(ori_ori_n405_), .C(ori_ori_n402_), .D(ori_ori_n48_), .Y(ori_ori_n408_));
  OAI210     o392(.A0(ori_ori_n399_), .A1(ori_ori_n395_), .B0(ori_ori_n408_), .Y(ori_ori_n409_));
  NOi31      o393(.An(ori_ori_n396_), .B(ori_ori_n31_), .C(x8), .Y(ori_ori_n410_));
  AOI210     o394(.A0(ori_ori_n36_), .A1(x9), .B0(ori_ori_n127_), .Y(ori_ori_n411_));
  NO3        o395(.A(ori_ori_n411_), .B(ori_ori_n117_), .C(ori_ori_n41_), .Y(ori_ori_n412_));
  NOi31      o396(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n413_));
  AOI210     o397(.A0(ori_ori_n265_), .A1(ori_ori_n58_), .B0(ori_ori_n116_), .Y(ori_ori_n414_));
  NO2        o398(.A(ori_ori_n414_), .B(x3), .Y(ori_ori_n415_));
  NO3        o399(.A(ori_ori_n415_), .B(ori_ori_n412_), .C(x2), .Y(ori_ori_n416_));
  OAI220     o400(.A0(ori_ori_n343_), .A1(ori_ori_n299_), .B0(ori_ori_n295_), .B1(ori_ori_n41_), .Y(ori_ori_n417_));
  AOI210     o401(.A0(x9), .A1(ori_ori_n46_), .B0(ori_ori_n379_), .Y(ori_ori_n418_));
  AOI220     o402(.A0(ori_ori_n418_), .A1(ori_ori_n85_), .B0(ori_ori_n417_), .B1(ori_ori_n147_), .Y(ori_ori_n419_));
  NO2        o403(.A(ori_ori_n419_), .B(ori_ori_n52_), .Y(ori_ori_n420_));
  NO3        o404(.A(ori_ori_n420_), .B(ori_ori_n416_), .C(ori_ori_n410_), .Y(ori_ori_n421_));
  AOI210     o405(.A0(ori_ori_n421_), .A1(ori_ori_n409_), .B0(ori_ori_n24_), .Y(ori_ori_n422_));
  NA4        o406(.A(ori_ori_n30_), .B(ori_ori_n85_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n423_));
  NO3        o407(.A(ori_ori_n60_), .B(x4), .C(x1), .Y(ori_ori_n424_));
  NO3        o408(.A(ori_ori_n66_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n425_));
  AOI220     o409(.A0(ori_ori_n425_), .A1(ori_ori_n266_), .B0(ori_ori_n424_), .B1(ori_ori_n387_), .Y(ori_ori_n426_));
  NO2        o410(.A(ori_ori_n426_), .B(ori_ori_n97_), .Y(ori_ori_n427_));
  NO3        o411(.A(ori_ori_n270_), .B(ori_ori_n171_), .C(ori_ori_n38_), .Y(ori_ori_n428_));
  OAI210     o412(.A0(ori_ori_n428_), .A1(ori_ori_n427_), .B0(x7), .Y(ori_ori_n429_));
  NA2        o413(.A(ori_ori_n222_), .B(x7), .Y(ori_ori_n430_));
  NA3        o414(.A(ori_ori_n430_), .B(ori_ori_n146_), .C(ori_ori_n128_), .Y(ori_ori_n431_));
  NA3        o415(.A(ori_ori_n431_), .B(ori_ori_n429_), .C(ori_ori_n423_), .Y(ori_ori_n432_));
  OAI210     o416(.A0(ori_ori_n432_), .A1(ori_ori_n422_), .B0(ori_ori_n34_), .Y(ori_ori_n433_));
  NO2        o417(.A(ori_ori_n406_), .B(ori_ori_n201_), .Y(ori_ori_n434_));
  NO4        o418(.A(ori_ori_n434_), .B(ori_ori_n75_), .C(x4), .D(ori_ori_n52_), .Y(ori_ori_n435_));
  NA2        o419(.A(ori_ori_n253_), .B(ori_ori_n21_), .Y(ori_ori_n436_));
  NO2        o420(.A(ori_ori_n155_), .B(ori_ori_n129_), .Y(ori_ori_n437_));
  NA2        o421(.A(ori_ori_n437_), .B(ori_ori_n436_), .Y(ori_ori_n438_));
  AOI210     o422(.A0(ori_ori_n438_), .A1(ori_ori_n162_), .B0(ori_ori_n27_), .Y(ori_ori_n439_));
  AOI220     o423(.A0(ori_ori_n355_), .A1(ori_ori_n85_), .B0(ori_ori_n144_), .B1(ori_ori_n195_), .Y(ori_ori_n440_));
  NA3        o424(.A(ori_ori_n440_), .B(ori_ori_n400_), .C(ori_ori_n83_), .Y(ori_ori_n441_));
  NA2        o425(.A(ori_ori_n441_), .B(ori_ori_n172_), .Y(ori_ori_n442_));
  OAI220     o426(.A0(x3), .A1(ori_ori_n67_), .B0(ori_ori_n155_), .B1(ori_ori_n41_), .Y(ori_ori_n443_));
  NA2        o427(.A(x3), .B(ori_ori_n52_), .Y(ori_ori_n444_));
  OAI210     o428(.A0(ori_ori_n143_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n445_));
  NO3        o429(.A(ori_ori_n413_), .B(x3), .C(ori_ori_n52_), .Y(ori_ori_n446_));
  NA2        o430(.A(ori_ori_n446_), .B(ori_ori_n445_), .Y(ori_ori_n447_));
  OAI210     o431(.A0(ori_ori_n148_), .A1(ori_ori_n444_), .B0(ori_ori_n447_), .Y(ori_ori_n448_));
  AOI220     o432(.A0(ori_ori_n448_), .A1(x0), .B0(ori_ori_n443_), .B1(ori_ori_n129_), .Y(ori_ori_n449_));
  AOI210     o433(.A0(ori_ori_n449_), .A1(ori_ori_n442_), .B0(ori_ori_n230_), .Y(ori_ori_n450_));
  NO3        o434(.A(ori_ori_n450_), .B(ori_ori_n439_), .C(ori_ori_n435_), .Y(ori_ori_n451_));
  NA3        o435(.A(ori_ori_n451_), .B(ori_ori_n433_), .C(ori_ori_n392_), .Y(ori_ori_n452_));
  AOI210     o436(.A0(ori_ori_n375_), .A1(ori_ori_n24_), .B0(ori_ori_n452_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO4        m012(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .D(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  AN2        m021(.A(x8), .B(x7), .Y(mai_mai_n38_));
  NA3        m022(.A(mai_mai_n38_), .B(mai_mai_n37_), .C(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m023(.A(x4), .B(x3), .Y(mai_mai_n40_));
  AOI210     m024(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(x2), .B(x0), .Y(mai_mai_n42_));
  INV        m026(.A(x3), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n44_));
  INV        m028(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n46_));
  OAI210     m030(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n42_), .Y(mai_mai_n47_));
  INV        m031(.A(x4), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n49_), .B(x2), .Y(mai_mai_n50_));
  OAI210     m034(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n47_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n38_), .B(mai_mai_n37_), .Y(mai_mai_n52_));
  AOI220     m036(.A0(mai_mai_n52_), .A1(mai_mai_n35_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n53_));
  INV        m037(.A(x2), .Y(mai_mai_n54_));
  NO2        m038(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n55_));
  NA2        m039(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  OAI210     m041(.A0(mai_mai_n53_), .A1(mai_mai_n32_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  NO3        m042(.A(mai_mai_n58_), .B(mai_mai_n51_), .C(mai_mai_n41_), .Y(mai01));
  NA2        m043(.A(x8), .B(x7), .Y(mai_mai_n60_));
  NA2        m044(.A(mai_mai_n43_), .B(x1), .Y(mai_mai_n61_));
  INV        m045(.A(x9), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n62_), .B(mai_mai_n36_), .Y(mai_mai_n63_));
  INV        m047(.A(mai_mai_n63_), .Y(mai_mai_n64_));
  NO2        m048(.A(x7), .B(x6), .Y(mai_mai_n65_));
  NO2        m049(.A(mai_mai_n61_), .B(x5), .Y(mai_mai_n66_));
  NO2        m050(.A(x8), .B(x2), .Y(mai_mai_n67_));
  INV        m051(.A(mai_mai_n67_), .Y(mai_mai_n68_));
  NO2        m052(.A(mai_mai_n68_), .B(x1), .Y(mai_mai_n69_));
  OA210      m053(.A0(mai_mai_n69_), .A1(mai_mai_n66_), .B0(mai_mai_n65_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n44_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n71_));
  OAI210     m055(.A0(mai_mai_n56_), .A1(mai_mai_n20_), .B0(mai_mai_n71_), .Y(mai_mai_n72_));
  NAi31      m056(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n73_));
  OAI220     m057(.A0(mai_mai_n73_), .A1(mai_mai_n43_), .B0(mai_mai_n72_), .B1(mai_mai_n70_), .Y(mai_mai_n74_));
  NA2        m058(.A(mai_mai_n74_), .B(x4), .Y(mai_mai_n75_));
  NA2        m059(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n76_));
  OAI210     m060(.A0(mai_mai_n76_), .A1(mai_mai_n56_), .B0(x0), .Y(mai_mai_n77_));
  NA2        m061(.A(x5), .B(x3), .Y(mai_mai_n78_));
  NO2        m062(.A(x8), .B(x6), .Y(mai_mai_n79_));
  NO4        m063(.A(mai_mai_n79_), .B(mai_mai_n78_), .C(mai_mai_n65_), .D(mai_mai_n54_), .Y(mai_mai_n80_));
  NAi21      m064(.An(x4), .B(x3), .Y(mai_mai_n81_));
  INV        m065(.A(mai_mai_n81_), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(mai_mai_n22_), .Y(mai_mai_n83_));
  NO2        m067(.A(x4), .B(x2), .Y(mai_mai_n84_));
  NO2        m068(.A(mai_mai_n84_), .B(x3), .Y(mai_mai_n85_));
  NO3        m069(.A(mai_mai_n85_), .B(mai_mai_n83_), .C(mai_mai_n18_), .Y(mai_mai_n86_));
  NO3        m070(.A(mai_mai_n86_), .B(mai_mai_n80_), .C(mai_mai_n77_), .Y(mai_mai_n87_));
  NO4        m071(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n43_), .D(x1), .Y(mai_mai_n88_));
  NA2        m072(.A(mai_mai_n62_), .B(mai_mai_n48_), .Y(mai_mai_n89_));
  INV        m073(.A(mai_mai_n89_), .Y(mai_mai_n90_));
  NA2        m074(.A(mai_mai_n88_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  NA2        m075(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n92_), .B(mai_mai_n25_), .Y(mai_mai_n93_));
  INV        m077(.A(x8), .Y(mai_mai_n94_));
  NA2        m078(.A(x2), .B(x1), .Y(mai_mai_n95_));
  INV        m079(.A(mai_mai_n93_), .Y(mai_mai_n96_));
  NO2        m080(.A(mai_mai_n96_), .B(mai_mai_n26_), .Y(mai_mai_n97_));
  AOI210     m081(.A0(mai_mai_n56_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n98_));
  OAI210     m082(.A0(mai_mai_n45_), .A1(mai_mai_n37_), .B0(mai_mai_n48_), .Y(mai_mai_n99_));
  NO3        m083(.A(mai_mai_n99_), .B(mai_mai_n98_), .C(mai_mai_n97_), .Y(mai_mai_n100_));
  NA2        m084(.A(x4), .B(mai_mai_n43_), .Y(mai_mai_n101_));
  NO2        m085(.A(mai_mai_n48_), .B(mai_mai_n54_), .Y(mai_mai_n102_));
  OAI210     m086(.A0(mai_mai_n102_), .A1(mai_mai_n43_), .B0(mai_mai_n18_), .Y(mai_mai_n103_));
  AOI210     m087(.A0(mai_mai_n101_), .A1(mai_mai_n52_), .B0(mai_mai_n103_), .Y(mai_mai_n104_));
  NO2        m088(.A(x3), .B(x2), .Y(mai_mai_n105_));
  NA3        m089(.A(mai_mai_n105_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n106_));
  AOI210     m090(.A0(x8), .A1(x6), .B0(mai_mai_n106_), .Y(mai_mai_n107_));
  NA2        m091(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n108_));
  OAI210     m092(.A0(mai_mai_n108_), .A1(mai_mai_n40_), .B0(mai_mai_n17_), .Y(mai_mai_n109_));
  NO4        m093(.A(mai_mai_n109_), .B(mai_mai_n107_), .C(mai_mai_n104_), .D(mai_mai_n100_), .Y(mai_mai_n110_));
  AO220      m094(.A0(mai_mai_n110_), .A1(mai_mai_n91_), .B0(mai_mai_n87_), .B1(mai_mai_n75_), .Y(mai02));
  NO2        m095(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n112_));
  NO2        m096(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n113_));
  NA2        m097(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n114_));
  NA2        m098(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n115_));
  OAI210     m099(.A0(mai_mai_n89_), .A1(mai_mai_n114_), .B0(mai_mai_n115_), .Y(mai_mai_n116_));
  AOI220     m100(.A0(mai_mai_n116_), .A1(mai_mai_n113_), .B0(mai_mai_n112_), .B1(x4), .Y(mai_mai_n117_));
  NO3        m101(.A(mai_mai_n117_), .B(x7), .C(x5), .Y(mai_mai_n118_));
  NA2        m102(.A(x9), .B(x2), .Y(mai_mai_n119_));
  OR2        m103(.A(x8), .B(x0), .Y(mai_mai_n120_));
  INV        m104(.A(mai_mai_n120_), .Y(mai_mai_n121_));
  NAi21      m105(.An(x2), .B(x8), .Y(mai_mai_n122_));
  INV        m106(.A(mai_mai_n122_), .Y(mai_mai_n123_));
  OAI220     m107(.A0(mai_mai_n123_), .A1(mai_mai_n121_), .B0(mai_mai_n119_), .B1(x7), .Y(mai_mai_n124_));
  NO2        m108(.A(x4), .B(x1), .Y(mai_mai_n125_));
  NA3        m109(.A(mai_mai_n125_), .B(mai_mai_n124_), .C(mai_mai_n60_), .Y(mai_mai_n126_));
  NOi21      m110(.An(x0), .B(x1), .Y(mai_mai_n127_));
  NOi21      m111(.An(x0), .B(x4), .Y(mai_mai_n128_));
  NAi21      m112(.An(x8), .B(x7), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n129_), .B(mai_mai_n62_), .Y(mai_mai_n130_));
  NA2        m114(.A(mai_mai_n130_), .B(mai_mai_n128_), .Y(mai_mai_n131_));
  AOI210     m115(.A0(mai_mai_n131_), .A1(mai_mai_n126_), .B0(mai_mai_n78_), .Y(mai_mai_n132_));
  NO2        m116(.A(x5), .B(mai_mai_n48_), .Y(mai_mai_n133_));
  NA2        m117(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n134_));
  AOI210     m118(.A0(mai_mai_n134_), .A1(mai_mai_n108_), .B0(mai_mai_n115_), .Y(mai_mai_n135_));
  OAI210     m119(.A0(mai_mai_n135_), .A1(mai_mai_n35_), .B0(mai_mai_n133_), .Y(mai_mai_n136_));
  NAi21      m120(.An(x0), .B(x4), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n137_), .B(x1), .Y(mai_mai_n138_));
  NO2        m122(.A(x7), .B(x0), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n84_), .B(mai_mai_n102_), .Y(mai_mai_n140_));
  NO2        m124(.A(mai_mai_n140_), .B(x3), .Y(mai_mai_n141_));
  OAI210     m125(.A0(mai_mai_n139_), .A1(mai_mai_n138_), .B0(mai_mai_n141_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n21_), .B(mai_mai_n43_), .Y(mai_mai_n143_));
  NA2        m127(.A(x5), .B(x0), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n145_));
  NA3        m129(.A(mai_mai_n145_), .B(mai_mai_n144_), .C(mai_mai_n143_), .Y(mai_mai_n146_));
  NA4        m130(.A(mai_mai_n146_), .B(mai_mai_n142_), .C(mai_mai_n136_), .D(mai_mai_n36_), .Y(mai_mai_n147_));
  NO3        m131(.A(mai_mai_n147_), .B(mai_mai_n132_), .C(mai_mai_n118_), .Y(mai_mai_n148_));
  NO3        m132(.A(mai_mai_n78_), .B(mai_mai_n76_), .C(mai_mai_n24_), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n150_));
  NA2        m134(.A(x7), .B(x3), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n101_), .B(x5), .Y(mai_mai_n152_));
  NO2        m136(.A(x9), .B(x7), .Y(mai_mai_n153_));
  NOi21      m137(.An(x8), .B(x0), .Y(mai_mai_n154_));
  OA210      m138(.A0(mai_mai_n153_), .A1(x1), .B0(mai_mai_n154_), .Y(mai_mai_n155_));
  NO2        m139(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n156_));
  INV        m140(.A(x7), .Y(mai_mai_n157_));
  NA2        m141(.A(mai_mai_n157_), .B(mai_mai_n18_), .Y(mai_mai_n158_));
  AOI220     m142(.A0(mai_mai_n158_), .A1(mai_mai_n156_), .B0(mai_mai_n112_), .B1(mai_mai_n38_), .Y(mai_mai_n159_));
  NO2        m143(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n160_), .B(mai_mai_n128_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n161_), .B(mai_mai_n159_), .Y(mai_mai_n162_));
  AOI210     m146(.A0(mai_mai_n155_), .A1(mai_mai_n152_), .B0(mai_mai_n162_), .Y(mai_mai_n163_));
  OAI210     m147(.A0(mai_mai_n151_), .A1(mai_mai_n50_), .B0(mai_mai_n163_), .Y(mai_mai_n164_));
  NA2        m148(.A(x5), .B(x1), .Y(mai_mai_n165_));
  INV        m149(.A(mai_mai_n165_), .Y(mai_mai_n166_));
  AOI210     m150(.A0(mai_mai_n166_), .A1(mai_mai_n128_), .B0(mai_mai_n36_), .Y(mai_mai_n167_));
  NAi21      m151(.An(x2), .B(x7), .Y(mai_mai_n168_));
  NO2        m152(.A(mai_mai_n168_), .B(mai_mai_n48_), .Y(mai_mai_n169_));
  NA2        m153(.A(mai_mai_n169_), .B(mai_mai_n66_), .Y(mai_mai_n170_));
  NAi31      m154(.An(mai_mai_n78_), .B(mai_mai_n38_), .C(mai_mai_n35_), .Y(mai_mai_n171_));
  NA3        m155(.A(mai_mai_n171_), .B(mai_mai_n170_), .C(mai_mai_n167_), .Y(mai_mai_n172_));
  NO3        m156(.A(mai_mai_n172_), .B(mai_mai_n164_), .C(mai_mai_n149_), .Y(mai_mai_n173_));
  NO2        m157(.A(mai_mai_n173_), .B(mai_mai_n148_), .Y(mai_mai_n174_));
  NO2        m158(.A(mai_mai_n144_), .B(mai_mai_n140_), .Y(mai_mai_n175_));
  NA2        m159(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n176_));
  NA2        m160(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n177_));
  NA3        m161(.A(mai_mai_n177_), .B(mai_mai_n176_), .C(mai_mai_n24_), .Y(mai_mai_n178_));
  AN2        m162(.A(mai_mai_n178_), .B(mai_mai_n145_), .Y(mai_mai_n179_));
  NA2        m163(.A(x8), .B(x0), .Y(mai_mai_n180_));
  NO2        m164(.A(mai_mai_n157_), .B(mai_mai_n25_), .Y(mai_mai_n181_));
  NO2        m165(.A(mai_mai_n127_), .B(x4), .Y(mai_mai_n182_));
  NA2        m166(.A(mai_mai_n182_), .B(mai_mai_n181_), .Y(mai_mai_n183_));
  AOI210     m167(.A0(mai_mai_n180_), .A1(mai_mai_n134_), .B0(mai_mai_n183_), .Y(mai_mai_n184_));
  NA2        m168(.A(x2), .B(x0), .Y(mai_mai_n185_));
  NA2        m169(.A(x4), .B(x1), .Y(mai_mai_n186_));
  NAi21      m170(.An(mai_mai_n125_), .B(mai_mai_n186_), .Y(mai_mai_n187_));
  NOi31      m171(.An(mai_mai_n187_), .B(mai_mai_n160_), .C(mai_mai_n185_), .Y(mai_mai_n188_));
  NO4        m172(.A(mai_mai_n188_), .B(mai_mai_n184_), .C(mai_mai_n179_), .D(mai_mai_n175_), .Y(mai_mai_n189_));
  NO2        m173(.A(mai_mai_n189_), .B(mai_mai_n43_), .Y(mai_mai_n190_));
  NO2        m174(.A(mai_mai_n178_), .B(mai_mai_n76_), .Y(mai_mai_n191_));
  INV        m175(.A(mai_mai_n133_), .Y(mai_mai_n192_));
  NO2        m176(.A(mai_mai_n108_), .B(mai_mai_n17_), .Y(mai_mai_n193_));
  AOI210     m177(.A0(mai_mai_n35_), .A1(mai_mai_n94_), .B0(mai_mai_n193_), .Y(mai_mai_n194_));
  NO3        m178(.A(mai_mai_n194_), .B(mai_mai_n192_), .C(x7), .Y(mai_mai_n195_));
  NA3        m179(.A(mai_mai_n187_), .B(mai_mai_n192_), .C(mai_mai_n42_), .Y(mai_mai_n196_));
  OAI210     m180(.A0(mai_mai_n177_), .A1(mai_mai_n140_), .B0(mai_mai_n196_), .Y(mai_mai_n197_));
  NO3        m181(.A(mai_mai_n197_), .B(mai_mai_n195_), .C(mai_mai_n191_), .Y(mai_mai_n198_));
  NO2        m182(.A(mai_mai_n198_), .B(x3), .Y(mai_mai_n199_));
  NO3        m183(.A(mai_mai_n199_), .B(mai_mai_n190_), .C(mai_mai_n174_), .Y(mai03));
  NO2        m184(.A(mai_mai_n48_), .B(x3), .Y(mai_mai_n201_));
  NO2        m185(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n202_));
  NO2        m186(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n203_));
  NO2        m187(.A(mai_mai_n78_), .B(x6), .Y(mai_mai_n204_));
  NA2        m188(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n205_));
  NO2        m189(.A(mai_mai_n205_), .B(x4), .Y(mai_mai_n206_));
  NO2        m190(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n207_));
  AO220      m191(.A0(mai_mai_n207_), .A1(mai_mai_n206_), .B0(mai_mai_n204_), .B1(mai_mai_n55_), .Y(mai_mai_n208_));
  INV        m192(.A(mai_mai_n208_), .Y(mai_mai_n209_));
  NA2        m193(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n210_));
  NA2        m194(.A(mai_mai_n205_), .B(mai_mai_n81_), .Y(mai_mai_n211_));
  AOI210     m195(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n185_), .Y(mai_mai_n212_));
  NA2        m196(.A(mai_mai_n212_), .B(mai_mai_n211_), .Y(mai_mai_n213_));
  NO2        m197(.A(x5), .B(x1), .Y(mai_mai_n214_));
  AOI220     m198(.A0(mai_mai_n214_), .A1(mai_mai_n17_), .B0(mai_mai_n105_), .B1(x5), .Y(mai_mai_n215_));
  NO2        m199(.A(mai_mai_n210_), .B(mai_mai_n176_), .Y(mai_mai_n216_));
  NO3        m200(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n217_));
  NO2        m201(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  OAI210     m202(.A0(mai_mai_n215_), .A1(mai_mai_n64_), .B0(mai_mai_n218_), .Y(mai_mai_n219_));
  NA2        m203(.A(mai_mai_n219_), .B(mai_mai_n48_), .Y(mai_mai_n220_));
  NA3        m204(.A(mai_mai_n220_), .B(mai_mai_n213_), .C(mai_mai_n209_), .Y(mai_mai_n221_));
  NO2        m205(.A(mai_mai_n48_), .B(mai_mai_n43_), .Y(mai_mai_n222_));
  NA2        m206(.A(mai_mai_n222_), .B(mai_mai_n19_), .Y(mai_mai_n223_));
  NO2        m207(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n224_));
  NO2        m208(.A(mai_mai_n224_), .B(x6), .Y(mai_mai_n225_));
  NOi21      m209(.An(mai_mai_n84_), .B(mai_mai_n225_), .Y(mai_mai_n226_));
  NA2        m210(.A(mai_mai_n62_), .B(mai_mai_n94_), .Y(mai_mai_n227_));
  NA3        m211(.A(mai_mai_n227_), .B(mai_mai_n224_), .C(x6), .Y(mai_mai_n228_));
  AOI210     m212(.A0(mai_mai_n228_), .A1(mai_mai_n226_), .B0(mai_mai_n157_), .Y(mai_mai_n229_));
  AO210      m213(.A0(mai_mai_n229_), .A1(mai_mai_n223_), .B0(mai_mai_n181_), .Y(mai_mai_n230_));
  NA2        m214(.A(mai_mai_n43_), .B(mai_mai_n54_), .Y(mai_mai_n231_));
  OAI210     m215(.A0(mai_mai_n231_), .A1(mai_mai_n25_), .B0(mai_mai_n177_), .Y(mai_mai_n232_));
  NO2        m216(.A(mai_mai_n186_), .B(x6), .Y(mai_mai_n233_));
  AOI220     m217(.A0(mai_mai_n233_), .A1(mai_mai_n232_), .B0(mai_mai_n145_), .B1(mai_mai_n93_), .Y(mai_mai_n234_));
  NA2        m218(.A(x6), .B(mai_mai_n48_), .Y(mai_mai_n235_));
  OAI210     m219(.A0(mai_mai_n121_), .A1(mai_mai_n79_), .B0(x4), .Y(mai_mai_n236_));
  AOI210     m220(.A0(mai_mai_n236_), .A1(mai_mai_n235_), .B0(mai_mai_n78_), .Y(mai_mai_n237_));
  NO2        m221(.A(mai_mai_n62_), .B(x6), .Y(mai_mai_n238_));
  NO2        m222(.A(mai_mai_n165_), .B(mai_mai_n43_), .Y(mai_mai_n239_));
  OAI210     m223(.A0(mai_mai_n239_), .A1(mai_mai_n216_), .B0(mai_mai_n238_), .Y(mai_mai_n240_));
  NA2        m224(.A(mai_mai_n202_), .B(mai_mai_n138_), .Y(mai_mai_n241_));
  NA3        m225(.A(mai_mai_n210_), .B(mai_mai_n133_), .C(x6), .Y(mai_mai_n242_));
  OAI210     m226(.A0(mai_mai_n94_), .A1(mai_mai_n36_), .B0(mai_mai_n66_), .Y(mai_mai_n243_));
  NA4        m227(.A(mai_mai_n243_), .B(mai_mai_n242_), .C(mai_mai_n241_), .D(mai_mai_n240_), .Y(mai_mai_n244_));
  OAI210     m228(.A0(mai_mai_n244_), .A1(mai_mai_n237_), .B0(x2), .Y(mai_mai_n245_));
  NA3        m229(.A(mai_mai_n245_), .B(mai_mai_n234_), .C(mai_mai_n230_), .Y(mai_mai_n246_));
  AOI210     m230(.A0(mai_mai_n221_), .A1(x8), .B0(mai_mai_n246_), .Y(mai_mai_n247_));
  NO2        m231(.A(mai_mai_n94_), .B(x3), .Y(mai_mai_n248_));
  NA2        m232(.A(mai_mai_n248_), .B(mai_mai_n206_), .Y(mai_mai_n249_));
  NO3        m233(.A(mai_mai_n92_), .B(mai_mai_n79_), .C(mai_mai_n25_), .Y(mai_mai_n250_));
  AOI210     m234(.A0(mai_mai_n225_), .A1(mai_mai_n160_), .B0(mai_mai_n250_), .Y(mai_mai_n251_));
  AOI210     m235(.A0(mai_mai_n251_), .A1(mai_mai_n249_), .B0(x2), .Y(mai_mai_n252_));
  NO2        m236(.A(x4), .B(mai_mai_n54_), .Y(mai_mai_n253_));
  AOI220     m237(.A0(mai_mai_n206_), .A1(mai_mai_n193_), .B0(mai_mai_n253_), .B1(mai_mai_n66_), .Y(mai_mai_n254_));
  NA2        m238(.A(mai_mai_n62_), .B(x6), .Y(mai_mai_n255_));
  NA2        m239(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n256_));
  NO2        m240(.A(mai_mai_n256_), .B(mai_mai_n25_), .Y(mai_mai_n257_));
  NA2        m241(.A(mai_mai_n257_), .B(mai_mai_n125_), .Y(mai_mai_n258_));
  NA2        m242(.A(mai_mai_n210_), .B(x6), .Y(mai_mai_n259_));
  NO2        m243(.A(mai_mai_n210_), .B(x6), .Y(mai_mai_n260_));
  INV        m244(.A(mai_mai_n260_), .Y(mai_mai_n261_));
  NA3        m245(.A(mai_mai_n261_), .B(mai_mai_n259_), .C(mai_mai_n150_), .Y(mai_mai_n262_));
  NA4        m246(.A(mai_mai_n262_), .B(mai_mai_n258_), .C(mai_mai_n254_), .D(mai_mai_n157_), .Y(mai_mai_n263_));
  NO2        m247(.A(mai_mai_n144_), .B(mai_mai_n18_), .Y(mai_mai_n264_));
  NAi21      m248(.An(x1), .B(x4), .Y(mai_mai_n265_));
  AOI210     m249(.A0(x3), .A1(x2), .B0(mai_mai_n48_), .Y(mai_mai_n266_));
  OAI210     m250(.A0(mai_mai_n144_), .A1(x3), .B0(mai_mai_n266_), .Y(mai_mai_n267_));
  NA2        m251(.A(mai_mai_n267_), .B(mai_mai_n265_), .Y(mai_mai_n268_));
  INV        m252(.A(mai_mai_n268_), .Y(mai_mai_n269_));
  NA2        m253(.A(mai_mai_n62_), .B(x2), .Y(mai_mai_n270_));
  NO3        m254(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n271_));
  NA2        m255(.A(mai_mai_n108_), .B(mai_mai_n25_), .Y(mai_mai_n272_));
  NA2        m256(.A(x6), .B(x2), .Y(mai_mai_n273_));
  NO2        m257(.A(mai_mai_n273_), .B(mai_mai_n176_), .Y(mai_mai_n274_));
  AOI210     m258(.A0(mai_mai_n272_), .A1(mai_mai_n271_), .B0(mai_mai_n274_), .Y(mai_mai_n275_));
  OAI220     m259(.A0(mai_mai_n275_), .A1(mai_mai_n43_), .B0(mai_mai_n182_), .B1(mai_mai_n46_), .Y(mai_mai_n276_));
  NA2        m260(.A(mai_mai_n276_), .B(mai_mai_n269_), .Y(mai_mai_n277_));
  NA2        m261(.A(x9), .B(mai_mai_n43_), .Y(mai_mai_n278_));
  NO2        m262(.A(mai_mai_n278_), .B(mai_mai_n205_), .Y(mai_mai_n279_));
  OR3        m263(.A(mai_mai_n279_), .B(mai_mai_n204_), .C(mai_mai_n152_), .Y(mai_mai_n280_));
  NA2        m264(.A(x4), .B(x0), .Y(mai_mai_n281_));
  NO3        m265(.A(mai_mai_n73_), .B(mai_mai_n281_), .C(x6), .Y(mai_mai_n282_));
  AOI210     m266(.A0(mai_mai_n280_), .A1(mai_mai_n42_), .B0(mai_mai_n282_), .Y(mai_mai_n283_));
  AOI210     m267(.A0(mai_mai_n283_), .A1(mai_mai_n277_), .B0(x8), .Y(mai_mai_n284_));
  INV        m268(.A(mai_mai_n255_), .Y(mai_mai_n285_));
  OAI210     m269(.A0(mai_mai_n264_), .A1(mai_mai_n214_), .B0(mai_mai_n285_), .Y(mai_mai_n286_));
  INV        m270(.A(mai_mai_n180_), .Y(mai_mai_n287_));
  OAI210     m271(.A0(mai_mai_n287_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n288_));
  AOI210     m272(.A0(mai_mai_n288_), .A1(mai_mai_n286_), .B0(mai_mai_n231_), .Y(mai_mai_n289_));
  NO4        m273(.A(mai_mai_n289_), .B(mai_mai_n284_), .C(mai_mai_n263_), .D(mai_mai_n252_), .Y(mai_mai_n290_));
  INV        m274(.A(x1), .Y(mai_mai_n291_));
  NO3        m275(.A(mai_mai_n291_), .B(x3), .C(mai_mai_n36_), .Y(mai_mai_n292_));
  OAI210     m276(.A0(mai_mai_n292_), .A1(mai_mai_n260_), .B0(x2), .Y(mai_mai_n293_));
  OAI210     m277(.A0(mai_mai_n287_), .A1(x6), .B0(mai_mai_n44_), .Y(mai_mai_n294_));
  AOI210     m278(.A0(mai_mai_n294_), .A1(mai_mai_n293_), .B0(mai_mai_n192_), .Y(mai_mai_n295_));
  NOi21      m279(.An(mai_mai_n273_), .B(mai_mai_n17_), .Y(mai_mai_n296_));
  NA3        m280(.A(mai_mai_n296_), .B(mai_mai_n214_), .C(mai_mai_n40_), .Y(mai_mai_n297_));
  AOI210     m281(.A0(mai_mai_n36_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n298_));
  NA3        m282(.A(mai_mai_n298_), .B(mai_mai_n166_), .C(mai_mai_n32_), .Y(mai_mai_n299_));
  NA2        m283(.A(x3), .B(x2), .Y(mai_mai_n300_));
  AOI220     m284(.A0(mai_mai_n300_), .A1(mai_mai_n231_), .B0(mai_mai_n299_), .B1(mai_mai_n297_), .Y(mai_mai_n301_));
  NAi21      m285(.An(x4), .B(x0), .Y(mai_mai_n302_));
  NO3        m286(.A(mai_mai_n302_), .B(mai_mai_n44_), .C(x2), .Y(mai_mai_n303_));
  OAI210     m287(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n303_), .Y(mai_mai_n304_));
  OAI220     m288(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n305_));
  NO2        m289(.A(x9), .B(x8), .Y(mai_mai_n306_));
  NA3        m290(.A(mai_mai_n306_), .B(mai_mai_n36_), .C(mai_mai_n54_), .Y(mai_mai_n307_));
  OAI210     m291(.A0(mai_mai_n298_), .A1(mai_mai_n296_), .B0(mai_mai_n307_), .Y(mai_mai_n308_));
  AOI220     m292(.A0(mai_mai_n308_), .A1(mai_mai_n82_), .B0(mai_mai_n305_), .B1(mai_mai_n31_), .Y(mai_mai_n309_));
  AOI210     m293(.A0(mai_mai_n309_), .A1(mai_mai_n304_), .B0(mai_mai_n25_), .Y(mai_mai_n310_));
  NA3        m294(.A(mai_mai_n36_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n311_));
  OAI210     m295(.A0(mai_mai_n298_), .A1(mai_mai_n296_), .B0(mai_mai_n311_), .Y(mai_mai_n312_));
  INV        m296(.A(mai_mai_n216_), .Y(mai_mai_n313_));
  NA2        m297(.A(mai_mai_n36_), .B(mai_mai_n43_), .Y(mai_mai_n314_));
  OR2        m298(.A(mai_mai_n314_), .B(mai_mai_n281_), .Y(mai_mai_n315_));
  OAI220     m299(.A0(mai_mai_n315_), .A1(mai_mai_n165_), .B0(mai_mai_n235_), .B1(mai_mai_n313_), .Y(mai_mai_n316_));
  AO210      m300(.A0(mai_mai_n312_), .A1(mai_mai_n152_), .B0(mai_mai_n316_), .Y(mai_mai_n317_));
  NO4        m301(.A(mai_mai_n317_), .B(mai_mai_n310_), .C(mai_mai_n301_), .D(mai_mai_n295_), .Y(mai_mai_n318_));
  OAI210     m302(.A0(mai_mai_n290_), .A1(mai_mai_n247_), .B0(mai_mai_n318_), .Y(mai04));
  OAI210     m303(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n320_));
  NA3        m304(.A(mai_mai_n320_), .B(mai_mai_n271_), .C(mai_mai_n85_), .Y(mai_mai_n321_));
  NO2        m305(.A(x2), .B(x1), .Y(mai_mai_n322_));
  OAI210     m306(.A0(mai_mai_n256_), .A1(mai_mai_n322_), .B0(mai_mai_n36_), .Y(mai_mai_n323_));
  NO2        m307(.A(mai_mai_n322_), .B(mai_mai_n302_), .Y(mai_mai_n324_));
  AOI210     m308(.A0(mai_mai_n62_), .A1(x4), .B0(mai_mai_n114_), .Y(mai_mai_n325_));
  OAI210     m309(.A0(mai_mai_n325_), .A1(mai_mai_n324_), .B0(mai_mai_n248_), .Y(mai_mai_n326_));
  NO2        m310(.A(mai_mai_n270_), .B(mai_mai_n92_), .Y(mai_mai_n327_));
  NO2        m311(.A(mai_mai_n327_), .B(mai_mai_n36_), .Y(mai_mai_n328_));
  NO2        m312(.A(mai_mai_n300_), .B(mai_mai_n207_), .Y(mai_mai_n329_));
  NA2        m313(.A(mai_mai_n329_), .B(mai_mai_n94_), .Y(mai_mai_n330_));
  NA3        m314(.A(mai_mai_n330_), .B(mai_mai_n328_), .C(mai_mai_n326_), .Y(mai_mai_n331_));
  NA2        m315(.A(mai_mai_n331_), .B(mai_mai_n323_), .Y(mai_mai_n332_));
  NO3        m316(.A(mai_mai_n255_), .B(mai_mai_n122_), .C(mai_mai_n18_), .Y(mai_mai_n333_));
  INV        m317(.A(mai_mai_n333_), .Y(mai_mai_n334_));
  OAI210     m318(.A0(mai_mai_n120_), .A1(mai_mai_n108_), .B0(mai_mai_n180_), .Y(mai_mai_n335_));
  NA3        m319(.A(mai_mai_n335_), .B(x6), .C(x3), .Y(mai_mai_n336_));
  NOi21      m320(.An(mai_mai_n154_), .B(mai_mai_n134_), .Y(mai_mai_n337_));
  AOI210     m321(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n338_));
  OAI220     m322(.A0(mai_mai_n338_), .A1(mai_mai_n314_), .B0(mai_mai_n270_), .B1(mai_mai_n311_), .Y(mai_mai_n339_));
  AOI210     m323(.A0(mai_mai_n337_), .A1(mai_mai_n63_), .B0(mai_mai_n339_), .Y(mai_mai_n340_));
  NA2        m324(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n341_));
  OAI210     m325(.A0(mai_mai_n108_), .A1(mai_mai_n17_), .B0(mai_mai_n341_), .Y(mai_mai_n342_));
  NA2        m326(.A(mai_mai_n342_), .B(mai_mai_n79_), .Y(mai_mai_n343_));
  NA4        m327(.A(mai_mai_n343_), .B(mai_mai_n340_), .C(mai_mai_n336_), .D(mai_mai_n334_), .Y(mai_mai_n344_));
  OAI210     m328(.A0(mai_mai_n113_), .A1(x3), .B0(mai_mai_n303_), .Y(mai_mai_n345_));
  NA2        m329(.A(mai_mai_n345_), .B(mai_mai_n157_), .Y(mai_mai_n346_));
  AOI210     m330(.A0(mai_mai_n344_), .A1(x4), .B0(mai_mai_n346_), .Y(mai_mai_n347_));
  NA2        m331(.A(mai_mai_n324_), .B(mai_mai_n94_), .Y(mai_mai_n348_));
  NOi21      m332(.An(x4), .B(x0), .Y(mai_mai_n349_));
  XO2        m333(.A(x4), .B(x0), .Y(mai_mai_n350_));
  OAI210     m334(.A0(mai_mai_n350_), .A1(mai_mai_n119_), .B0(mai_mai_n265_), .Y(mai_mai_n351_));
  AOI220     m335(.A0(mai_mai_n351_), .A1(x8), .B0(mai_mai_n349_), .B1(mai_mai_n95_), .Y(mai_mai_n352_));
  AOI210     m336(.A0(mai_mai_n352_), .A1(mai_mai_n348_), .B0(x3), .Y(mai_mai_n353_));
  INV        m337(.A(mai_mai_n95_), .Y(mai_mai_n354_));
  NO2        m338(.A(mai_mai_n94_), .B(x4), .Y(mai_mai_n355_));
  AOI220     m339(.A0(mai_mai_n355_), .A1(mai_mai_n44_), .B0(mai_mai_n128_), .B1(mai_mai_n354_), .Y(mai_mai_n356_));
  NO2        m340(.A(mai_mai_n350_), .B(x2), .Y(mai_mai_n357_));
  NO3        m341(.A(mai_mai_n227_), .B(mai_mai_n28_), .C(mai_mai_n24_), .Y(mai_mai_n358_));
  NO2        m342(.A(mai_mai_n358_), .B(mai_mai_n357_), .Y(mai_mai_n359_));
  NA4        m343(.A(mai_mai_n359_), .B(mai_mai_n356_), .C(mai_mai_n223_), .D(x6), .Y(mai_mai_n360_));
  OAI220     m344(.A0(mai_mai_n302_), .A1(mai_mai_n92_), .B0(mai_mai_n185_), .B1(mai_mai_n94_), .Y(mai_mai_n361_));
  NO2        m345(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n362_));
  OR2        m346(.A(mai_mai_n355_), .B(mai_mai_n362_), .Y(mai_mai_n363_));
  NO2        m347(.A(mai_mai_n154_), .B(mai_mai_n108_), .Y(mai_mai_n364_));
  AOI220     m348(.A0(mai_mai_n364_), .A1(mai_mai_n363_), .B0(mai_mai_n361_), .B1(mai_mai_n61_), .Y(mai_mai_n365_));
  NO2        m349(.A(mai_mai_n154_), .B(mai_mai_n81_), .Y(mai_mai_n366_));
  NO2        m350(.A(mai_mai_n35_), .B(x2), .Y(mai_mai_n367_));
  NOi21      m351(.An(mai_mai_n125_), .B(mai_mai_n27_), .Y(mai_mai_n368_));
  AOI210     m352(.A0(mai_mai_n367_), .A1(mai_mai_n366_), .B0(mai_mai_n368_), .Y(mai_mai_n369_));
  OAI210     m353(.A0(mai_mai_n365_), .A1(mai_mai_n62_), .B0(mai_mai_n369_), .Y(mai_mai_n370_));
  OAI220     m354(.A0(mai_mai_n370_), .A1(x6), .B0(mai_mai_n360_), .B1(mai_mai_n353_), .Y(mai_mai_n371_));
  NA2        m355(.A(mai_mai_n48_), .B(mai_mai_n42_), .Y(mai_mai_n372_));
  OAI210     m356(.A0(mai_mai_n372_), .A1(mai_mai_n94_), .B0(mai_mai_n315_), .Y(mai_mai_n373_));
  AOI210     m357(.A0(mai_mai_n373_), .A1(mai_mai_n18_), .B0(mai_mai_n157_), .Y(mai_mai_n374_));
  AO220      m358(.A0(mai_mai_n374_), .A1(mai_mai_n371_), .B0(mai_mai_n347_), .B1(mai_mai_n332_), .Y(mai_mai_n375_));
  NA2        m359(.A(mai_mai_n367_), .B(x6), .Y(mai_mai_n376_));
  AOI210     m360(.A0(x6), .A1(x1), .B0(mai_mai_n156_), .Y(mai_mai_n377_));
  NA2        m361(.A(mai_mai_n355_), .B(x0), .Y(mai_mai_n378_));
  NA2        m362(.A(mai_mai_n84_), .B(x6), .Y(mai_mai_n379_));
  OAI210     m363(.A0(mai_mai_n378_), .A1(mai_mai_n377_), .B0(mai_mai_n379_), .Y(mai_mai_n380_));
  AOI220     m364(.A0(mai_mai_n380_), .A1(mai_mai_n376_), .B0(mai_mai_n217_), .B1(mai_mai_n49_), .Y(mai_mai_n381_));
  NA3        m365(.A(mai_mai_n381_), .B(mai_mai_n375_), .C(mai_mai_n321_), .Y(mai_mai_n382_));
  AOI210     m366(.A0(mai_mai_n203_), .A1(x8), .B0(mai_mai_n113_), .Y(mai_mai_n383_));
  NA2        m367(.A(mai_mai_n383_), .B(mai_mai_n341_), .Y(mai_mai_n384_));
  NA3        m368(.A(mai_mai_n384_), .B(mai_mai_n201_), .C(mai_mai_n157_), .Y(mai_mai_n385_));
  OAI210     m369(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n231_), .Y(mai_mai_n386_));
  AO220      m370(.A0(mai_mai_n386_), .A1(mai_mai_n153_), .B0(mai_mai_n112_), .B1(x4), .Y(mai_mai_n387_));
  NA3        m371(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n388_));
  NO2        m372(.A(mai_mai_n388_), .B(mai_mai_n354_), .Y(mai_mai_n389_));
  AOI210     m373(.A0(mai_mai_n387_), .A1(mai_mai_n121_), .B0(mai_mai_n389_), .Y(mai_mai_n390_));
  AOI210     m374(.A0(mai_mai_n390_), .A1(mai_mai_n385_), .B0(mai_mai_n25_), .Y(mai_mai_n391_));
  NA3        m375(.A(mai_mai_n123_), .B(mai_mai_n222_), .C(x0), .Y(mai_mai_n392_));
  AOI210     m376(.A0(mai_mai_n122_), .A1(mai_mai_n120_), .B0(mai_mai_n42_), .Y(mai_mai_n393_));
  NOi31      m377(.An(mai_mai_n393_), .B(mai_mai_n362_), .C(mai_mai_n186_), .Y(mai_mai_n394_));
  NA2        m378(.A(mai_mai_n394_), .B(mai_mai_n153_), .Y(mai_mai_n395_));
  NAi31      m379(.An(mai_mai_n50_), .B(mai_mai_n291_), .C(mai_mai_n181_), .Y(mai_mai_n396_));
  NA3        m380(.A(mai_mai_n396_), .B(mai_mai_n395_), .C(mai_mai_n392_), .Y(mai_mai_n397_));
  OAI210     m381(.A0(mai_mai_n397_), .A1(mai_mai_n391_), .B0(x6), .Y(mai_mai_n398_));
  NA2        m382(.A(mai_mai_n48_), .B(mai_mai_n139_), .Y(mai_mai_n399_));
  NA3        m383(.A(mai_mai_n55_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n400_));
  AOI220     m384(.A0(mai_mai_n400_), .A1(mai_mai_n399_), .B0(mai_mai_n40_), .B1(mai_mai_n32_), .Y(mai_mai_n401_));
  NO2        m385(.A(mai_mai_n157_), .B(x0), .Y(mai_mai_n402_));
  AOI220     m386(.A0(mai_mai_n402_), .A1(mai_mai_n222_), .B0(mai_mai_n201_), .B1(mai_mai_n157_), .Y(mai_mai_n403_));
  AOI210     m387(.A0(mai_mai_n130_), .A1(mai_mai_n253_), .B0(x1), .Y(mai_mai_n404_));
  OAI210     m388(.A0(mai_mai_n403_), .A1(x8), .B0(mai_mai_n404_), .Y(mai_mai_n405_));
  NAi31      m389(.An(x2), .B(x8), .C(x0), .Y(mai_mai_n406_));
  OAI210     m390(.A0(mai_mai_n406_), .A1(x4), .B0(mai_mai_n168_), .Y(mai_mai_n407_));
  NA3        m391(.A(mai_mai_n407_), .B(mai_mai_n151_), .C(x9), .Y(mai_mai_n408_));
  NO4        m392(.A(mai_mai_n129_), .B(mai_mai_n302_), .C(x9), .D(x2), .Y(mai_mai_n409_));
  NO2        m393(.A(mai_mai_n409_), .B(mai_mai_n18_), .Y(mai_mai_n410_));
  NO3        m394(.A(x9), .B(mai_mai_n157_), .C(x0), .Y(mai_mai_n411_));
  AOI220     m395(.A0(mai_mai_n411_), .A1(mai_mai_n248_), .B0(mai_mai_n366_), .B1(mai_mai_n157_), .Y(mai_mai_n412_));
  NA4        m396(.A(mai_mai_n412_), .B(mai_mai_n410_), .C(mai_mai_n408_), .D(mai_mai_n50_), .Y(mai_mai_n413_));
  OAI210     m397(.A0(mai_mai_n405_), .A1(mai_mai_n401_), .B0(mai_mai_n413_), .Y(mai_mai_n414_));
  NOi31      m398(.An(mai_mai_n402_), .B(mai_mai_n32_), .C(x8), .Y(mai_mai_n415_));
  AOI210     m399(.A0(mai_mai_n38_), .A1(x9), .B0(mai_mai_n137_), .Y(mai_mai_n416_));
  NO2        m400(.A(mai_mai_n416_), .B(mai_mai_n43_), .Y(mai_mai_n417_));
  NOi31      m401(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n418_));
  INV        m402(.A(mai_mai_n418_), .Y(mai_mai_n419_));
  AOI210     m403(.A0(mai_mai_n265_), .A1(mai_mai_n60_), .B0(mai_mai_n127_), .Y(mai_mai_n420_));
  OAI210     m404(.A0(mai_mai_n420_), .A1(x3), .B0(mai_mai_n419_), .Y(mai_mai_n421_));
  NO3        m405(.A(mai_mai_n421_), .B(mai_mai_n417_), .C(x2), .Y(mai_mai_n422_));
  OAI220     m406(.A0(mai_mai_n350_), .A1(mai_mai_n306_), .B0(mai_mai_n302_), .B1(mai_mai_n43_), .Y(mai_mai_n423_));
  AOI210     m407(.A0(x9), .A1(mai_mai_n48_), .B0(mai_mai_n388_), .Y(mai_mai_n424_));
  AOI220     m408(.A0(mai_mai_n424_), .A1(mai_mai_n94_), .B0(mai_mai_n423_), .B1(mai_mai_n157_), .Y(mai_mai_n425_));
  NO2        m409(.A(mai_mai_n425_), .B(mai_mai_n54_), .Y(mai_mai_n426_));
  NO3        m410(.A(mai_mai_n426_), .B(mai_mai_n422_), .C(mai_mai_n415_), .Y(mai_mai_n427_));
  AOI210     m411(.A0(mai_mai_n427_), .A1(mai_mai_n414_), .B0(mai_mai_n25_), .Y(mai_mai_n428_));
  NO3        m412(.A(mai_mai_n62_), .B(x4), .C(x1), .Y(mai_mai_n429_));
  NO3        m413(.A(mai_mai_n67_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n430_));
  AOI220     m414(.A0(mai_mai_n430_), .A1(mai_mai_n266_), .B0(mai_mai_n429_), .B1(mai_mai_n393_), .Y(mai_mai_n431_));
  NO2        m415(.A(mai_mai_n431_), .B(mai_mai_n105_), .Y(mai_mai_n432_));
  NO3        m416(.A(mai_mai_n270_), .B(mai_mai_n180_), .C(mai_mai_n40_), .Y(mai_mai_n433_));
  OAI210     m417(.A0(mai_mai_n433_), .A1(mai_mai_n432_), .B0(x7), .Y(mai_mai_n434_));
  NA2        m418(.A(mai_mai_n227_), .B(x7), .Y(mai_mai_n435_));
  NA3        m419(.A(mai_mai_n435_), .B(mai_mai_n156_), .C(mai_mai_n138_), .Y(mai_mai_n436_));
  NA2        m420(.A(mai_mai_n436_), .B(mai_mai_n434_), .Y(mai_mai_n437_));
  OAI210     m421(.A0(mai_mai_n437_), .A1(mai_mai_n428_), .B0(mai_mai_n36_), .Y(mai_mai_n438_));
  NO2        m422(.A(mai_mai_n411_), .B(mai_mai_n207_), .Y(mai_mai_n439_));
  NO4        m423(.A(mai_mai_n439_), .B(mai_mai_n78_), .C(x4), .D(mai_mai_n54_), .Y(mai_mai_n440_));
  NA2        m424(.A(mai_mai_n256_), .B(mai_mai_n21_), .Y(mai_mai_n441_));
  NO2        m425(.A(mai_mai_n165_), .B(mai_mai_n139_), .Y(mai_mai_n442_));
  NA2        m426(.A(mai_mai_n442_), .B(mai_mai_n441_), .Y(mai_mai_n443_));
  AOI210     m427(.A0(mai_mai_n443_), .A1(mai_mai_n171_), .B0(mai_mai_n28_), .Y(mai_mai_n444_));
  AOI220     m428(.A0(mai_mai_n362_), .A1(mai_mai_n94_), .B0(mai_mai_n154_), .B1(mai_mai_n203_), .Y(mai_mai_n445_));
  NA3        m429(.A(mai_mai_n445_), .B(mai_mai_n406_), .C(mai_mai_n92_), .Y(mai_mai_n446_));
  NA2        m430(.A(mai_mai_n446_), .B(mai_mai_n181_), .Y(mai_mai_n447_));
  OAI220     m431(.A0(mai_mai_n278_), .A1(mai_mai_n68_), .B0(mai_mai_n165_), .B1(mai_mai_n43_), .Y(mai_mai_n448_));
  NA2        m432(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n449_));
  AOI210     m433(.A0(mai_mai_n168_), .A1(mai_mai_n27_), .B0(mai_mai_n73_), .Y(mai_mai_n450_));
  OAI210     m434(.A0(mai_mai_n153_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n451_));
  NO3        m435(.A(mai_mai_n418_), .B(x3), .C(mai_mai_n54_), .Y(mai_mai_n452_));
  AOI210     m436(.A0(mai_mai_n452_), .A1(mai_mai_n451_), .B0(mai_mai_n450_), .Y(mai_mai_n453_));
  OAI210     m437(.A0(mai_mai_n158_), .A1(mai_mai_n449_), .B0(mai_mai_n453_), .Y(mai_mai_n454_));
  AOI220     m438(.A0(mai_mai_n454_), .A1(x0), .B0(mai_mai_n448_), .B1(mai_mai_n139_), .Y(mai_mai_n455_));
  AOI210     m439(.A0(mai_mai_n455_), .A1(mai_mai_n447_), .B0(mai_mai_n235_), .Y(mai_mai_n456_));
  NA2        m440(.A(x9), .B(x5), .Y(mai_mai_n457_));
  NO4        m441(.A(mai_mai_n108_), .B(mai_mai_n457_), .C(mai_mai_n60_), .D(mai_mai_n32_), .Y(mai_mai_n458_));
  NO4        m442(.A(mai_mai_n458_), .B(mai_mai_n456_), .C(mai_mai_n444_), .D(mai_mai_n440_), .Y(mai_mai_n459_));
  NA3        m443(.A(mai_mai_n459_), .B(mai_mai_n438_), .C(mai_mai_n398_), .Y(mai_mai_n460_));
  AOI210     m444(.A0(mai_mai_n382_), .A1(mai_mai_n25_), .B0(mai_mai_n460_), .Y(mai05));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  INV        u012(.A(men_men_n24_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  OA210      u015(.A0(men_men_n31_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n32_));
  NOi31      u016(.An(men_men_n23_), .B(men_men_n32_), .C(men_men_n29_), .Y(men00));
  NO2        u017(.A(x1), .B(x0), .Y(men_men_n34_));
  INV        u018(.A(x6), .Y(men_men_n35_));
  NO2        u019(.A(men_men_n35_), .B(men_men_n25_), .Y(men_men_n36_));
  AN2        u020(.A(x8), .B(x7), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  NO2        u022(.A(men_men_n23_), .B(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n36_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n50_));
  AOI220     u034(.A0(men_men_n50_), .A1(men_men_n34_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n51_));
  INV        u035(.A(x2), .Y(men_men_n52_));
  NO2        u036(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  OAI210     u039(.A0(men_men_n51_), .A1(men_men_n31_), .B0(men_men_n55_), .Y(men_men_n56_));
  NO3        u040(.A(men_men_n56_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u041(.A(x8), .B(x7), .Y(men_men_n58_));
  NA2        u042(.A(men_men_n41_), .B(x1), .Y(men_men_n59_));
  INV        u043(.A(x9), .Y(men_men_n60_));
  NO2        u044(.A(men_men_n60_), .B(men_men_n35_), .Y(men_men_n61_));
  INV        u045(.A(men_men_n61_), .Y(men_men_n62_));
  NO3        u046(.A(men_men_n62_), .B(men_men_n59_), .C(men_men_n58_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n59_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  NO2        u051(.A(men_men_n67_), .B(x1), .Y(men_men_n68_));
  OA210      u052(.A0(men_men_n68_), .A1(men_men_n65_), .B0(men_men_n64_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n42_), .A1(men_men_n25_), .B0(men_men_n52_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n54_), .A1(men_men_n20_), .B0(men_men_n70_), .Y(men_men_n71_));
  NAi31      u055(.An(x1), .B(x9), .C(x5), .Y(men_men_n72_));
  OAI220     u056(.A0(men_men_n72_), .A1(men_men_n41_), .B0(men_men_n71_), .B1(men_men_n69_), .Y(men_men_n73_));
  OAI210     u057(.A0(men_men_n73_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n74_));
  NA2        u058(.A(men_men_n46_), .B(x2), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n76_));
  NA2        u060(.A(x5), .B(x3), .Y(men_men_n77_));
  NO2        u061(.A(x8), .B(x6), .Y(men_men_n78_));
  NO4        u062(.A(men_men_n78_), .B(men_men_n77_), .C(men_men_n64_), .D(men_men_n52_), .Y(men_men_n79_));
  NAi21      u063(.An(x4), .B(x3), .Y(men_men_n80_));
  INV        u064(.A(men_men_n80_), .Y(men_men_n81_));
  NO2        u065(.A(men_men_n81_), .B(men_men_n22_), .Y(men_men_n82_));
  NO2        u066(.A(x4), .B(x2), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n83_), .B(x3), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n82_), .C(men_men_n18_), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n85_), .B(men_men_n79_), .C(men_men_n76_), .Y(men_men_n86_));
  NO4        u070(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .D(x1), .Y(men_men_n87_));
  NA2        u071(.A(men_men_n60_), .B(men_men_n46_), .Y(men_men_n88_));
  INV        u072(.A(men_men_n88_), .Y(men_men_n89_));
  OAI210     u073(.A0(men_men_n87_), .A1(men_men_n65_), .B0(men_men_n89_), .Y(men_men_n90_));
  NA2        u074(.A(x3), .B(men_men_n18_), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n25_), .Y(men_men_n92_));
  INV        u076(.A(x8), .Y(men_men_n93_));
  NA2        u077(.A(x2), .B(x1), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n92_), .Y(men_men_n96_));
  NO2        u080(.A(men_men_n96_), .B(men_men_n26_), .Y(men_men_n97_));
  AOI210     u081(.A0(men_men_n54_), .A1(men_men_n25_), .B0(men_men_n52_), .Y(men_men_n98_));
  OAI210     u082(.A0(men_men_n43_), .A1(men_men_n36_), .B0(men_men_n46_), .Y(men_men_n99_));
  NO3        u083(.A(men_men_n99_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n100_));
  NA2        u084(.A(x4), .B(men_men_n41_), .Y(men_men_n101_));
  NO2        u085(.A(men_men_n46_), .B(men_men_n52_), .Y(men_men_n102_));
  NA2        u086(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n103_));
  AOI210     u087(.A0(men_men_n101_), .A1(men_men_n50_), .B0(men_men_n103_), .Y(men_men_n104_));
  NO2        u088(.A(x3), .B(x2), .Y(men_men_n105_));
  NA3        u089(.A(men_men_n105_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n106_));
  INV        u090(.A(men_men_n106_), .Y(men_men_n107_));
  NA2        u091(.A(men_men_n52_), .B(x1), .Y(men_men_n108_));
  OAI210     u092(.A0(men_men_n108_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n109_));
  NO4        u093(.A(men_men_n109_), .B(men_men_n107_), .C(men_men_n104_), .D(men_men_n100_), .Y(men_men_n110_));
  AO220      u094(.A0(men_men_n110_), .A1(men_men_n90_), .B0(men_men_n86_), .B1(men_men_n74_), .Y(men02));
  NO2        u095(.A(x3), .B(men_men_n52_), .Y(men_men_n112_));
  NO2        u096(.A(x8), .B(men_men_n18_), .Y(men_men_n113_));
  NA2        u097(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n114_));
  NA2        u098(.A(men_men_n41_), .B(x0), .Y(men_men_n115_));
  OAI210     u099(.A0(men_men_n88_), .A1(men_men_n114_), .B0(men_men_n115_), .Y(men_men_n116_));
  AOI220     u100(.A0(men_men_n116_), .A1(men_men_n113_), .B0(men_men_n112_), .B1(x4), .Y(men_men_n117_));
  NO3        u101(.A(men_men_n117_), .B(x7), .C(x5), .Y(men_men_n118_));
  NA2        u102(.A(x9), .B(x2), .Y(men_men_n119_));
  OR2        u103(.A(x8), .B(x0), .Y(men_men_n120_));
  INV        u104(.A(men_men_n120_), .Y(men_men_n121_));
  NAi21      u105(.An(x2), .B(x8), .Y(men_men_n122_));
  INV        u106(.A(men_men_n122_), .Y(men_men_n123_));
  NO2        u107(.A(men_men_n123_), .B(men_men_n121_), .Y(men_men_n124_));
  NO2        u108(.A(x4), .B(x1), .Y(men_men_n125_));
  NA3        u109(.A(men_men_n125_), .B(men_men_n124_), .C(men_men_n58_), .Y(men_men_n126_));
  NOi21      u110(.An(x0), .B(x1), .Y(men_men_n127_));
  NO3        u111(.A(x9), .B(x8), .C(x7), .Y(men_men_n128_));
  NOi21      u112(.An(x0), .B(x4), .Y(men_men_n129_));
  NA2        u113(.A(men_men_n128_), .B(men_men_n127_), .Y(men_men_n130_));
  AOI210     u114(.A0(men_men_n130_), .A1(men_men_n126_), .B0(men_men_n77_), .Y(men_men_n131_));
  NO2        u115(.A(x5), .B(men_men_n46_), .Y(men_men_n132_));
  NA2        u116(.A(x2), .B(men_men_n18_), .Y(men_men_n133_));
  AOI210     u117(.A0(men_men_n133_), .A1(men_men_n108_), .B0(men_men_n115_), .Y(men_men_n134_));
  OAI210     u118(.A0(men_men_n134_), .A1(men_men_n34_), .B0(men_men_n132_), .Y(men_men_n135_));
  NAi21      u119(.An(x0), .B(x4), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n136_), .B(x1), .Y(men_men_n137_));
  NO2        u121(.A(x7), .B(x0), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n83_), .B(men_men_n102_), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n139_), .B(x3), .Y(men_men_n140_));
  OAI210     u124(.A0(men_men_n138_), .A1(men_men_n137_), .B0(men_men_n140_), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n21_), .B(men_men_n41_), .Y(men_men_n142_));
  NA2        u126(.A(x5), .B(x0), .Y(men_men_n143_));
  NO2        u127(.A(men_men_n46_), .B(x2), .Y(men_men_n144_));
  NA3        u128(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n142_), .Y(men_men_n145_));
  NA4        u129(.A(men_men_n145_), .B(men_men_n141_), .C(men_men_n135_), .D(men_men_n35_), .Y(men_men_n146_));
  NO3        u130(.A(men_men_n146_), .B(men_men_n131_), .C(men_men_n118_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n77_), .B(men_men_n75_), .C(men_men_n24_), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n149_));
  AOI220     u133(.A0(men_men_n127_), .A1(men_men_n149_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n150_));
  NO3        u134(.A(men_men_n150_), .B(men_men_n58_), .C(men_men_n60_), .Y(men_men_n151_));
  NA2        u135(.A(x7), .B(x3), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n101_), .B(x5), .Y(men_men_n153_));
  NO2        u137(.A(x9), .B(x7), .Y(men_men_n154_));
  NOi21      u138(.An(x8), .B(x0), .Y(men_men_n155_));
  NO2        u139(.A(men_men_n41_), .B(x2), .Y(men_men_n156_));
  INV        u140(.A(x7), .Y(men_men_n157_));
  NA2        u141(.A(men_men_n157_), .B(men_men_n18_), .Y(men_men_n158_));
  AOI220     u142(.A0(men_men_n158_), .A1(men_men_n156_), .B0(men_men_n112_), .B1(men_men_n37_), .Y(men_men_n159_));
  NO2        u143(.A(men_men_n25_), .B(x4), .Y(men_men_n160_));
  NO2        u144(.A(men_men_n160_), .B(men_men_n129_), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n161_), .B(men_men_n159_), .Y(men_men_n162_));
  INV        u146(.A(men_men_n162_), .Y(men_men_n163_));
  OAI210     u147(.A0(men_men_n152_), .A1(men_men_n48_), .B0(men_men_n163_), .Y(men_men_n164_));
  NA2        u148(.A(x5), .B(x1), .Y(men_men_n165_));
  INV        u149(.A(men_men_n165_), .Y(men_men_n166_));
  AOI210     u150(.A0(men_men_n166_), .A1(men_men_n129_), .B0(men_men_n35_), .Y(men_men_n167_));
  NO2        u151(.A(men_men_n60_), .B(men_men_n93_), .Y(men_men_n168_));
  NAi21      u152(.An(x2), .B(x7), .Y(men_men_n169_));
  NO3        u153(.A(men_men_n169_), .B(men_men_n168_), .C(men_men_n46_), .Y(men_men_n170_));
  NA2        u154(.A(men_men_n170_), .B(men_men_n65_), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n171_), .B(men_men_n167_), .Y(men_men_n172_));
  NO4        u156(.A(men_men_n172_), .B(men_men_n164_), .C(men_men_n151_), .D(men_men_n148_), .Y(men_men_n173_));
  NO2        u157(.A(men_men_n173_), .B(men_men_n147_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n143_), .B(men_men_n139_), .Y(men_men_n175_));
  NA2        u159(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n176_));
  NA2        u160(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n177_));
  NA3        u161(.A(men_men_n177_), .B(men_men_n176_), .C(men_men_n24_), .Y(men_men_n178_));
  AN2        u162(.A(men_men_n178_), .B(men_men_n144_), .Y(men_men_n179_));
  NA2        u163(.A(x8), .B(x0), .Y(men_men_n180_));
  NO2        u164(.A(men_men_n157_), .B(men_men_n25_), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n127_), .B(x4), .Y(men_men_n182_));
  NA2        u166(.A(men_men_n182_), .B(men_men_n181_), .Y(men_men_n183_));
  AOI210     u167(.A0(men_men_n180_), .A1(men_men_n133_), .B0(men_men_n183_), .Y(men_men_n184_));
  NA2        u168(.A(x2), .B(x0), .Y(men_men_n185_));
  NA2        u169(.A(x4), .B(x1), .Y(men_men_n186_));
  NAi21      u170(.An(men_men_n125_), .B(men_men_n186_), .Y(men_men_n187_));
  NOi31      u171(.An(men_men_n187_), .B(men_men_n160_), .C(men_men_n185_), .Y(men_men_n188_));
  NO4        u172(.A(men_men_n188_), .B(men_men_n184_), .C(men_men_n179_), .D(men_men_n175_), .Y(men_men_n189_));
  NO2        u173(.A(men_men_n189_), .B(men_men_n41_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n178_), .B(men_men_n75_), .Y(men_men_n191_));
  INV        u175(.A(men_men_n132_), .Y(men_men_n192_));
  NO2        u176(.A(men_men_n108_), .B(men_men_n17_), .Y(men_men_n193_));
  AOI210     u177(.A0(men_men_n34_), .A1(men_men_n93_), .B0(men_men_n193_), .Y(men_men_n194_));
  NO3        u178(.A(men_men_n194_), .B(men_men_n192_), .C(x7), .Y(men_men_n195_));
  NA3        u179(.A(men_men_n187_), .B(men_men_n192_), .C(men_men_n40_), .Y(men_men_n196_));
  OAI210     u180(.A0(men_men_n177_), .A1(men_men_n139_), .B0(men_men_n196_), .Y(men_men_n197_));
  NO3        u181(.A(men_men_n197_), .B(men_men_n195_), .C(men_men_n191_), .Y(men_men_n198_));
  NO2        u182(.A(men_men_n198_), .B(x3), .Y(men_men_n199_));
  NO3        u183(.A(men_men_n199_), .B(men_men_n190_), .C(men_men_n174_), .Y(men03));
  NO2        u184(.A(men_men_n46_), .B(x3), .Y(men_men_n201_));
  NO2        u185(.A(x6), .B(men_men_n25_), .Y(men_men_n202_));
  INV        u186(.A(men_men_n202_), .Y(men_men_n203_));
  NO2        u187(.A(men_men_n52_), .B(x1), .Y(men_men_n204_));
  OAI210     u188(.A0(men_men_n204_), .A1(men_men_n25_), .B0(men_men_n61_), .Y(men_men_n205_));
  OAI220     u189(.A0(men_men_n205_), .A1(men_men_n17_), .B0(men_men_n203_), .B1(men_men_n108_), .Y(men_men_n206_));
  NA2        u190(.A(men_men_n206_), .B(men_men_n201_), .Y(men_men_n207_));
  NO2        u191(.A(men_men_n77_), .B(x6), .Y(men_men_n208_));
  NA2        u192(.A(x6), .B(men_men_n25_), .Y(men_men_n209_));
  NO2        u193(.A(men_men_n209_), .B(x4), .Y(men_men_n210_));
  NO2        u194(.A(men_men_n18_), .B(x0), .Y(men_men_n211_));
  AO220      u195(.A0(men_men_n211_), .A1(men_men_n210_), .B0(men_men_n208_), .B1(men_men_n53_), .Y(men_men_n212_));
  NA2        u196(.A(men_men_n212_), .B(men_men_n60_), .Y(men_men_n213_));
  NA2        u197(.A(x3), .B(men_men_n17_), .Y(men_men_n214_));
  NO2        u198(.A(men_men_n214_), .B(men_men_n209_), .Y(men_men_n215_));
  NA2        u199(.A(x9), .B(men_men_n52_), .Y(men_men_n216_));
  NA2        u200(.A(men_men_n216_), .B(x4), .Y(men_men_n217_));
  NA2        u201(.A(men_men_n209_), .B(men_men_n80_), .Y(men_men_n218_));
  AOI210     u202(.A0(men_men_n25_), .A1(x3), .B0(men_men_n185_), .Y(men_men_n219_));
  AOI220     u203(.A0(men_men_n219_), .A1(men_men_n218_), .B0(men_men_n217_), .B1(men_men_n215_), .Y(men_men_n220_));
  NO3        u204(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n221_));
  NO2        u205(.A(x5), .B(x1), .Y(men_men_n222_));
  AOI220     u206(.A0(men_men_n222_), .A1(men_men_n17_), .B0(men_men_n105_), .B1(x5), .Y(men_men_n223_));
  NO2        u207(.A(men_men_n214_), .B(men_men_n176_), .Y(men_men_n224_));
  NO3        u208(.A(x3), .B(x2), .C(x1), .Y(men_men_n225_));
  NO2        u209(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  OAI210     u210(.A0(men_men_n223_), .A1(men_men_n62_), .B0(men_men_n226_), .Y(men_men_n227_));
  AOI220     u211(.A0(men_men_n227_), .A1(men_men_n46_), .B0(men_men_n221_), .B1(men_men_n132_), .Y(men_men_n228_));
  NA4        u212(.A(men_men_n228_), .B(men_men_n220_), .C(men_men_n213_), .D(men_men_n207_), .Y(men_men_n229_));
  NO2        u213(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n230_));
  NA2        u214(.A(men_men_n230_), .B(men_men_n19_), .Y(men_men_n231_));
  NO2        u215(.A(x3), .B(men_men_n17_), .Y(men_men_n232_));
  NO2        u216(.A(men_men_n232_), .B(x6), .Y(men_men_n233_));
  NOi21      u217(.An(men_men_n83_), .B(men_men_n233_), .Y(men_men_n234_));
  NA2        u218(.A(men_men_n60_), .B(men_men_n93_), .Y(men_men_n235_));
  NA3        u219(.A(men_men_n235_), .B(men_men_n232_), .C(x6), .Y(men_men_n236_));
  AOI210     u220(.A0(men_men_n236_), .A1(men_men_n234_), .B0(men_men_n157_), .Y(men_men_n237_));
  AO210      u221(.A0(men_men_n237_), .A1(men_men_n231_), .B0(men_men_n181_), .Y(men_men_n238_));
  NA2        u222(.A(men_men_n41_), .B(men_men_n52_), .Y(men_men_n239_));
  NA2        u223(.A(men_men_n144_), .B(men_men_n92_), .Y(men_men_n240_));
  NA2        u224(.A(x6), .B(men_men_n46_), .Y(men_men_n241_));
  OAI210     u225(.A0(men_men_n121_), .A1(men_men_n78_), .B0(x4), .Y(men_men_n242_));
  AOI210     u226(.A0(men_men_n242_), .A1(men_men_n241_), .B0(men_men_n77_), .Y(men_men_n243_));
  NA2        u227(.A(men_men_n202_), .B(men_men_n137_), .Y(men_men_n244_));
  NA3        u228(.A(men_men_n214_), .B(men_men_n132_), .C(x6), .Y(men_men_n245_));
  OAI210     u229(.A0(men_men_n93_), .A1(men_men_n35_), .B0(men_men_n65_), .Y(men_men_n246_));
  NA3        u230(.A(men_men_n246_), .B(men_men_n245_), .C(men_men_n244_), .Y(men_men_n247_));
  OAI210     u231(.A0(men_men_n247_), .A1(men_men_n243_), .B0(x2), .Y(men_men_n248_));
  NA3        u232(.A(men_men_n248_), .B(men_men_n240_), .C(men_men_n238_), .Y(men_men_n249_));
  AOI210     u233(.A0(men_men_n229_), .A1(x8), .B0(men_men_n249_), .Y(men_men_n250_));
  NO2        u234(.A(men_men_n93_), .B(x3), .Y(men_men_n251_));
  NA2        u235(.A(men_men_n251_), .B(men_men_n210_), .Y(men_men_n252_));
  NO3        u236(.A(men_men_n91_), .B(men_men_n78_), .C(men_men_n25_), .Y(men_men_n253_));
  AOI210     u237(.A0(men_men_n233_), .A1(men_men_n160_), .B0(men_men_n253_), .Y(men_men_n254_));
  AOI210     u238(.A0(men_men_n254_), .A1(men_men_n252_), .B0(x2), .Y(men_men_n255_));
  NO2        u239(.A(x4), .B(men_men_n52_), .Y(men_men_n256_));
  AOI220     u240(.A0(men_men_n210_), .A1(men_men_n193_), .B0(men_men_n256_), .B1(men_men_n65_), .Y(men_men_n257_));
  NA2        u241(.A(men_men_n60_), .B(x6), .Y(men_men_n258_));
  NA3        u242(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n259_));
  AOI210     u243(.A0(men_men_n259_), .A1(men_men_n143_), .B0(men_men_n258_), .Y(men_men_n260_));
  NA2        u244(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n261_));
  NO2        u245(.A(men_men_n261_), .B(men_men_n25_), .Y(men_men_n262_));
  OAI210     u246(.A0(men_men_n262_), .A1(men_men_n260_), .B0(men_men_n125_), .Y(men_men_n263_));
  NA2        u247(.A(men_men_n214_), .B(x6), .Y(men_men_n264_));
  NO2        u248(.A(men_men_n214_), .B(x6), .Y(men_men_n265_));
  NAi21      u249(.An(men_men_n168_), .B(men_men_n265_), .Y(men_men_n266_));
  NA3        u250(.A(men_men_n266_), .B(men_men_n264_), .C(men_men_n149_), .Y(men_men_n267_));
  NA4        u251(.A(men_men_n267_), .B(men_men_n263_), .C(men_men_n257_), .D(men_men_n157_), .Y(men_men_n268_));
  NA2        u252(.A(men_men_n202_), .B(men_men_n232_), .Y(men_men_n269_));
  NO2        u253(.A(x9), .B(x6), .Y(men_men_n270_));
  NO2        u254(.A(men_men_n143_), .B(men_men_n18_), .Y(men_men_n271_));
  NAi21      u255(.An(men_men_n271_), .B(men_men_n259_), .Y(men_men_n272_));
  NAi21      u256(.An(x1), .B(x4), .Y(men_men_n273_));
  AOI210     u257(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n274_));
  OAI210     u258(.A0(men_men_n143_), .A1(x3), .B0(men_men_n274_), .Y(men_men_n275_));
  AOI220     u259(.A0(men_men_n275_), .A1(men_men_n273_), .B0(men_men_n272_), .B1(men_men_n270_), .Y(men_men_n276_));
  NA2        u260(.A(men_men_n276_), .B(men_men_n269_), .Y(men_men_n277_));
  NA2        u261(.A(men_men_n60_), .B(x2), .Y(men_men_n278_));
  NO2        u262(.A(men_men_n278_), .B(men_men_n269_), .Y(men_men_n279_));
  NO3        u263(.A(x9), .B(x6), .C(x0), .Y(men_men_n280_));
  NA2        u264(.A(men_men_n108_), .B(men_men_n25_), .Y(men_men_n281_));
  NA2        u265(.A(x6), .B(x2), .Y(men_men_n282_));
  NO2        u266(.A(men_men_n282_), .B(men_men_n176_), .Y(men_men_n283_));
  AOI210     u267(.A0(men_men_n281_), .A1(men_men_n280_), .B0(men_men_n283_), .Y(men_men_n284_));
  OAI220     u268(.A0(men_men_n284_), .A1(men_men_n41_), .B0(men_men_n182_), .B1(men_men_n44_), .Y(men_men_n285_));
  OAI210     u269(.A0(men_men_n285_), .A1(men_men_n279_), .B0(men_men_n277_), .Y(men_men_n286_));
  NA2        u270(.A(x9), .B(men_men_n41_), .Y(men_men_n287_));
  NO2        u271(.A(men_men_n287_), .B(men_men_n209_), .Y(men_men_n288_));
  OR3        u272(.A(men_men_n288_), .B(men_men_n208_), .C(men_men_n153_), .Y(men_men_n289_));
  NA2        u273(.A(x4), .B(x0), .Y(men_men_n290_));
  NO3        u274(.A(men_men_n72_), .B(men_men_n290_), .C(x6), .Y(men_men_n291_));
  AOI210     u275(.A0(men_men_n289_), .A1(men_men_n40_), .B0(men_men_n291_), .Y(men_men_n292_));
  AOI210     u276(.A0(men_men_n292_), .A1(men_men_n286_), .B0(x8), .Y(men_men_n293_));
  INV        u277(.A(men_men_n180_), .Y(men_men_n294_));
  OAI210     u278(.A0(men_men_n294_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n295_));
  NO2        u279(.A(men_men_n295_), .B(men_men_n239_), .Y(men_men_n296_));
  NO4        u280(.A(men_men_n296_), .B(men_men_n293_), .C(men_men_n268_), .D(men_men_n255_), .Y(men_men_n297_));
  NO2        u281(.A(men_men_n168_), .B(x1), .Y(men_men_n298_));
  NO3        u282(.A(men_men_n298_), .B(x3), .C(men_men_n35_), .Y(men_men_n299_));
  OAI210     u283(.A0(men_men_n299_), .A1(men_men_n265_), .B0(x2), .Y(men_men_n300_));
  OAI210     u284(.A0(men_men_n294_), .A1(x6), .B0(men_men_n42_), .Y(men_men_n301_));
  AOI210     u285(.A0(men_men_n301_), .A1(men_men_n300_), .B0(men_men_n192_), .Y(men_men_n302_));
  NOi21      u286(.An(men_men_n282_), .B(men_men_n17_), .Y(men_men_n303_));
  NA3        u287(.A(men_men_n303_), .B(men_men_n222_), .C(men_men_n38_), .Y(men_men_n304_));
  AOI210     u288(.A0(men_men_n35_), .A1(men_men_n52_), .B0(x0), .Y(men_men_n305_));
  NA3        u289(.A(men_men_n305_), .B(men_men_n166_), .C(men_men_n31_), .Y(men_men_n306_));
  NA2        u290(.A(x3), .B(x2), .Y(men_men_n307_));
  AOI220     u291(.A0(men_men_n307_), .A1(men_men_n239_), .B0(men_men_n306_), .B1(men_men_n304_), .Y(men_men_n308_));
  NAi21      u292(.An(x4), .B(x0), .Y(men_men_n309_));
  NO3        u293(.A(men_men_n309_), .B(men_men_n42_), .C(x2), .Y(men_men_n310_));
  OAI210     u294(.A0(x6), .A1(men_men_n18_), .B0(men_men_n310_), .Y(men_men_n311_));
  OAI220     u295(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n312_));
  NO2        u296(.A(x9), .B(x8), .Y(men_men_n313_));
  NO2        u297(.A(men_men_n305_), .B(men_men_n303_), .Y(men_men_n314_));
  AOI220     u298(.A0(men_men_n314_), .A1(men_men_n81_), .B0(men_men_n312_), .B1(men_men_n30_), .Y(men_men_n315_));
  AOI210     u299(.A0(men_men_n315_), .A1(men_men_n311_), .B0(men_men_n25_), .Y(men_men_n316_));
  NA3        u300(.A(men_men_n35_), .B(x1), .C(men_men_n17_), .Y(men_men_n317_));
  OAI210     u301(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n317_), .Y(men_men_n318_));
  INV        u302(.A(men_men_n224_), .Y(men_men_n319_));
  NA2        u303(.A(men_men_n35_), .B(men_men_n41_), .Y(men_men_n320_));
  OR2        u304(.A(men_men_n320_), .B(men_men_n290_), .Y(men_men_n321_));
  OAI220     u305(.A0(men_men_n321_), .A1(men_men_n165_), .B0(men_men_n241_), .B1(men_men_n319_), .Y(men_men_n322_));
  AO210      u306(.A0(men_men_n318_), .A1(men_men_n153_), .B0(men_men_n322_), .Y(men_men_n323_));
  NO4        u307(.A(men_men_n323_), .B(men_men_n316_), .C(men_men_n308_), .D(men_men_n302_), .Y(men_men_n324_));
  OAI210     u308(.A0(men_men_n297_), .A1(men_men_n250_), .B0(men_men_n324_), .Y(men04));
  OAI210     u309(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n326_));
  NA3        u310(.A(men_men_n326_), .B(men_men_n280_), .C(men_men_n84_), .Y(men_men_n327_));
  NO2        u311(.A(x2), .B(x1), .Y(men_men_n328_));
  OAI210     u312(.A0(men_men_n261_), .A1(men_men_n328_), .B0(men_men_n35_), .Y(men_men_n329_));
  NO2        u313(.A(men_men_n328_), .B(men_men_n309_), .Y(men_men_n330_));
  AOI210     u314(.A0(men_men_n60_), .A1(x4), .B0(men_men_n114_), .Y(men_men_n331_));
  OAI210     u315(.A0(men_men_n331_), .A1(men_men_n330_), .B0(men_men_n251_), .Y(men_men_n332_));
  NO2        u316(.A(men_men_n278_), .B(men_men_n91_), .Y(men_men_n333_));
  NO2        u317(.A(men_men_n333_), .B(men_men_n35_), .Y(men_men_n334_));
  NO2        u318(.A(men_men_n307_), .B(men_men_n211_), .Y(men_men_n335_));
  NA2        u319(.A(x9), .B(x0), .Y(men_men_n336_));
  AOI210     u320(.A0(men_men_n91_), .A1(men_men_n75_), .B0(men_men_n336_), .Y(men_men_n337_));
  OAI210     u321(.A0(men_men_n337_), .A1(men_men_n335_), .B0(men_men_n93_), .Y(men_men_n338_));
  NA3        u322(.A(men_men_n338_), .B(men_men_n334_), .C(men_men_n332_), .Y(men_men_n339_));
  NA2        u323(.A(men_men_n339_), .B(men_men_n329_), .Y(men_men_n340_));
  NO2        u324(.A(men_men_n216_), .B(men_men_n115_), .Y(men_men_n341_));
  NO3        u325(.A(men_men_n258_), .B(men_men_n122_), .C(men_men_n18_), .Y(men_men_n342_));
  NO2        u326(.A(men_men_n342_), .B(men_men_n341_), .Y(men_men_n343_));
  OAI210     u327(.A0(men_men_n120_), .A1(men_men_n108_), .B0(men_men_n180_), .Y(men_men_n344_));
  NA3        u328(.A(men_men_n344_), .B(x6), .C(x3), .Y(men_men_n345_));
  NOi21      u329(.An(men_men_n155_), .B(men_men_n133_), .Y(men_men_n346_));
  AOI210     u330(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n347_));
  OAI220     u331(.A0(men_men_n347_), .A1(men_men_n320_), .B0(men_men_n278_), .B1(men_men_n317_), .Y(men_men_n348_));
  AOI210     u332(.A0(men_men_n346_), .A1(men_men_n61_), .B0(men_men_n348_), .Y(men_men_n349_));
  NA2        u333(.A(x2), .B(men_men_n17_), .Y(men_men_n350_));
  OAI210     u334(.A0(men_men_n108_), .A1(men_men_n17_), .B0(men_men_n350_), .Y(men_men_n351_));
  AOI220     u335(.A0(men_men_n351_), .A1(men_men_n78_), .B0(men_men_n333_), .B1(men_men_n93_), .Y(men_men_n352_));
  NA4        u336(.A(men_men_n352_), .B(men_men_n349_), .C(men_men_n345_), .D(men_men_n343_), .Y(men_men_n353_));
  OAI210     u337(.A0(men_men_n113_), .A1(x3), .B0(men_men_n310_), .Y(men_men_n354_));
  NA3        u338(.A(men_men_n235_), .B(men_men_n221_), .C(men_men_n83_), .Y(men_men_n355_));
  NA3        u339(.A(men_men_n355_), .B(men_men_n354_), .C(men_men_n157_), .Y(men_men_n356_));
  AOI210     u340(.A0(men_men_n353_), .A1(x4), .B0(men_men_n356_), .Y(men_men_n357_));
  NA3        u341(.A(men_men_n330_), .B(men_men_n216_), .C(men_men_n93_), .Y(men_men_n358_));
  NOi21      u342(.An(x4), .B(x0), .Y(men_men_n359_));
  XO2        u343(.A(x4), .B(x0), .Y(men_men_n360_));
  OAI210     u344(.A0(men_men_n360_), .A1(men_men_n119_), .B0(men_men_n273_), .Y(men_men_n361_));
  AOI220     u345(.A0(men_men_n361_), .A1(x8), .B0(men_men_n359_), .B1(men_men_n94_), .Y(men_men_n362_));
  AOI210     u346(.A0(men_men_n362_), .A1(men_men_n358_), .B0(x3), .Y(men_men_n363_));
  INV        u347(.A(men_men_n94_), .Y(men_men_n364_));
  NO2        u348(.A(men_men_n93_), .B(x4), .Y(men_men_n365_));
  AOI220     u349(.A0(men_men_n365_), .A1(men_men_n42_), .B0(men_men_n129_), .B1(men_men_n364_), .Y(men_men_n366_));
  NO3        u350(.A(men_men_n360_), .B(men_men_n168_), .C(x2), .Y(men_men_n367_));
  INV        u351(.A(men_men_n367_), .Y(men_men_n368_));
  NA4        u352(.A(men_men_n368_), .B(men_men_n366_), .C(men_men_n231_), .D(x6), .Y(men_men_n369_));
  OAI220     u353(.A0(men_men_n309_), .A1(men_men_n91_), .B0(men_men_n185_), .B1(men_men_n93_), .Y(men_men_n370_));
  NO2        u354(.A(men_men_n41_), .B(x0), .Y(men_men_n371_));
  NA2        u355(.A(men_men_n370_), .B(men_men_n59_), .Y(men_men_n372_));
  NO2        u356(.A(men_men_n155_), .B(men_men_n80_), .Y(men_men_n373_));
  NO2        u357(.A(men_men_n34_), .B(x2), .Y(men_men_n374_));
  NOi21      u358(.An(men_men_n125_), .B(men_men_n27_), .Y(men_men_n375_));
  AOI210     u359(.A0(men_men_n374_), .A1(men_men_n373_), .B0(men_men_n375_), .Y(men_men_n376_));
  OAI210     u360(.A0(men_men_n372_), .A1(men_men_n60_), .B0(men_men_n376_), .Y(men_men_n377_));
  OAI220     u361(.A0(men_men_n377_), .A1(x6), .B0(men_men_n369_), .B1(men_men_n363_), .Y(men_men_n378_));
  OAI210     u362(.A0(men_men_n61_), .A1(men_men_n46_), .B0(men_men_n40_), .Y(men_men_n379_));
  OAI210     u363(.A0(men_men_n379_), .A1(men_men_n93_), .B0(men_men_n321_), .Y(men_men_n380_));
  AOI210     u364(.A0(men_men_n380_), .A1(men_men_n18_), .B0(men_men_n157_), .Y(men_men_n381_));
  AO220      u365(.A0(men_men_n381_), .A1(men_men_n378_), .B0(men_men_n357_), .B1(men_men_n340_), .Y(men_men_n382_));
  NA2        u366(.A(men_men_n374_), .B(x6), .Y(men_men_n383_));
  AOI210     u367(.A0(x6), .A1(x1), .B0(men_men_n156_), .Y(men_men_n384_));
  NA2        u368(.A(men_men_n365_), .B(x0), .Y(men_men_n385_));
  NA2        u369(.A(men_men_n83_), .B(x6), .Y(men_men_n386_));
  OAI210     u370(.A0(men_men_n385_), .A1(men_men_n384_), .B0(men_men_n386_), .Y(men_men_n387_));
  AOI220     u371(.A0(men_men_n387_), .A1(men_men_n383_), .B0(men_men_n225_), .B1(men_men_n47_), .Y(men_men_n388_));
  NA3        u372(.A(men_men_n388_), .B(men_men_n382_), .C(men_men_n327_), .Y(men_men_n389_));
  AOI210     u373(.A0(men_men_n204_), .A1(x8), .B0(men_men_n113_), .Y(men_men_n390_));
  NA2        u374(.A(men_men_n390_), .B(men_men_n350_), .Y(men_men_n391_));
  NA3        u375(.A(men_men_n391_), .B(men_men_n201_), .C(men_men_n157_), .Y(men_men_n392_));
  OAI210     u376(.A0(men_men_n28_), .A1(x1), .B0(men_men_n239_), .Y(men_men_n393_));
  AO220      u377(.A0(men_men_n393_), .A1(men_men_n154_), .B0(men_men_n112_), .B1(x4), .Y(men_men_n394_));
  NA3        u378(.A(x7), .B(x3), .C(x0), .Y(men_men_n395_));
  NA2        u379(.A(men_men_n230_), .B(x0), .Y(men_men_n396_));
  OAI220     u380(.A0(men_men_n396_), .A1(men_men_n216_), .B0(men_men_n395_), .B1(men_men_n364_), .Y(men_men_n397_));
  AOI210     u381(.A0(men_men_n394_), .A1(men_men_n121_), .B0(men_men_n397_), .Y(men_men_n398_));
  AOI210     u382(.A0(men_men_n398_), .A1(men_men_n392_), .B0(men_men_n25_), .Y(men_men_n399_));
  NA3        u383(.A(men_men_n123_), .B(men_men_n230_), .C(x0), .Y(men_men_n400_));
  OAI210     u384(.A0(men_men_n201_), .A1(men_men_n66_), .B0(men_men_n211_), .Y(men_men_n401_));
  NA3        u385(.A(men_men_n204_), .B(men_men_n232_), .C(x8), .Y(men_men_n402_));
  AOI210     u386(.A0(men_men_n402_), .A1(men_men_n401_), .B0(men_men_n25_), .Y(men_men_n403_));
  NA2        u387(.A(men_men_n403_), .B(men_men_n154_), .Y(men_men_n404_));
  NAi31      u388(.An(men_men_n48_), .B(men_men_n298_), .C(men_men_n181_), .Y(men_men_n405_));
  NA3        u389(.A(men_men_n405_), .B(men_men_n404_), .C(men_men_n400_), .Y(men_men_n406_));
  OAI210     u390(.A0(men_men_n406_), .A1(men_men_n399_), .B0(x6), .Y(men_men_n407_));
  OAI210     u391(.A0(men_men_n168_), .A1(men_men_n46_), .B0(men_men_n138_), .Y(men_men_n408_));
  NA3        u392(.A(men_men_n53_), .B(men_men_n37_), .C(men_men_n30_), .Y(men_men_n409_));
  AOI220     u393(.A0(men_men_n409_), .A1(men_men_n408_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n410_));
  NO2        u394(.A(men_men_n157_), .B(x0), .Y(men_men_n411_));
  AOI220     u395(.A0(men_men_n411_), .A1(men_men_n230_), .B0(men_men_n201_), .B1(men_men_n157_), .Y(men_men_n412_));
  INV        u396(.A(x1), .Y(men_men_n413_));
  OAI210     u397(.A0(men_men_n412_), .A1(x8), .B0(men_men_n413_), .Y(men_men_n414_));
  NOi21      u398(.An(men_men_n128_), .B(men_men_n185_), .Y(men_men_n415_));
  NO2        u399(.A(men_men_n415_), .B(men_men_n18_), .Y(men_men_n416_));
  NO3        u400(.A(x9), .B(men_men_n157_), .C(x0), .Y(men_men_n417_));
  AOI220     u401(.A0(men_men_n417_), .A1(men_men_n251_), .B0(men_men_n373_), .B1(men_men_n157_), .Y(men_men_n418_));
  NA3        u402(.A(men_men_n418_), .B(men_men_n416_), .C(men_men_n48_), .Y(men_men_n419_));
  OAI210     u403(.A0(men_men_n414_), .A1(men_men_n410_), .B0(men_men_n419_), .Y(men_men_n420_));
  NOi31      u404(.An(men_men_n411_), .B(men_men_n31_), .C(x8), .Y(men_men_n421_));
  AOI210     u405(.A0(men_men_n37_), .A1(x9), .B0(men_men_n136_), .Y(men_men_n422_));
  NO3        u406(.A(men_men_n422_), .B(men_men_n128_), .C(men_men_n41_), .Y(men_men_n423_));
  NOi31      u407(.An(x1), .B(x8), .C(x7), .Y(men_men_n424_));
  AOI220     u408(.A0(men_men_n424_), .A1(men_men_n359_), .B0(men_men_n129_), .B1(x3), .Y(men_men_n425_));
  AOI210     u409(.A0(men_men_n273_), .A1(men_men_n58_), .B0(men_men_n127_), .Y(men_men_n426_));
  OAI210     u410(.A0(men_men_n426_), .A1(x3), .B0(men_men_n425_), .Y(men_men_n427_));
  NO3        u411(.A(men_men_n427_), .B(men_men_n423_), .C(x2), .Y(men_men_n428_));
  OAI220     u412(.A0(men_men_n360_), .A1(men_men_n313_), .B0(men_men_n309_), .B1(men_men_n41_), .Y(men_men_n429_));
  INV        u413(.A(men_men_n395_), .Y(men_men_n430_));
  AOI220     u414(.A0(men_men_n430_), .A1(men_men_n93_), .B0(men_men_n429_), .B1(men_men_n157_), .Y(men_men_n431_));
  NO2        u415(.A(men_men_n431_), .B(men_men_n52_), .Y(men_men_n432_));
  NO3        u416(.A(men_men_n432_), .B(men_men_n428_), .C(men_men_n421_), .Y(men_men_n433_));
  AOI210     u417(.A0(men_men_n433_), .A1(men_men_n420_), .B0(men_men_n25_), .Y(men_men_n434_));
  NA4        u418(.A(men_men_n30_), .B(men_men_n93_), .C(x2), .D(men_men_n17_), .Y(men_men_n435_));
  NO3        u419(.A(men_men_n66_), .B(men_men_n18_), .C(x0), .Y(men_men_n436_));
  NA2        u420(.A(men_men_n436_), .B(men_men_n274_), .Y(men_men_n437_));
  NO2        u421(.A(men_men_n437_), .B(men_men_n105_), .Y(men_men_n438_));
  NO3        u422(.A(men_men_n278_), .B(men_men_n180_), .C(men_men_n38_), .Y(men_men_n439_));
  OAI210     u423(.A0(men_men_n439_), .A1(men_men_n438_), .B0(x7), .Y(men_men_n440_));
  NA2        u424(.A(men_men_n235_), .B(x7), .Y(men_men_n441_));
  NA3        u425(.A(men_men_n441_), .B(men_men_n156_), .C(men_men_n137_), .Y(men_men_n442_));
  NA3        u426(.A(men_men_n442_), .B(men_men_n440_), .C(men_men_n435_), .Y(men_men_n443_));
  OAI210     u427(.A0(men_men_n443_), .A1(men_men_n434_), .B0(men_men_n35_), .Y(men_men_n444_));
  NO2        u428(.A(men_men_n417_), .B(men_men_n211_), .Y(men_men_n445_));
  NO4        u429(.A(men_men_n445_), .B(men_men_n77_), .C(x4), .D(men_men_n52_), .Y(men_men_n446_));
  AOI220     u430(.A0(men_men_n371_), .A1(men_men_n93_), .B0(men_men_n155_), .B1(men_men_n204_), .Y(men_men_n447_));
  NA2        u431(.A(men_men_n447_), .B(men_men_n91_), .Y(men_men_n448_));
  NA2        u432(.A(men_men_n448_), .B(men_men_n181_), .Y(men_men_n449_));
  OAI220     u433(.A0(men_men_n287_), .A1(men_men_n67_), .B0(men_men_n165_), .B1(men_men_n41_), .Y(men_men_n450_));
  NA2        u434(.A(x3), .B(men_men_n52_), .Y(men_men_n451_));
  AOI210     u435(.A0(men_men_n169_), .A1(men_men_n27_), .B0(men_men_n72_), .Y(men_men_n452_));
  OAI210     u436(.A0(men_men_n154_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n453_));
  NO3        u437(.A(men_men_n424_), .B(x3), .C(men_men_n52_), .Y(men_men_n454_));
  AOI210     u438(.A0(men_men_n454_), .A1(men_men_n453_), .B0(men_men_n452_), .Y(men_men_n455_));
  OAI210     u439(.A0(men_men_n158_), .A1(men_men_n451_), .B0(men_men_n455_), .Y(men_men_n456_));
  AOI220     u440(.A0(men_men_n456_), .A1(x0), .B0(men_men_n450_), .B1(men_men_n138_), .Y(men_men_n457_));
  AOI210     u441(.A0(men_men_n457_), .A1(men_men_n449_), .B0(men_men_n241_), .Y(men_men_n458_));
  INV        u442(.A(x5), .Y(men_men_n459_));
  NO4        u443(.A(men_men_n108_), .B(men_men_n459_), .C(men_men_n58_), .D(men_men_n31_), .Y(men_men_n460_));
  NO3        u444(.A(men_men_n460_), .B(men_men_n458_), .C(men_men_n446_), .Y(men_men_n461_));
  NA3        u445(.A(men_men_n461_), .B(men_men_n444_), .C(men_men_n407_), .Y(men_men_n462_));
  AOI210     u446(.A0(men_men_n389_), .A1(men_men_n25_), .B0(men_men_n462_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule