//Benchmark atmr_intb_466_0.0313

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n349_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n364_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n419_, mai_mai_n420_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n368_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  AOI220     o035(.A0(x11), .A1(ori_ori_n48_), .B0(x10), .B1(ori_ori_n57_), .Y(ori_ori_n58_));
  INV        o036(.A(ori_ori_n55_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(ori_ori_n24_), .Y(ori_ori_n61_));
  OAI220     o039(.A0(ori_ori_n61_), .A1(ori_ori_n59_), .B0(ori_ori_n58_), .B1(ori_ori_n56_), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n63_));
  OAI210     o041(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n63_), .Y(ori_ori_n64_));
  AOI220     o042(.A0(ori_ori_n64_), .A1(ori_ori_n55_), .B0(ori_ori_n62_), .B1(ori_ori_n31_), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n65_), .B(x05), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n57_), .B(ori_ori_n23_), .Y(ori_ori_n67_));
  NA2        o045(.A(x09), .B(x05), .Y(ori_ori_n68_));
  NA2        o046(.A(x10), .B(x06), .Y(ori_ori_n69_));
  NA3        o047(.A(ori_ori_n69_), .B(ori_ori_n68_), .C(ori_ori_n28_), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n57_), .B(ori_ori_n41_), .Y(ori_ori_n71_));
  OAI210     o049(.A0(ori_ori_n70_), .A1(ori_ori_n67_), .B0(x03), .Y(ori_ori_n72_));
  NOi31      o050(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n73_));
  INV        o051(.A(ori_ori_n24_), .Y(ori_ori_n74_));
  NO2        o052(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n75_), .B(ori_ori_n36_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n75_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n77_));
  INV        o055(.A(ori_ori_n77_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n79_));
  NO2        o057(.A(x08), .B(x01), .Y(ori_ori_n80_));
  OAI210     o058(.A0(ori_ori_n80_), .A1(ori_ori_n79_), .B0(ori_ori_n35_), .Y(ori_ori_n81_));
  NA2        o059(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n82_));
  NO3        o060(.A(ori_ori_n81_), .B(ori_ori_n78_), .C(ori_ori_n74_), .Y(ori_ori_n83_));
  AN2        o061(.A(ori_ori_n83_), .B(ori_ori_n72_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n81_), .Y(ori_ori_n85_));
  NA2        o063(.A(x11), .B(x00), .Y(ori_ori_n86_));
  NO2        o064(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n87_));
  NOi21      o065(.An(ori_ori_n86_), .B(ori_ori_n87_), .Y(ori_ori_n88_));
  INV        o066(.A(ori_ori_n88_), .Y(ori_ori_n89_));
  NOi21      o067(.An(x01), .B(x10), .Y(ori_ori_n90_));
  NO2        o068(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n91_));
  NO3        o069(.A(ori_ori_n91_), .B(ori_ori_n90_), .C(x06), .Y(ori_ori_n92_));
  NA2        o070(.A(ori_ori_n92_), .B(ori_ori_n27_), .Y(ori_ori_n93_));
  OAI210     o071(.A0(ori_ori_n89_), .A1(x07), .B0(ori_ori_n93_), .Y(ori_ori_n94_));
  NO3        o072(.A(ori_ori_n94_), .B(ori_ori_n84_), .C(ori_ori_n66_), .Y(ori01));
  INV        o073(.A(x12), .Y(ori_ori_n96_));
  INV        o074(.A(x13), .Y(ori_ori_n97_));
  NA2        o075(.A(x08), .B(x04), .Y(ori_ori_n98_));
  NA2        o076(.A(ori_ori_n90_), .B(ori_ori_n28_), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n99_), .B(ori_ori_n68_), .Y(ori_ori_n100_));
  NO2        o078(.A(x10), .B(x01), .Y(ori_ori_n101_));
  NO2        o079(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n102_));
  NO2        o080(.A(ori_ori_n102_), .B(ori_ori_n101_), .Y(ori_ori_n103_));
  NA2        o081(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n104_), .B(ori_ori_n36_), .Y(ori_ori_n105_));
  AOI210     o083(.A0(ori_ori_n105_), .A1(ori_ori_n103_), .B0(ori_ori_n100_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(ori_ori_n97_), .Y(ori_ori_n107_));
  NO2        o085(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n108_));
  NOi21      o086(.An(ori_ori_n108_), .B(ori_ori_n54_), .Y(ori_ori_n109_));
  INV        o087(.A(x13), .Y(ori_ori_n110_));
  NA2        o088(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n111_));
  NA2        o089(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n112_));
  NO2        o090(.A(ori_ori_n112_), .B(x05), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n35_), .B(ori_ori_n53_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n114_), .B(ori_ori_n97_), .Y(ori_ori_n115_));
  AOI210     o093(.A0(ori_ori_n115_), .A1(ori_ori_n76_), .B0(ori_ori_n109_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n116_), .B(ori_ori_n69_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n118_));
  NA2        o096(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n122_), .B(ori_ori_n120_), .Y(ori_ori_n123_));
  NO3        o101(.A(ori_ori_n123_), .B(x06), .C(x03), .Y(ori_ori_n124_));
  NO3        o102(.A(ori_ori_n124_), .B(ori_ori_n117_), .C(ori_ori_n107_), .Y(ori_ori_n125_));
  NA2        o103(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n126_));
  OAI210     o104(.A0(ori_ori_n80_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n127_), .B(ori_ori_n126_), .Y(ori_ori_n128_));
  NO2        o106(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n130_));
  NO2        o108(.A(x09), .B(x05), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n131_), .B(ori_ori_n47_), .Y(ori_ori_n132_));
  NO2        o110(.A(ori_ori_n103_), .B(ori_ori_n49_), .Y(ori_ori_n133_));
  NA2        o111(.A(x09), .B(x00), .Y(ori_ori_n134_));
  NA2        o112(.A(ori_ori_n108_), .B(ori_ori_n134_), .Y(ori_ori_n135_));
  NA2        o113(.A(ori_ori_n73_), .B(ori_ori_n50_), .Y(ori_ori_n136_));
  AOI210     o114(.A0(ori_ori_n136_), .A1(ori_ori_n135_), .B0(ori_ori_n130_), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n137_), .B(ori_ori_n133_), .Y(ori_ori_n138_));
  NO2        o116(.A(x03), .B(x02), .Y(ori_ori_n139_));
  NA2        o117(.A(ori_ori_n81_), .B(ori_ori_n97_), .Y(ori_ori_n140_));
  OAI210     o118(.A0(ori_ori_n140_), .A1(ori_ori_n109_), .B0(ori_ori_n139_), .Y(ori_ori_n141_));
  OA210      o119(.A0(ori_ori_n138_), .A1(x11), .B0(ori_ori_n141_), .Y(ori_ori_n142_));
  OAI210     o120(.A0(ori_ori_n125_), .A1(ori_ori_n23_), .B0(ori_ori_n142_), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n103_), .B(ori_ori_n40_), .Y(ori_ori_n144_));
  NAi21      o122(.An(x06), .B(x10), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n144_), .B(ori_ori_n41_), .Y(ori_ori_n146_));
  NO2        o124(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n147_));
  NA2        o125(.A(ori_ori_n97_), .B(x01), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n148_), .B(x08), .Y(ori_ori_n149_));
  OAI210     o127(.A0(x05), .A1(ori_ori_n149_), .B0(ori_ori_n50_), .Y(ori_ori_n150_));
  AOI210     o128(.A0(ori_ori_n150_), .A1(ori_ori_n147_), .B0(ori_ori_n48_), .Y(ori_ori_n151_));
  AOI210     o129(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n152_));
  OAI210     o130(.A0(ori_ori_n151_), .A1(ori_ori_n146_), .B0(ori_ori_n152_), .Y(ori_ori_n153_));
  NA2        o131(.A(x10), .B(x05), .Y(ori_ori_n154_));
  NO2        o132(.A(x09), .B(x01), .Y(ori_ori_n155_));
  INV        o133(.A(ori_ori_n25_), .Y(ori_ori_n156_));
  NAi21      o134(.An(x13), .B(x00), .Y(ori_ori_n157_));
  AOI210     o135(.A0(ori_ori_n29_), .A1(ori_ori_n48_), .B0(ori_ori_n157_), .Y(ori_ori_n158_));
  AOI220     o136(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(ori_ori_n159_));
  OAI210     o137(.A0(ori_ori_n154_), .A1(ori_ori_n35_), .B0(ori_ori_n159_), .Y(ori_ori_n160_));
  AN2        o138(.A(ori_ori_n160_), .B(ori_ori_n158_), .Y(ori_ori_n161_));
  NO2        o139(.A(ori_ori_n157_), .B(ori_ori_n36_), .Y(ori_ori_n162_));
  INV        o140(.A(ori_ori_n162_), .Y(ori_ori_n163_));
  OAI210     o141(.A0(ori_ori_n406_), .A1(ori_ori_n161_), .B0(ori_ori_n156_), .Y(ori_ori_n164_));
  NOi21      o142(.An(x09), .B(x00), .Y(ori_ori_n165_));
  NO3        o143(.A(ori_ori_n79_), .B(ori_ori_n165_), .C(ori_ori_n47_), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n166_), .B(ori_ori_n119_), .Y(ori_ori_n167_));
  NA2        o145(.A(x10), .B(x08), .Y(ori_ori_n168_));
  INV        o146(.A(ori_ori_n168_), .Y(ori_ori_n169_));
  NA2        o147(.A(x06), .B(x05), .Y(ori_ori_n170_));
  OAI210     o148(.A0(ori_ori_n170_), .A1(ori_ori_n35_), .B0(ori_ori_n96_), .Y(ori_ori_n171_));
  AOI210     o149(.A0(ori_ori_n169_), .A1(ori_ori_n54_), .B0(ori_ori_n171_), .Y(ori_ori_n172_));
  NA2        o150(.A(ori_ori_n172_), .B(ori_ori_n167_), .Y(ori_ori_n173_));
  NO2        o151(.A(ori_ori_n97_), .B(x12), .Y(ori_ori_n174_));
  AOI210     o152(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n174_), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n90_), .B(ori_ori_n50_), .Y(ori_ori_n176_));
  NO2        o154(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n177_));
  NA2        o155(.A(ori_ori_n177_), .B(x02), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n178_), .B(ori_ori_n176_), .Y(ori_ori_n179_));
  AOI210     o157(.A0(ori_ori_n175_), .A1(ori_ori_n173_), .B0(ori_ori_n179_), .Y(ori_ori_n180_));
  NA3        o158(.A(ori_ori_n180_), .B(ori_ori_n164_), .C(ori_ori_n153_), .Y(ori_ori_n181_));
  AOI210     o159(.A0(ori_ori_n143_), .A1(ori_ori_n96_), .B0(ori_ori_n181_), .Y(ori_ori_n182_));
  INV        o160(.A(ori_ori_n70_), .Y(ori_ori_n183_));
  NA2        o161(.A(ori_ori_n183_), .B(ori_ori_n128_), .Y(ori_ori_n184_));
  NA2        o162(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n185_));
  NA2        o163(.A(ori_ori_n185_), .B(ori_ori_n127_), .Y(ori_ori_n186_));
  NO2        o164(.A(ori_ori_n118_), .B(x06), .Y(ori_ori_n187_));
  INV        o165(.A(ori_ori_n187_), .Y(ori_ori_n188_));
  AOI210     o166(.A0(ori_ori_n188_), .A1(ori_ori_n184_), .B0(x12), .Y(ori_ori_n189_));
  INV        o167(.A(ori_ori_n73_), .Y(ori_ori_n190_));
  NO2        o168(.A(ori_ori_n90_), .B(x06), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n191_), .B(ori_ori_n41_), .Y(ori_ori_n192_));
  INV        o170(.A(ori_ori_n130_), .Y(ori_ori_n193_));
  OAI210     o171(.A0(ori_ori_n193_), .A1(ori_ori_n192_), .B0(x02), .Y(ori_ori_n194_));
  AOI210     o172(.A0(ori_ori_n194_), .A1(ori_ori_n53_), .B0(ori_ori_n23_), .Y(ori_ori_n195_));
  OAI210     o173(.A0(ori_ori_n189_), .A1(ori_ori_n53_), .B0(ori_ori_n195_), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n130_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n198_));
  OAI210     o176(.A0(ori_ori_n75_), .A1(ori_ori_n36_), .B0(ori_ori_n111_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n97_), .B(x03), .Y(ori_ori_n200_));
  NA2        o178(.A(ori_ori_n200_), .B(ori_ori_n199_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n202_));
  INV        o180(.A(ori_ori_n145_), .Y(ori_ori_n203_));
  NOi21      o181(.An(x13), .B(x04), .Y(ori_ori_n204_));
  NO3        o182(.A(ori_ori_n204_), .B(ori_ori_n73_), .C(ori_ori_n165_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n205_), .B(x05), .Y(ori_ori_n206_));
  AOI220     o184(.A0(ori_ori_n206_), .A1(ori_ori_n202_), .B0(ori_ori_n203_), .B1(ori_ori_n53_), .Y(ori_ori_n207_));
  OAI210     o185(.A0(ori_ori_n201_), .A1(ori_ori_n197_), .B0(ori_ori_n207_), .Y(ori_ori_n208_));
  INV        o186(.A(ori_ori_n87_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n209_), .B(x12), .Y(ori_ori_n210_));
  NA2        o188(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n212_));
  OAI210     o190(.A0(ori_ori_n212_), .A1(ori_ori_n160_), .B0(ori_ori_n158_), .Y(ori_ori_n213_));
  AOI210     o191(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n214_));
  NO2        o192(.A(x06), .B(x00), .Y(ori_ori_n215_));
  NO3        o193(.A(ori_ori_n215_), .B(ori_ori_n214_), .C(ori_ori_n41_), .Y(ori_ori_n216_));
  OAI210     o194(.A0(ori_ori_n98_), .A1(ori_ori_n134_), .B0(ori_ori_n69_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n217_), .B(ori_ori_n216_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n219_), .B(x03), .Y(ori_ori_n220_));
  OA210      o198(.A0(ori_ori_n220_), .A1(ori_ori_n218_), .B0(ori_ori_n213_), .Y(ori_ori_n221_));
  NA2        o199(.A(x13), .B(ori_ori_n96_), .Y(ori_ori_n222_));
  NA3        o200(.A(ori_ori_n222_), .B(ori_ori_n171_), .C(ori_ori_n88_), .Y(ori_ori_n223_));
  OAI210     o201(.A0(ori_ori_n221_), .A1(ori_ori_n211_), .B0(ori_ori_n223_), .Y(ori_ori_n224_));
  AOI210     o202(.A0(ori_ori_n210_), .A1(ori_ori_n208_), .B0(ori_ori_n224_), .Y(ori_ori_n225_));
  AOI210     o203(.A0(ori_ori_n225_), .A1(ori_ori_n196_), .B0(x07), .Y(ori_ori_n226_));
  NA2        o204(.A(ori_ori_n68_), .B(ori_ori_n29_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n204_), .B(ori_ori_n165_), .Y(ori_ori_n228_));
  AOI210     o206(.A0(ori_ori_n228_), .A1(ori_ori_n136_), .B0(ori_ori_n227_), .Y(ori_ori_n229_));
  NO2        o207(.A(ori_ori_n97_), .B(x06), .Y(ori_ori_n230_));
  INV        o208(.A(ori_ori_n230_), .Y(ori_ori_n231_));
  NO2        o209(.A(x08), .B(x05), .Y(ori_ori_n232_));
  NO2        o210(.A(ori_ori_n232_), .B(ori_ori_n214_), .Y(ori_ori_n233_));
  NA2        o211(.A(x13), .B(ori_ori_n31_), .Y(ori_ori_n234_));
  OAI210     o212(.A0(ori_ori_n233_), .A1(ori_ori_n231_), .B0(ori_ori_n234_), .Y(ori_ori_n235_));
  NO2        o213(.A(x12), .B(x02), .Y(ori_ori_n236_));
  INV        o214(.A(ori_ori_n236_), .Y(ori_ori_n237_));
  NO2        o215(.A(ori_ori_n237_), .B(ori_ori_n209_), .Y(ori_ori_n238_));
  OA210      o216(.A0(ori_ori_n235_), .A1(ori_ori_n229_), .B0(ori_ori_n238_), .Y(ori_ori_n239_));
  NA2        o217(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n240_));
  NO2        o218(.A(ori_ori_n240_), .B(x01), .Y(ori_ori_n241_));
  NOi21      o219(.An(ori_ori_n80_), .B(ori_ori_n111_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n242_), .B(ori_ori_n241_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n243_), .B(ori_ori_n29_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n230_), .B(ori_ori_n199_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n97_), .B(x04), .Y(ori_ori_n246_));
  OAI210     o224(.A0(x02), .A1(ori_ori_n110_), .B0(ori_ori_n245_), .Y(ori_ori_n247_));
  NO3        o225(.A(ori_ori_n86_), .B(x12), .C(x03), .Y(ori_ori_n248_));
  OAI210     o226(.A0(ori_ori_n247_), .A1(ori_ori_n244_), .B0(ori_ori_n248_), .Y(ori_ori_n249_));
  AOI210     o227(.A0(ori_ori_n176_), .A1(ori_ori_n170_), .B0(ori_ori_n98_), .Y(ori_ori_n250_));
  NOi21      o228(.An(ori_ori_n227_), .B(ori_ori_n191_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n252_));
  OAI210     o230(.A0(ori_ori_n251_), .A1(ori_ori_n250_), .B0(ori_ori_n252_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n254_));
  NO2        o232(.A(ori_ori_n211_), .B(ori_ori_n28_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n197_), .B(ori_ori_n255_), .Y(ori_ori_n256_));
  NA3        o234(.A(ori_ori_n256_), .B(ori_ori_n253_), .C(ori_ori_n249_), .Y(ori_ori_n257_));
  NO3        o235(.A(ori_ori_n257_), .B(ori_ori_n239_), .C(ori_ori_n226_), .Y(ori_ori_n258_));
  OAI210     o236(.A0(ori_ori_n182_), .A1(ori_ori_n57_), .B0(ori_ori_n258_), .Y(ori02));
  AOI210     o237(.A0(ori_ori_n126_), .A1(ori_ori_n81_), .B0(ori_ori_n121_), .Y(ori_ori_n260_));
  NOi21      o238(.An(ori_ori_n205_), .B(ori_ori_n155_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n97_), .B(ori_ori_n35_), .Y(ori_ori_n262_));
  NA3        o240(.A(ori_ori_n262_), .B(ori_ori_n169_), .C(ori_ori_n52_), .Y(ori_ori_n263_));
  OAI210     o241(.A0(ori_ori_n261_), .A1(ori_ori_n32_), .B0(ori_ori_n263_), .Y(ori_ori_n264_));
  OAI210     o242(.A0(ori_ori_n264_), .A1(ori_ori_n260_), .B0(ori_ori_n154_), .Y(ori_ori_n265_));
  INV        o243(.A(ori_ori_n154_), .Y(ori_ori_n266_));
  OAI220     o244(.A0(ori_ori_n50_), .A1(ori_ori_n97_), .B0(ori_ori_n81_), .B1(ori_ori_n50_), .Y(ori_ori_n267_));
  AOI220     o245(.A0(ori_ori_n267_), .A1(ori_ori_n266_), .B0(ori_ori_n140_), .B1(ori_ori_n139_), .Y(ori_ori_n268_));
  AOI210     o246(.A0(ori_ori_n268_), .A1(ori_ori_n265_), .B0(ori_ori_n48_), .Y(ori_ori_n269_));
  NO2        o247(.A(x05), .B(x02), .Y(ori_ori_n270_));
  OAI210     o248(.A0(ori_ori_n186_), .A1(ori_ori_n165_), .B0(ori_ori_n270_), .Y(ori_ori_n271_));
  AOI220     o249(.A0(ori_ori_n232_), .A1(ori_ori_n54_), .B0(ori_ori_n52_), .B1(ori_ori_n36_), .Y(ori_ori_n272_));
  NOi21      o250(.An(ori_ori_n262_), .B(ori_ori_n272_), .Y(ori_ori_n273_));
  INV        o251(.A(ori_ori_n273_), .Y(ori_ori_n274_));
  AOI210     o252(.A0(ori_ori_n274_), .A1(ori_ori_n271_), .B0(ori_ori_n130_), .Y(ori_ori_n275_));
  NAi21      o253(.An(ori_ori_n206_), .B(ori_ori_n201_), .Y(ori_ori_n276_));
  NO2        o254(.A(ori_ori_n219_), .B(ori_ori_n47_), .Y(ori_ori_n277_));
  NA2        o255(.A(ori_ori_n277_), .B(ori_ori_n276_), .Y(ori_ori_n278_));
  AN2        o256(.A(ori_ori_n200_), .B(ori_ori_n199_), .Y(ori_ori_n279_));
  OAI210     o257(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n280_));
  NA2        o258(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n281_));
  OA210      o259(.A0(ori_ori_n281_), .A1(x08), .B0(ori_ori_n132_), .Y(ori_ori_n282_));
  AOI210     o260(.A0(ori_ori_n282_), .A1(ori_ori_n127_), .B0(ori_ori_n280_), .Y(ori_ori_n283_));
  OAI210     o261(.A0(ori_ori_n283_), .A1(ori_ori_n279_), .B0(ori_ori_n91_), .Y(ori_ori_n284_));
  NA3        o262(.A(ori_ori_n91_), .B(ori_ori_n80_), .C(ori_ori_n198_), .Y(ori_ori_n285_));
  NA3        o263(.A(ori_ori_n90_), .B(ori_ori_n79_), .C(ori_ori_n42_), .Y(ori_ori_n286_));
  AOI210     o264(.A0(ori_ori_n286_), .A1(ori_ori_n285_), .B0(x04), .Y(ori_ori_n287_));
  INV        o265(.A(ori_ori_n139_), .Y(ori_ori_n288_));
  OAI220     o266(.A0(ori_ori_n233_), .A1(ori_ori_n99_), .B0(ori_ori_n288_), .B1(ori_ori_n120_), .Y(ori_ori_n289_));
  AOI210     o267(.A0(ori_ori_n289_), .A1(x13), .B0(ori_ori_n287_), .Y(ori_ori_n290_));
  NA3        o268(.A(ori_ori_n290_), .B(ori_ori_n284_), .C(ori_ori_n278_), .Y(ori_ori_n291_));
  NO3        o269(.A(ori_ori_n291_), .B(ori_ori_n275_), .C(ori_ori_n269_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n129_), .B(x03), .Y(ori_ori_n293_));
  INV        o271(.A(ori_ori_n157_), .Y(ori_ori_n294_));
  OAI210     o272(.A0(ori_ori_n50_), .A1(ori_ori_n35_), .B0(ori_ori_n36_), .Y(ori_ori_n295_));
  AOI220     o273(.A0(ori_ori_n295_), .A1(ori_ori_n294_), .B0(ori_ori_n177_), .B1(x08), .Y(ori_ori_n296_));
  OAI210     o274(.A0(ori_ori_n296_), .A1(ori_ori_n254_), .B0(ori_ori_n293_), .Y(ori_ori_n297_));
  NA2        o275(.A(ori_ori_n297_), .B(ori_ori_n101_), .Y(ori_ori_n298_));
  INV        o276(.A(ori_ori_n52_), .Y(ori_ori_n299_));
  OAI220     o277(.A0(ori_ori_n246_), .A1(ori_ori_n299_), .B0(ori_ori_n121_), .B1(ori_ori_n28_), .Y(ori_ori_n300_));
  NA2        o278(.A(ori_ori_n300_), .B(ori_ori_n102_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n246_), .B(ori_ori_n96_), .Y(ori_ori_n302_));
  NA2        o280(.A(ori_ori_n96_), .B(ori_ori_n41_), .Y(ori_ori_n303_));
  NA3        o281(.A(ori_ori_n303_), .B(ori_ori_n302_), .C(ori_ori_n120_), .Y(ori_ori_n304_));
  NA4        o282(.A(ori_ori_n304_), .B(ori_ori_n301_), .C(ori_ori_n298_), .D(ori_ori_n48_), .Y(ori_ori_n305_));
  INV        o283(.A(ori_ori_n177_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n307_));
  OAI220     o285(.A0(ori_ori_n307_), .A1(ori_ori_n407_), .B0(ori_ori_n306_), .B1(ori_ori_n55_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n308_), .B(x02), .Y(ori_ori_n309_));
  INV        o287(.A(ori_ori_n212_), .Y(ori_ori_n310_));
  NA2        o288(.A(ori_ori_n174_), .B(x04), .Y(ori_ori_n311_));
  NO2        o289(.A(ori_ori_n311_), .B(ori_ori_n310_), .Y(ori_ori_n312_));
  NO3        o290(.A(ori_ori_n159_), .B(x13), .C(ori_ori_n31_), .Y(ori_ori_n313_));
  OAI210     o291(.A0(ori_ori_n313_), .A1(ori_ori_n312_), .B0(ori_ori_n91_), .Y(ori_ori_n314_));
  NO3        o292(.A(ori_ori_n174_), .B(ori_ori_n147_), .C(ori_ori_n51_), .Y(ori_ori_n315_));
  OAI210     o293(.A0(ori_ori_n134_), .A1(ori_ori_n36_), .B0(ori_ori_n96_), .Y(ori_ori_n316_));
  OAI210     o294(.A0(ori_ori_n316_), .A1(ori_ori_n166_), .B0(ori_ori_n315_), .Y(ori_ori_n317_));
  NA4        o295(.A(ori_ori_n317_), .B(ori_ori_n314_), .C(ori_ori_n309_), .D(x06), .Y(ori_ori_n318_));
  NA2        o296(.A(x09), .B(x03), .Y(ori_ori_n319_));
  OAI220     o297(.A0(ori_ori_n319_), .A1(ori_ori_n119_), .B0(ori_ori_n185_), .B1(ori_ori_n60_), .Y(ori_ori_n320_));
  OAI220     o298(.A0(ori_ori_n148_), .A1(x09), .B0(x08), .B1(ori_ori_n41_), .Y(ori_ori_n321_));
  NA2        o299(.A(ori_ori_n321_), .B(ori_ori_n197_), .Y(ori_ori_n322_));
  NO3        o300(.A(ori_ori_n108_), .B(ori_ori_n119_), .C(ori_ori_n38_), .Y(ori_ori_n323_));
  INV        o301(.A(ori_ori_n323_), .Y(ori_ori_n324_));
  OAI210     o302(.A0(ori_ori_n322_), .A1(ori_ori_n28_), .B0(ori_ori_n324_), .Y(ori_ori_n325_));
  AO220      o303(.A0(ori_ori_n325_), .A1(x04), .B0(ori_ori_n320_), .B1(x05), .Y(ori_ori_n326_));
  AOI210     o304(.A0(ori_ori_n318_), .A1(ori_ori_n305_), .B0(ori_ori_n326_), .Y(ori_ori_n327_));
  OAI210     o305(.A0(ori_ori_n292_), .A1(x12), .B0(ori_ori_n327_), .Y(ori03));
  OR2        o306(.A(ori_ori_n42_), .B(ori_ori_n198_), .Y(ori_ori_n329_));
  AOI210     o307(.A0(ori_ori_n140_), .A1(ori_ori_n96_), .B0(ori_ori_n329_), .Y(ori_ori_n330_));
  AO210      o308(.A0(ori_ori_n310_), .A1(ori_ori_n82_), .B0(ori_ori_n311_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n174_), .B(ori_ori_n139_), .Y(ori_ori_n332_));
  NA3        o310(.A(ori_ori_n332_), .B(ori_ori_n331_), .C(ori_ori_n178_), .Y(ori_ori_n333_));
  OAI210     o311(.A0(ori_ori_n333_), .A1(ori_ori_n330_), .B0(x05), .Y(ori_ori_n334_));
  NA2        o312(.A(ori_ori_n329_), .B(x05), .Y(ori_ori_n335_));
  AOI210     o313(.A0(ori_ori_n127_), .A1(ori_ori_n190_), .B0(ori_ori_n335_), .Y(ori_ori_n336_));
  AOI210     o314(.A0(ori_ori_n200_), .A1(ori_ori_n76_), .B0(ori_ori_n113_), .Y(ori_ori_n337_));
  OAI220     o315(.A0(ori_ori_n337_), .A1(ori_ori_n55_), .B0(ori_ori_n281_), .B1(ori_ori_n272_), .Y(ori_ori_n338_));
  OAI210     o316(.A0(ori_ori_n338_), .A1(ori_ori_n336_), .B0(ori_ori_n96_), .Y(ori_ori_n339_));
  AOI210     o317(.A0(ori_ori_n132_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n340_));
  NO2        o318(.A(ori_ori_n155_), .B(ori_ori_n122_), .Y(ori_ori_n341_));
  OAI220     o319(.A0(ori_ori_n341_), .A1(ori_ori_n37_), .B0(ori_ori_n135_), .B1(x13), .Y(ori_ori_n342_));
  OAI210     o320(.A0(ori_ori_n342_), .A1(ori_ori_n340_), .B0(x04), .Y(ori_ori_n343_));
  NO3        o321(.A(ori_ori_n303_), .B(ori_ori_n81_), .C(ori_ori_n55_), .Y(ori_ori_n344_));
  AOI210     o322(.A0(ori_ori_n163_), .A1(ori_ori_n96_), .B0(ori_ori_n132_), .Y(ori_ori_n345_));
  OA210      o323(.A0(ori_ori_n149_), .A1(x12), .B0(ori_ori_n122_), .Y(ori_ori_n346_));
  NO3        o324(.A(ori_ori_n346_), .B(ori_ori_n345_), .C(ori_ori_n344_), .Y(ori_ori_n347_));
  NA4        o325(.A(ori_ori_n347_), .B(ori_ori_n343_), .C(ori_ori_n339_), .D(ori_ori_n334_), .Y(ori04));
  NO2        o326(.A(ori_ori_n85_), .B(ori_ori_n39_), .Y(ori_ori_n349_));
  XO2        o327(.A(ori_ori_n349_), .B(ori_ori_n222_), .Y(ori05));
  AOI210     o328(.A0(ori_ori_n68_), .A1(ori_ori_n51_), .B0(ori_ori_n187_), .Y(ori_ori_n351_));
  AOI210     o329(.A0(ori_ori_n351_), .A1(ori_ori_n280_), .B0(ori_ori_n25_), .Y(ori_ori_n352_));
  NA3        o330(.A(ori_ori_n130_), .B(ori_ori_n121_), .C(ori_ori_n31_), .Y(ori_ori_n353_));
  NA2        o331(.A(ori_ori_n203_), .B(ori_ori_n53_), .Y(ori_ori_n354_));
  AOI210     o332(.A0(ori_ori_n354_), .A1(ori_ori_n353_), .B0(ori_ori_n24_), .Y(ori_ori_n355_));
  OAI210     o333(.A0(ori_ori_n355_), .A1(ori_ori_n352_), .B0(ori_ori_n96_), .Y(ori_ori_n356_));
  NA2        o334(.A(x11), .B(ori_ori_n31_), .Y(ori_ori_n357_));
  NA2        o335(.A(ori_ori_n23_), .B(ori_ori_n28_), .Y(ori_ori_n358_));
  NA2        o336(.A(ori_ori_n227_), .B(x03), .Y(ori_ori_n359_));
  OAI220     o337(.A0(ori_ori_n359_), .A1(ori_ori_n358_), .B0(ori_ori_n357_), .B1(ori_ori_n77_), .Y(ori_ori_n360_));
  OAI210     o338(.A0(ori_ori_n26_), .A1(ori_ori_n96_), .B0(x07), .Y(ori_ori_n361_));
  AOI210     o339(.A0(ori_ori_n360_), .A1(x06), .B0(ori_ori_n361_), .Y(ori_ori_n362_));
  AOI210     o340(.A0(ori_ori_n77_), .A1(ori_ori_n31_), .B0(ori_ori_n51_), .Y(ori_ori_n363_));
  NO3        o341(.A(ori_ori_n363_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n364_));
  AOI210     o342(.A0(ori_ori_n405_), .A1(ori_ori_n359_), .B0(ori_ori_n230_), .Y(ori_ori_n365_));
  OR2        o343(.A(ori_ori_n365_), .B(ori_ori_n211_), .Y(ori_ori_n366_));
  NA2        o344(.A(ori_ori_n215_), .B(ori_ori_n209_), .Y(ori_ori_n367_));
  NA2        o345(.A(ori_ori_n367_), .B(ori_ori_n366_), .Y(ori_ori_n368_));
  OAI210     o346(.A0(ori_ori_n368_), .A1(ori_ori_n364_), .B0(ori_ori_n96_), .Y(ori_ori_n369_));
  NA2        o347(.A(ori_ori_n33_), .B(ori_ori_n96_), .Y(ori_ori_n370_));
  AOI210     o348(.A0(ori_ori_n370_), .A1(ori_ori_n87_), .B0(x07), .Y(ori_ori_n371_));
  AOI220     o349(.A0(ori_ori_n371_), .A1(ori_ori_n369_), .B0(ori_ori_n362_), .B1(ori_ori_n356_), .Y(ori_ori_n372_));
  AOI210     o350(.A0(ori_ori_n311_), .A1(ori_ori_n104_), .B0(ori_ori_n236_), .Y(ori_ori_n373_));
  NOi21      o351(.An(ori_ori_n293_), .B(ori_ori_n122_), .Y(ori_ori_n374_));
  NO2        o352(.A(ori_ori_n374_), .B(ori_ori_n237_), .Y(ori_ori_n375_));
  OAI210     o353(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n376_));
  AOI210     o354(.A0(ori_ori_n222_), .A1(ori_ori_n47_), .B0(ori_ori_n376_), .Y(ori_ori_n377_));
  NO4        o355(.A(ori_ori_n377_), .B(ori_ori_n375_), .C(ori_ori_n373_), .D(x08), .Y(ori_ori_n378_));
  NO2        o356(.A(ori_ori_n121_), .B(ori_ori_n28_), .Y(ori_ori_n379_));
  NO2        o357(.A(ori_ori_n379_), .B(ori_ori_n241_), .Y(ori_ori_n380_));
  OR3        o358(.A(ori_ori_n380_), .B(x12), .C(x03), .Y(ori_ori_n381_));
  NA3        o359(.A(ori_ori_n306_), .B(ori_ori_n114_), .C(x12), .Y(ori_ori_n382_));
  AO210      o360(.A0(ori_ori_n306_), .A1(ori_ori_n114_), .B0(ori_ori_n222_), .Y(ori_ori_n383_));
  NA4        o361(.A(ori_ori_n383_), .B(ori_ori_n382_), .C(ori_ori_n381_), .D(x08), .Y(ori_ori_n384_));
  INV        o362(.A(ori_ori_n384_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n378_), .B(ori_ori_n385_), .Y(ori_ori_n386_));
  INV        o364(.A(x03), .Y(ori_ori_n387_));
  NO2        o365(.A(ori_ori_n131_), .B(ori_ori_n43_), .Y(ori_ori_n388_));
  OAI210     o366(.A0(ori_ori_n388_), .A1(ori_ori_n387_), .B0(ori_ori_n162_), .Y(ori_ori_n389_));
  NA3        o367(.A(ori_ori_n380_), .B(ori_ori_n374_), .C(ori_ori_n302_), .Y(ori_ori_n390_));
  INV        o368(.A(x14), .Y(ori_ori_n391_));
  NO3        o369(.A(ori_ori_n148_), .B(ori_ori_n71_), .C(ori_ori_n53_), .Y(ori_ori_n392_));
  NO2        o370(.A(ori_ori_n392_), .B(ori_ori_n391_), .Y(ori_ori_n393_));
  NA3        o371(.A(ori_ori_n393_), .B(ori_ori_n390_), .C(ori_ori_n389_), .Y(ori_ori_n394_));
  AOI220     o372(.A0(ori_ori_n370_), .A1(ori_ori_n57_), .B0(ori_ori_n379_), .B1(ori_ori_n147_), .Y(ori_ori_n395_));
  NOi21      o373(.An(ori_ori_n246_), .B(ori_ori_n135_), .Y(ori_ori_n396_));
  NO3        o374(.A(ori_ori_n118_), .B(ori_ori_n24_), .C(x06), .Y(ori_ori_n397_));
  AOI210     o375(.A0(ori_ori_n252_), .A1(ori_ori_n203_), .B0(ori_ori_n397_), .Y(ori_ori_n398_));
  OAI210     o376(.A0(ori_ori_n44_), .A1(x04), .B0(ori_ori_n398_), .Y(ori_ori_n399_));
  OAI210     o377(.A0(ori_ori_n399_), .A1(ori_ori_n396_), .B0(ori_ori_n96_), .Y(ori_ori_n400_));
  OAI210     o378(.A0(ori_ori_n395_), .A1(ori_ori_n86_), .B0(ori_ori_n400_), .Y(ori_ori_n401_));
  NO4        o379(.A(ori_ori_n401_), .B(ori_ori_n394_), .C(ori_ori_n386_), .D(ori_ori_n372_), .Y(ori06));
  INV        o380(.A(x02), .Y(ori_ori_n405_));
  INV        o381(.A(ori_ori_n69_), .Y(ori_ori_n406_));
  INV        o382(.A(ori_ori_n40_), .Y(ori_ori_n407_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m046(.A0(mai_mai_n68_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x09), .B(x05), .Y(mai_mai_n71_));
  NA2        m049(.A(x10), .B(x06), .Y(mai_mai_n72_));
  NA3        m050(.A(mai_mai_n72_), .B(mai_mai_n71_), .C(mai_mai_n28_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n73_), .A1(x11), .B0(x03), .Y(mai_mai_n74_));
  NOi31      m052(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n75_));
  NO2        m053(.A(mai_mai_n419_), .B(mai_mai_n24_), .Y(mai_mai_n76_));
  NO2        m054(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n77_), .B(mai_mai_n36_), .Y(mai_mai_n78_));
  OAI210     m056(.A0(mai_mai_n77_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n79_));
  AOI210     m057(.A0(mai_mai_n78_), .A1(mai_mai_n48_), .B0(mai_mai_n79_), .Y(mai_mai_n80_));
  NO2        m058(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n81_));
  NO2        m059(.A(x08), .B(x01), .Y(mai_mai_n82_));
  OAI210     m060(.A0(mai_mai_n82_), .A1(mai_mai_n81_), .B0(mai_mai_n35_), .Y(mai_mai_n83_));
  NA2        m061(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n84_));
  NO3        m062(.A(mai_mai_n83_), .B(mai_mai_n80_), .C(mai_mai_n76_), .Y(mai_mai_n85_));
  AN2        m063(.A(mai_mai_n85_), .B(mai_mai_n74_), .Y(mai_mai_n86_));
  INV        m064(.A(mai_mai_n83_), .Y(mai_mai_n87_));
  NO2        m065(.A(x06), .B(x05), .Y(mai_mai_n88_));
  NA2        m066(.A(x11), .B(x00), .Y(mai_mai_n89_));
  NO2        m067(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n90_));
  NOi21      m068(.An(mai_mai_n89_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  AOI210     m069(.A0(mai_mai_n88_), .A1(mai_mai_n87_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NOi21      m070(.An(x01), .B(x10), .Y(mai_mai_n93_));
  NO2        m071(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n94_));
  NO3        m072(.A(mai_mai_n94_), .B(mai_mai_n93_), .C(x06), .Y(mai_mai_n95_));
  NA2        m073(.A(mai_mai_n95_), .B(mai_mai_n27_), .Y(mai_mai_n96_));
  OAI210     m074(.A0(mai_mai_n92_), .A1(x07), .B0(mai_mai_n96_), .Y(mai_mai_n97_));
  NO3        m075(.A(mai_mai_n97_), .B(mai_mai_n86_), .C(mai_mai_n70_), .Y(mai01));
  INV        m076(.A(x12), .Y(mai_mai_n99_));
  INV        m077(.A(x13), .Y(mai_mai_n100_));
  NA2        m078(.A(mai_mai_n93_), .B(mai_mai_n28_), .Y(mai_mai_n101_));
  NO2        m079(.A(x10), .B(x01), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NA2        m082(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n106_));
  NOi21      m084(.An(mai_mai_n106_), .B(mai_mai_n58_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n108_));
  NA3        m086(.A(x13), .B(mai_mai_n108_), .C(x06), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n109_), .B(mai_mai_n107_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n82_), .B(x13), .Y(mai_mai_n111_));
  NA2        m089(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n112_), .B(mai_mai_n111_), .Y(mai_mai_n113_));
  NA2        m091(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n114_), .B(x05), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n115_), .B(mai_mai_n113_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n117_));
  INV        m095(.A(mai_mai_n107_), .Y(mai_mai_n118_));
  AOI210     m096(.A0(mai_mai_n118_), .A1(mai_mai_n116_), .B0(mai_mai_n72_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n120_));
  NA2        m098(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n121_), .B(mai_mai_n120_), .Y(mai_mai_n122_));
  NA2        m100(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n36_), .B(x04), .Y(mai_mai_n124_));
  NA3        m102(.A(mai_mai_n124_), .B(mai_mai_n123_), .C(x13), .Y(mai_mai_n125_));
  NO3        m103(.A(mai_mai_n117_), .B(mai_mai_n77_), .C(mai_mai_n36_), .Y(mai_mai_n126_));
  NO2        m104(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n127_));
  NOi41      m105(.An(mai_mai_n125_), .B(mai_mai_n127_), .C(mai_mai_n126_), .D(mai_mai_n122_), .Y(mai_mai_n128_));
  NO3        m106(.A(mai_mai_n128_), .B(x06), .C(x03), .Y(mai_mai_n129_));
  NO3        m107(.A(mai_mai_n129_), .B(mai_mai_n119_), .C(mai_mai_n110_), .Y(mai_mai_n130_));
  NA2        m108(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n131_));
  OAI210     m109(.A0(mai_mai_n82_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n132_));
  NA2        m110(.A(mai_mai_n132_), .B(mai_mai_n131_), .Y(mai_mai_n133_));
  NO2        m111(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n134_));
  NA2        m112(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n135_));
  AOI210     m113(.A0(mai_mai_n135_), .A1(mai_mai_n49_), .B0(mai_mai_n134_), .Y(mai_mai_n136_));
  AN2        m114(.A(mai_mai_n136_), .B(mai_mai_n133_), .Y(mai_mai_n137_));
  NO2        m115(.A(x09), .B(x05), .Y(mai_mai_n138_));
  NA2        m116(.A(mai_mai_n138_), .B(mai_mai_n47_), .Y(mai_mai_n139_));
  AOI210     m117(.A0(mai_mai_n139_), .A1(mai_mai_n104_), .B0(mai_mai_n49_), .Y(mai_mai_n140_));
  NA2        m118(.A(x09), .B(x00), .Y(mai_mai_n141_));
  NA2        m119(.A(mai_mai_n106_), .B(mai_mai_n141_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n140_), .B(mai_mai_n137_), .Y(mai_mai_n143_));
  NO2        m121(.A(x03), .B(x02), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n83_), .B(mai_mai_n100_), .Y(mai_mai_n145_));
  OAI210     m123(.A0(mai_mai_n145_), .A1(mai_mai_n107_), .B0(mai_mai_n144_), .Y(mai_mai_n146_));
  OA210      m124(.A0(mai_mai_n143_), .A1(x11), .B0(mai_mai_n146_), .Y(mai_mai_n147_));
  OAI210     m125(.A0(mai_mai_n130_), .A1(mai_mai_n23_), .B0(mai_mai_n147_), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n104_), .B(mai_mai_n40_), .Y(mai_mai_n149_));
  NAi21      m127(.An(x06), .B(x10), .Y(mai_mai_n150_));
  NOi21      m128(.An(x01), .B(x13), .Y(mai_mai_n151_));
  NA2        m129(.A(mai_mai_n151_), .B(mai_mai_n150_), .Y(mai_mai_n152_));
  BUFFER     m130(.A(mai_mai_n152_), .Y(mai_mai_n153_));
  AOI210     m131(.A0(mai_mai_n153_), .A1(mai_mai_n149_), .B0(mai_mai_n41_), .Y(mai_mai_n154_));
  NO2        m132(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n100_), .B(x01), .Y(mai_mai_n156_));
  NO2        m134(.A(mai_mai_n156_), .B(x08), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n155_), .B(mai_mai_n48_), .Y(mai_mai_n158_));
  AOI210     m136(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n159_));
  OAI210     m137(.A0(mai_mai_n158_), .A1(mai_mai_n154_), .B0(mai_mai_n159_), .Y(mai_mai_n160_));
  NA2        m138(.A(x04), .B(x02), .Y(mai_mai_n161_));
  NA2        m139(.A(x10), .B(x05), .Y(mai_mai_n162_));
  NA2        m140(.A(x09), .B(x06), .Y(mai_mai_n163_));
  NO2        m141(.A(x09), .B(x01), .Y(mai_mai_n164_));
  NO2        m142(.A(mai_mai_n164_), .B(mai_mai_n31_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(x00), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n106_), .B(x08), .Y(mai_mai_n167_));
  OAI210     m145(.A0(mai_mai_n420_), .A1(x11), .B0(mai_mai_n166_), .Y(mai_mai_n168_));
  NAi21      m146(.An(mai_mai_n161_), .B(mai_mai_n168_), .Y(mai_mai_n169_));
  INV        m147(.A(mai_mai_n25_), .Y(mai_mai_n170_));
  NAi21      m148(.An(x13), .B(x00), .Y(mai_mai_n171_));
  AOI220     m149(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n172_));
  AN2        m150(.A(mai_mai_n72_), .B(mai_mai_n71_), .Y(mai_mai_n173_));
  NO2        m151(.A(mai_mai_n94_), .B(x06), .Y(mai_mai_n174_));
  NO2        m152(.A(mai_mai_n171_), .B(mai_mai_n36_), .Y(mai_mai_n175_));
  INV        m153(.A(mai_mai_n175_), .Y(mai_mai_n176_));
  OAI220     m154(.A0(mai_mai_n176_), .A1(mai_mai_n163_), .B0(mai_mai_n174_), .B1(mai_mai_n173_), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n177_), .B(mai_mai_n170_), .Y(mai_mai_n178_));
  NOi21      m156(.An(x09), .B(x00), .Y(mai_mai_n179_));
  NO3        m157(.A(mai_mai_n81_), .B(mai_mai_n179_), .C(mai_mai_n47_), .Y(mai_mai_n180_));
  NA2        m158(.A(mai_mai_n180_), .B(mai_mai_n121_), .Y(mai_mai_n181_));
  NA2        m159(.A(x10), .B(x08), .Y(mai_mai_n182_));
  INV        m160(.A(mai_mai_n182_), .Y(mai_mai_n183_));
  NA2        m161(.A(x06), .B(x05), .Y(mai_mai_n184_));
  OAI210     m162(.A0(mai_mai_n184_), .A1(mai_mai_n35_), .B0(mai_mai_n99_), .Y(mai_mai_n185_));
  AOI210     m163(.A0(mai_mai_n183_), .A1(mai_mai_n58_), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  NA2        m164(.A(mai_mai_n186_), .B(mai_mai_n181_), .Y(mai_mai_n187_));
  NO2        m165(.A(mai_mai_n100_), .B(x12), .Y(mai_mai_n188_));
  AOI210     m166(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n188_), .Y(mai_mai_n189_));
  NO2        m167(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n190_));
  NA2        m168(.A(mai_mai_n190_), .B(x02), .Y(mai_mai_n191_));
  NA2        m169(.A(mai_mai_n189_), .B(mai_mai_n187_), .Y(mai_mai_n192_));
  NA4        m170(.A(mai_mai_n192_), .B(mai_mai_n178_), .C(mai_mai_n169_), .D(mai_mai_n160_), .Y(mai_mai_n193_));
  AOI210     m171(.A0(mai_mai_n148_), .A1(mai_mai_n99_), .B0(mai_mai_n193_), .Y(mai_mai_n194_));
  INV        m172(.A(mai_mai_n73_), .Y(mai_mai_n195_));
  NA2        m173(.A(mai_mai_n195_), .B(mai_mai_n133_), .Y(mai_mai_n196_));
  NA2        m174(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n197_));
  NA2        m175(.A(mai_mai_n197_), .B(mai_mai_n132_), .Y(mai_mai_n198_));
  AOI210     m176(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n199_));
  NO2        m177(.A(mai_mai_n120_), .B(x06), .Y(mai_mai_n200_));
  AOI210     m178(.A0(mai_mai_n199_), .A1(mai_mai_n198_), .B0(mai_mai_n200_), .Y(mai_mai_n201_));
  AOI210     m179(.A0(mai_mai_n201_), .A1(mai_mai_n196_), .B0(x12), .Y(mai_mai_n202_));
  INV        m180(.A(mai_mai_n75_), .Y(mai_mai_n203_));
  NO2        m181(.A(x05), .B(mai_mai_n51_), .Y(mai_mai_n204_));
  OAI210     m182(.A0(mai_mai_n204_), .A1(mai_mai_n152_), .B0(mai_mai_n57_), .Y(mai_mai_n205_));
  NA2        m183(.A(mai_mai_n205_), .B(mai_mai_n203_), .Y(mai_mai_n206_));
  NO2        m184(.A(mai_mai_n93_), .B(x06), .Y(mai_mai_n207_));
  AOI210     m185(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n208_));
  NO3        m186(.A(mai_mai_n208_), .B(mai_mai_n207_), .C(mai_mai_n41_), .Y(mai_mai_n209_));
  NA4        m187(.A(mai_mai_n150_), .B(mai_mai_n56_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n210_));
  NA2        m188(.A(mai_mai_n210_), .B(mai_mai_n135_), .Y(mai_mai_n211_));
  OAI210     m189(.A0(mai_mai_n211_), .A1(mai_mai_n209_), .B0(x02), .Y(mai_mai_n212_));
  AOI210     m190(.A0(mai_mai_n212_), .A1(mai_mai_n206_), .B0(mai_mai_n23_), .Y(mai_mai_n213_));
  OAI210     m191(.A0(mai_mai_n202_), .A1(mai_mai_n57_), .B0(mai_mai_n213_), .Y(mai_mai_n214_));
  INV        m192(.A(mai_mai_n135_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n216_));
  OAI210     m194(.A0(mai_mai_n77_), .A1(mai_mai_n36_), .B0(mai_mai_n112_), .Y(mai_mai_n217_));
  NO2        m195(.A(mai_mai_n100_), .B(x03), .Y(mai_mai_n218_));
  AOI220     m196(.A0(mai_mai_n218_), .A1(mai_mai_n217_), .B0(mai_mai_n75_), .B1(mai_mai_n216_), .Y(mai_mai_n219_));
  NA2        m197(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n220_));
  INV        m198(.A(mai_mai_n150_), .Y(mai_mai_n221_));
  NOi21      m199(.An(x13), .B(x04), .Y(mai_mai_n222_));
  NO3        m200(.A(mai_mai_n222_), .B(mai_mai_n75_), .C(mai_mai_n179_), .Y(mai_mai_n223_));
  NO2        m201(.A(mai_mai_n223_), .B(x05), .Y(mai_mai_n224_));
  AOI220     m202(.A0(mai_mai_n224_), .A1(mai_mai_n220_), .B0(mai_mai_n221_), .B1(mai_mai_n57_), .Y(mai_mai_n225_));
  OAI210     m203(.A0(mai_mai_n219_), .A1(mai_mai_n215_), .B0(mai_mai_n225_), .Y(mai_mai_n226_));
  INV        m204(.A(mai_mai_n90_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n227_), .B(x12), .Y(mai_mai_n228_));
  NA2        m206(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n229_));
  NO2        m207(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n230_));
  AOI210     m208(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n231_));
  NO2        m209(.A(x06), .B(x00), .Y(mai_mai_n232_));
  NO3        m210(.A(mai_mai_n232_), .B(mai_mai_n231_), .C(mai_mai_n41_), .Y(mai_mai_n233_));
  INV        m211(.A(mai_mai_n72_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n234_), .B(mai_mai_n233_), .Y(mai_mai_n235_));
  NA2        m213(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n236_));
  NA2        m214(.A(mai_mai_n236_), .B(x03), .Y(mai_mai_n237_));
  OR2        m215(.A(mai_mai_n237_), .B(mai_mai_n235_), .Y(mai_mai_n238_));
  NA2        m216(.A(x13), .B(mai_mai_n99_), .Y(mai_mai_n239_));
  NA3        m217(.A(mai_mai_n239_), .B(mai_mai_n185_), .C(mai_mai_n91_), .Y(mai_mai_n240_));
  OAI210     m218(.A0(mai_mai_n238_), .A1(mai_mai_n229_), .B0(mai_mai_n240_), .Y(mai_mai_n241_));
  AOI210     m219(.A0(mai_mai_n228_), .A1(mai_mai_n226_), .B0(mai_mai_n241_), .Y(mai_mai_n242_));
  AOI210     m220(.A0(mai_mai_n242_), .A1(mai_mai_n214_), .B0(x07), .Y(mai_mai_n243_));
  NA2        m221(.A(mai_mai_n71_), .B(mai_mai_n29_), .Y(mai_mai_n244_));
  NOi31      m222(.An(mai_mai_n131_), .B(mai_mai_n222_), .C(mai_mai_n179_), .Y(mai_mai_n245_));
  NO2        m223(.A(mai_mai_n245_), .B(mai_mai_n244_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n100_), .B(x06), .Y(mai_mai_n247_));
  INV        m225(.A(mai_mai_n247_), .Y(mai_mai_n248_));
  NO2        m226(.A(x08), .B(x05), .Y(mai_mai_n249_));
  NO2        m227(.A(mai_mai_n249_), .B(mai_mai_n231_), .Y(mai_mai_n250_));
  OAI210     m228(.A0(mai_mai_n75_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n251_));
  OAI210     m229(.A0(mai_mai_n250_), .A1(mai_mai_n248_), .B0(mai_mai_n251_), .Y(mai_mai_n252_));
  NO2        m230(.A(x12), .B(x02), .Y(mai_mai_n253_));
  INV        m231(.A(mai_mai_n253_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n254_), .B(mai_mai_n227_), .Y(mai_mai_n255_));
  OA210      m233(.A0(mai_mai_n252_), .A1(mai_mai_n246_), .B0(mai_mai_n255_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n257_));
  NO2        m235(.A(mai_mai_n257_), .B(x01), .Y(mai_mai_n258_));
  NO2        m236(.A(mai_mai_n125_), .B(mai_mai_n29_), .Y(mai_mai_n259_));
  NA2        m237(.A(mai_mai_n247_), .B(mai_mai_n217_), .Y(mai_mai_n260_));
  NA2        m238(.A(mai_mai_n100_), .B(x04), .Y(mai_mai_n261_));
  NA2        m239(.A(mai_mai_n261_), .B(mai_mai_n28_), .Y(mai_mai_n262_));
  OAI210     m240(.A0(mai_mai_n262_), .A1(mai_mai_n111_), .B0(mai_mai_n260_), .Y(mai_mai_n263_));
  NO3        m241(.A(mai_mai_n89_), .B(x12), .C(x03), .Y(mai_mai_n264_));
  OAI210     m242(.A0(mai_mai_n263_), .A1(mai_mai_n259_), .B0(mai_mai_n264_), .Y(mai_mai_n265_));
  NOi21      m243(.An(mai_mai_n244_), .B(mai_mai_n207_), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n267_));
  NA2        m245(.A(mai_mai_n266_), .B(mai_mai_n267_), .Y(mai_mai_n268_));
  NO2        m246(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n269_));
  NO3        m247(.A(mai_mai_n269_), .B(mai_mai_n208_), .C(mai_mai_n174_), .Y(mai_mai_n270_));
  NO2        m248(.A(mai_mai_n229_), .B(mai_mai_n28_), .Y(mai_mai_n271_));
  OAI210     m249(.A0(mai_mai_n270_), .A1(mai_mai_n215_), .B0(mai_mai_n271_), .Y(mai_mai_n272_));
  NA3        m250(.A(mai_mai_n272_), .B(mai_mai_n268_), .C(mai_mai_n265_), .Y(mai_mai_n273_));
  NO3        m251(.A(mai_mai_n273_), .B(mai_mai_n256_), .C(mai_mai_n243_), .Y(mai_mai_n274_));
  OAI210     m252(.A0(mai_mai_n194_), .A1(mai_mai_n61_), .B0(mai_mai_n274_), .Y(mai02));
  AOI210     m253(.A0(mai_mai_n131_), .A1(mai_mai_n83_), .B0(mai_mai_n123_), .Y(mai_mai_n276_));
  NOi21      m254(.An(mai_mai_n223_), .B(mai_mai_n164_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n100_), .B(mai_mai_n35_), .Y(mai_mai_n278_));
  NA3        m256(.A(mai_mai_n278_), .B(mai_mai_n183_), .C(mai_mai_n56_), .Y(mai_mai_n279_));
  OAI210     m257(.A0(mai_mai_n277_), .A1(mai_mai_n32_), .B0(mai_mai_n279_), .Y(mai_mai_n280_));
  OAI210     m258(.A0(mai_mai_n280_), .A1(mai_mai_n276_), .B0(mai_mai_n162_), .Y(mai_mai_n281_));
  INV        m259(.A(mai_mai_n162_), .Y(mai_mai_n282_));
  AOI210     m260(.A0(mai_mai_n108_), .A1(mai_mai_n84_), .B0(mai_mai_n208_), .Y(mai_mai_n283_));
  NO2        m261(.A(mai_mai_n283_), .B(mai_mai_n100_), .Y(mai_mai_n284_));
  AOI220     m262(.A0(mai_mai_n284_), .A1(mai_mai_n282_), .B0(mai_mai_n145_), .B1(mai_mai_n144_), .Y(mai_mai_n285_));
  AOI210     m263(.A0(mai_mai_n285_), .A1(mai_mai_n281_), .B0(mai_mai_n48_), .Y(mai_mai_n286_));
  NO2        m264(.A(x05), .B(x02), .Y(mai_mai_n287_));
  OAI210     m265(.A0(mai_mai_n198_), .A1(mai_mai_n179_), .B0(mai_mai_n287_), .Y(mai_mai_n288_));
  AOI220     m266(.A0(mai_mai_n249_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n289_));
  NOi21      m267(.An(mai_mai_n278_), .B(mai_mai_n289_), .Y(mai_mai_n290_));
  AOI210     m268(.A0(mai_mai_n222_), .A1(mai_mai_n77_), .B0(mai_mai_n290_), .Y(mai_mai_n291_));
  AOI210     m269(.A0(mai_mai_n291_), .A1(mai_mai_n288_), .B0(mai_mai_n135_), .Y(mai_mai_n292_));
  NAi21      m270(.An(mai_mai_n224_), .B(mai_mai_n219_), .Y(mai_mai_n293_));
  NO2        m271(.A(mai_mai_n236_), .B(mai_mai_n47_), .Y(mai_mai_n294_));
  NA2        m272(.A(mai_mai_n294_), .B(mai_mai_n293_), .Y(mai_mai_n295_));
  AN2        m273(.A(mai_mai_n218_), .B(mai_mai_n217_), .Y(mai_mai_n296_));
  OAI210     m274(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n297_));
  NA2        m275(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n298_));
  OA210      m276(.A0(mai_mai_n298_), .A1(x08), .B0(mai_mai_n139_), .Y(mai_mai_n299_));
  AOI210     m277(.A0(mai_mai_n299_), .A1(mai_mai_n132_), .B0(mai_mai_n297_), .Y(mai_mai_n300_));
  OAI210     m278(.A0(mai_mai_n300_), .A1(mai_mai_n296_), .B0(mai_mai_n94_), .Y(mai_mai_n301_));
  INV        m279(.A(mai_mai_n144_), .Y(mai_mai_n302_));
  OAI220     m280(.A0(mai_mai_n250_), .A1(mai_mai_n101_), .B0(mai_mai_n302_), .B1(mai_mai_n122_), .Y(mai_mai_n303_));
  NA2        m281(.A(mai_mai_n303_), .B(x13), .Y(mai_mai_n304_));
  NA3        m282(.A(mai_mai_n304_), .B(mai_mai_n301_), .C(mai_mai_n295_), .Y(mai_mai_n305_));
  NO3        m283(.A(mai_mai_n305_), .B(mai_mai_n292_), .C(mai_mai_n286_), .Y(mai_mai_n306_));
  NA2        m284(.A(mai_mai_n134_), .B(x03), .Y(mai_mai_n307_));
  OAI210     m285(.A0(mai_mai_n171_), .A1(mai_mai_n269_), .B0(mai_mai_n307_), .Y(mai_mai_n308_));
  NA2        m286(.A(mai_mai_n308_), .B(mai_mai_n102_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n161_), .B(mai_mai_n156_), .Y(mai_mai_n310_));
  AN2        m288(.A(mai_mai_n310_), .B(mai_mai_n167_), .Y(mai_mai_n311_));
  INV        m289(.A(mai_mai_n56_), .Y(mai_mai_n312_));
  OAI220     m290(.A0(mai_mai_n261_), .A1(mai_mai_n312_), .B0(mai_mai_n123_), .B1(mai_mai_n28_), .Y(mai_mai_n313_));
  OAI210     m291(.A0(mai_mai_n313_), .A1(mai_mai_n311_), .B0(mai_mai_n103_), .Y(mai_mai_n314_));
  NA2        m292(.A(mai_mai_n261_), .B(mai_mai_n99_), .Y(mai_mai_n315_));
  NA2        m293(.A(mai_mai_n99_), .B(mai_mai_n41_), .Y(mai_mai_n316_));
  NA3        m294(.A(mai_mai_n316_), .B(mai_mai_n315_), .C(mai_mai_n122_), .Y(mai_mai_n317_));
  NA4        m295(.A(mai_mai_n317_), .B(mai_mai_n314_), .C(mai_mai_n309_), .D(mai_mai_n48_), .Y(mai_mai_n318_));
  INV        m296(.A(mai_mai_n190_), .Y(mai_mai_n319_));
  NO2        m297(.A(mai_mai_n157_), .B(mai_mai_n40_), .Y(mai_mai_n320_));
  NA2        m298(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n321_));
  OAI220     m299(.A0(mai_mai_n321_), .A1(mai_mai_n320_), .B0(mai_mai_n319_), .B1(mai_mai_n59_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n322_), .B(x02), .Y(mai_mai_n323_));
  INV        m301(.A(mai_mai_n230_), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n188_), .B(x04), .Y(mai_mai_n325_));
  NO2        m303(.A(mai_mai_n325_), .B(mai_mai_n324_), .Y(mai_mai_n326_));
  NO3        m304(.A(mai_mai_n172_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n327_));
  OAI210     m305(.A0(mai_mai_n327_), .A1(mai_mai_n326_), .B0(mai_mai_n94_), .Y(mai_mai_n328_));
  NO3        m306(.A(mai_mai_n188_), .B(mai_mai_n155_), .C(mai_mai_n52_), .Y(mai_mai_n329_));
  OAI210     m307(.A0(mai_mai_n141_), .A1(mai_mai_n36_), .B0(mai_mai_n99_), .Y(mai_mai_n330_));
  OAI210     m308(.A0(mai_mai_n330_), .A1(mai_mai_n180_), .B0(mai_mai_n329_), .Y(mai_mai_n331_));
  NA4        m309(.A(mai_mai_n331_), .B(mai_mai_n328_), .C(mai_mai_n323_), .D(x06), .Y(mai_mai_n332_));
  NA2        m310(.A(x09), .B(x03), .Y(mai_mai_n333_));
  OAI220     m311(.A0(mai_mai_n333_), .A1(mai_mai_n121_), .B0(mai_mai_n197_), .B1(mai_mai_n64_), .Y(mai_mai_n334_));
  OAI220     m312(.A0(mai_mai_n156_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n335_));
  NO3        m313(.A(mai_mai_n269_), .B(mai_mai_n120_), .C(x08), .Y(mai_mai_n336_));
  AOI210     m314(.A0(mai_mai_n335_), .A1(mai_mai_n215_), .B0(mai_mai_n336_), .Y(mai_mai_n337_));
  NO2        m315(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n338_));
  NA2        m316(.A(mai_mai_n329_), .B(mai_mai_n338_), .Y(mai_mai_n339_));
  OAI210     m317(.A0(mai_mai_n337_), .A1(mai_mai_n28_), .B0(mai_mai_n339_), .Y(mai_mai_n340_));
  AO220      m318(.A0(mai_mai_n340_), .A1(x04), .B0(mai_mai_n334_), .B1(x05), .Y(mai_mai_n341_));
  AOI210     m319(.A0(mai_mai_n332_), .A1(mai_mai_n318_), .B0(mai_mai_n341_), .Y(mai_mai_n342_));
  OAI210     m320(.A0(mai_mai_n306_), .A1(x12), .B0(mai_mai_n342_), .Y(mai03));
  OR2        m321(.A(mai_mai_n42_), .B(mai_mai_n216_), .Y(mai_mai_n344_));
  AOI210     m322(.A0(mai_mai_n145_), .A1(mai_mai_n99_), .B0(mai_mai_n344_), .Y(mai_mai_n345_));
  AO210      m323(.A0(mai_mai_n324_), .A1(mai_mai_n84_), .B0(mai_mai_n325_), .Y(mai_mai_n346_));
  NA2        m324(.A(mai_mai_n188_), .B(mai_mai_n144_), .Y(mai_mai_n347_));
  NA3        m325(.A(mai_mai_n347_), .B(mai_mai_n346_), .C(mai_mai_n191_), .Y(mai_mai_n348_));
  OAI210     m326(.A0(mai_mai_n348_), .A1(mai_mai_n345_), .B0(x05), .Y(mai_mai_n349_));
  NA2        m327(.A(mai_mai_n344_), .B(x05), .Y(mai_mai_n350_));
  AOI210     m328(.A0(mai_mai_n132_), .A1(mai_mai_n203_), .B0(mai_mai_n350_), .Y(mai_mai_n351_));
  AOI210     m329(.A0(mai_mai_n218_), .A1(mai_mai_n78_), .B0(mai_mai_n115_), .Y(mai_mai_n352_));
  OAI220     m330(.A0(mai_mai_n352_), .A1(mai_mai_n59_), .B0(mai_mai_n298_), .B1(mai_mai_n289_), .Y(mai_mai_n353_));
  OAI210     m331(.A0(mai_mai_n353_), .A1(mai_mai_n351_), .B0(mai_mai_n99_), .Y(mai_mai_n354_));
  AOI210     m332(.A0(mai_mai_n139_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n355_));
  NO2        m333(.A(mai_mai_n164_), .B(mai_mai_n127_), .Y(mai_mai_n356_));
  OAI220     m334(.A0(mai_mai_n356_), .A1(mai_mai_n37_), .B0(mai_mai_n142_), .B1(x13), .Y(mai_mai_n357_));
  OAI210     m335(.A0(mai_mai_n357_), .A1(mai_mai_n355_), .B0(x04), .Y(mai_mai_n358_));
  NO3        m336(.A(mai_mai_n316_), .B(mai_mai_n83_), .C(mai_mai_n59_), .Y(mai_mai_n359_));
  AOI210     m337(.A0(mai_mai_n176_), .A1(mai_mai_n99_), .B0(mai_mai_n139_), .Y(mai_mai_n360_));
  OA210      m338(.A0(mai_mai_n157_), .A1(x12), .B0(mai_mai_n127_), .Y(mai_mai_n361_));
  NO3        m339(.A(mai_mai_n361_), .B(mai_mai_n360_), .C(mai_mai_n359_), .Y(mai_mai_n362_));
  NA4        m340(.A(mai_mai_n362_), .B(mai_mai_n358_), .C(mai_mai_n354_), .D(mai_mai_n349_), .Y(mai04));
  NO2        m341(.A(mai_mai_n87_), .B(mai_mai_n39_), .Y(mai_mai_n364_));
  XO2        m342(.A(mai_mai_n364_), .B(mai_mai_n239_), .Y(mai05));
  NO2        m343(.A(mai_mai_n52_), .B(mai_mai_n200_), .Y(mai_mai_n366_));
  AOI210     m344(.A0(mai_mai_n366_), .A1(mai_mai_n297_), .B0(mai_mai_n25_), .Y(mai_mai_n367_));
  NO2        m345(.A(x06), .B(mai_mai_n24_), .Y(mai_mai_n368_));
  OAI210     m346(.A0(mai_mai_n368_), .A1(mai_mai_n367_), .B0(mai_mai_n99_), .Y(mai_mai_n369_));
  OAI210     m347(.A0(mai_mai_n26_), .A1(mai_mai_n99_), .B0(x07), .Y(mai_mai_n370_));
  INV        m348(.A(mai_mai_n370_), .Y(mai_mai_n371_));
  NA2        m349(.A(mai_mai_n151_), .B(x05), .Y(mai_mai_n372_));
  NA3        m350(.A(mai_mai_n372_), .B(mai_mai_n232_), .C(mai_mai_n227_), .Y(mai_mai_n373_));
  NO2        m351(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n374_));
  OR3        m352(.A(x06), .B(mai_mai_n374_), .C(mai_mai_n44_), .Y(mai_mai_n375_));
  NA3        m353(.A(mai_mai_n375_), .B(mai_mai_n373_), .C(mai_mai_n229_), .Y(mai_mai_n376_));
  NA2        m354(.A(mai_mai_n376_), .B(mai_mai_n99_), .Y(mai_mai_n377_));
  NA2        m355(.A(mai_mai_n33_), .B(mai_mai_n99_), .Y(mai_mai_n378_));
  AOI210     m356(.A0(mai_mai_n378_), .A1(mai_mai_n90_), .B0(x07), .Y(mai_mai_n379_));
  AOI220     m357(.A0(mai_mai_n379_), .A1(mai_mai_n377_), .B0(mai_mai_n371_), .B1(mai_mai_n369_), .Y(mai_mai_n380_));
  OR2        m358(.A(mai_mai_n257_), .B(mai_mai_n254_), .Y(mai_mai_n381_));
  NO2        m359(.A(x07), .B(mai_mai_n134_), .Y(mai_mai_n382_));
  OR2        m360(.A(mai_mai_n382_), .B(x03), .Y(mai_mai_n383_));
  NO2        m361(.A(x07), .B(x11), .Y(mai_mai_n384_));
  NO3        m362(.A(mai_mai_n384_), .B(mai_mai_n138_), .C(mai_mai_n28_), .Y(mai_mai_n385_));
  AOI220     m363(.A0(mai_mai_n385_), .A1(mai_mai_n383_), .B0(mai_mai_n381_), .B1(mai_mai_n47_), .Y(mai_mai_n386_));
  NA2        m364(.A(mai_mai_n386_), .B(mai_mai_n100_), .Y(mai_mai_n387_));
  AOI210     m365(.A0(mai_mai_n325_), .A1(mai_mai_n105_), .B0(mai_mai_n253_), .Y(mai_mai_n388_));
  NOi21      m366(.An(mai_mai_n307_), .B(mai_mai_n127_), .Y(mai_mai_n389_));
  NO2        m367(.A(mai_mai_n389_), .B(mai_mai_n254_), .Y(mai_mai_n390_));
  OAI210     m368(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n391_));
  AOI210     m369(.A0(mai_mai_n239_), .A1(mai_mai_n47_), .B0(mai_mai_n391_), .Y(mai_mai_n392_));
  NO4        m370(.A(mai_mai_n392_), .B(mai_mai_n390_), .C(mai_mai_n388_), .D(x08), .Y(mai_mai_n393_));
  NO2        m371(.A(x05), .B(x03), .Y(mai_mai_n394_));
  NO2        m372(.A(x13), .B(x12), .Y(mai_mai_n395_));
  NO2        m373(.A(mai_mai_n123_), .B(mai_mai_n28_), .Y(mai_mai_n396_));
  NO2        m374(.A(mai_mai_n396_), .B(mai_mai_n258_), .Y(mai_mai_n397_));
  NA3        m375(.A(mai_mai_n319_), .B(mai_mai_n117_), .C(x12), .Y(mai_mai_n398_));
  AO210      m376(.A0(mai_mai_n319_), .A1(mai_mai_n117_), .B0(mai_mai_n239_), .Y(mai_mai_n399_));
  NA3        m377(.A(mai_mai_n399_), .B(mai_mai_n398_), .C(x08), .Y(mai_mai_n400_));
  AOI210     m378(.A0(mai_mai_n395_), .A1(mai_mai_n394_), .B0(mai_mai_n400_), .Y(mai_mai_n401_));
  AOI210     m379(.A0(mai_mai_n393_), .A1(mai_mai_n387_), .B0(mai_mai_n401_), .Y(mai_mai_n402_));
  OAI210     m380(.A0(x07), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n403_));
  OAI220     m381(.A0(mai_mai_n162_), .A1(x02), .B0(mai_mai_n138_), .B1(mai_mai_n43_), .Y(mai_mai_n404_));
  OAI210     m382(.A0(mai_mai_n404_), .A1(mai_mai_n403_), .B0(mai_mai_n175_), .Y(mai_mai_n405_));
  NA3        m383(.A(mai_mai_n397_), .B(mai_mai_n389_), .C(mai_mai_n315_), .Y(mai_mai_n406_));
  INV        m384(.A(x14), .Y(mai_mai_n407_));
  NO3        m385(.A(mai_mai_n307_), .B(mai_mai_n101_), .C(x11), .Y(mai_mai_n408_));
  NO2        m386(.A(mai_mai_n408_), .B(mai_mai_n407_), .Y(mai_mai_n409_));
  NA3        m387(.A(mai_mai_n409_), .B(mai_mai_n406_), .C(mai_mai_n405_), .Y(mai_mai_n410_));
  NA2        m388(.A(mai_mai_n378_), .B(mai_mai_n61_), .Y(mai_mai_n411_));
  NOi21      m389(.An(mai_mai_n261_), .B(mai_mai_n142_), .Y(mai_mai_n412_));
  NO2        m390(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n413_));
  OAI210     m391(.A0(mai_mai_n413_), .A1(mai_mai_n412_), .B0(mai_mai_n99_), .Y(mai_mai_n414_));
  OAI210     m392(.A0(mai_mai_n411_), .A1(mai_mai_n89_), .B0(mai_mai_n414_), .Y(mai_mai_n415_));
  NO4        m393(.A(mai_mai_n415_), .B(mai_mai_n410_), .C(mai_mai_n402_), .D(mai_mai_n380_), .Y(mai06));
  INV        m394(.A(x07), .Y(mai_mai_n419_));
  INV        m395(.A(x01), .Y(mai_mai_n420_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  INV        u039(.A(men_men_n59_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n29_), .B(x02), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n24_), .Y(men_men_n64_));
  NO2        u042(.A(men_men_n64_), .B(men_men_n62_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n30_), .A1(x11), .B0(men_men_n66_), .Y(men_men_n67_));
  AOI220     u045(.A0(men_men_n67_), .A1(men_men_n59_), .B0(men_men_n65_), .B1(men_men_n31_), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n68_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x09), .Y(men_men_n70_));
  NO2        u048(.A(men_men_n61_), .B(men_men_n23_), .Y(men_men_n71_));
  NA2        u049(.A(x09), .B(x05), .Y(men_men_n72_));
  NA2        u050(.A(x10), .B(x06), .Y(men_men_n73_));
  NA2        u051(.A(men_men_n73_), .B(men_men_n72_), .Y(men_men_n74_));
  NO2        u052(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n75_));
  OAI210     u053(.A0(men_men_n74_), .A1(men_men_n71_), .B0(x03), .Y(men_men_n76_));
  NOi31      u054(.An(x08), .B(x04), .C(x00), .Y(men_men_n77_));
  NO2        u055(.A(x10), .B(x09), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n441_), .B(men_men_n24_), .Y(men_men_n79_));
  NO2        u057(.A(x09), .B(men_men_n41_), .Y(men_men_n80_));
  NO2        u058(.A(men_men_n80_), .B(men_men_n36_), .Y(men_men_n81_));
  OAI210     u059(.A0(men_men_n80_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n82_));
  AOI210     u060(.A0(men_men_n81_), .A1(men_men_n48_), .B0(men_men_n82_), .Y(men_men_n83_));
  NO2        u061(.A(men_men_n36_), .B(x00), .Y(men_men_n84_));
  NO2        u062(.A(x08), .B(x01), .Y(men_men_n85_));
  OAI210     u063(.A0(men_men_n85_), .A1(men_men_n84_), .B0(men_men_n35_), .Y(men_men_n86_));
  NA2        u064(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n87_));
  NO3        u065(.A(men_men_n86_), .B(men_men_n83_), .C(men_men_n79_), .Y(men_men_n88_));
  AN2        u066(.A(men_men_n88_), .B(men_men_n76_), .Y(men_men_n89_));
  INV        u067(.A(men_men_n86_), .Y(men_men_n90_));
  NO2        u068(.A(x06), .B(x05), .Y(men_men_n91_));
  NA2        u069(.A(x11), .B(x00), .Y(men_men_n92_));
  NO2        u070(.A(x11), .B(men_men_n47_), .Y(men_men_n93_));
  NOi21      u071(.An(men_men_n92_), .B(men_men_n93_), .Y(men_men_n94_));
  NOi21      u072(.An(x01), .B(x10), .Y(men_men_n95_));
  NO2        u073(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n96_));
  NO3        u074(.A(men_men_n96_), .B(men_men_n95_), .C(x06), .Y(men_men_n97_));
  NA2        u075(.A(men_men_n97_), .B(men_men_n27_), .Y(men_men_n98_));
  OAI210     u076(.A0(men_men_n444_), .A1(x07), .B0(men_men_n98_), .Y(men_men_n99_));
  NO3        u077(.A(men_men_n99_), .B(men_men_n89_), .C(men_men_n69_), .Y(men01));
  INV        u078(.A(x12), .Y(men_men_n101_));
  INV        u079(.A(x13), .Y(men_men_n102_));
  NA2        u080(.A(men_men_n446_), .B(men_men_n70_), .Y(men_men_n103_));
  NA2        u081(.A(x08), .B(x04), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n104_), .B(men_men_n57_), .Y(men_men_n105_));
  NA2        u083(.A(men_men_n105_), .B(men_men_n103_), .Y(men_men_n106_));
  NA2        u084(.A(men_men_n95_), .B(men_men_n28_), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n107_), .B(men_men_n72_), .Y(men_men_n108_));
  NO2        u086(.A(x10), .B(x01), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n29_), .B(x00), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n110_), .B(men_men_n109_), .Y(men_men_n111_));
  NA2        u089(.A(x04), .B(men_men_n28_), .Y(men_men_n112_));
  NO3        u090(.A(men_men_n112_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n113_));
  AOI210     u091(.A0(men_men_n113_), .A1(men_men_n111_), .B0(men_men_n108_), .Y(men_men_n114_));
  AOI210     u092(.A0(men_men_n114_), .A1(men_men_n106_), .B0(men_men_n102_), .Y(men_men_n115_));
  NO2        u093(.A(men_men_n56_), .B(x05), .Y(men_men_n116_));
  NOi21      u094(.An(men_men_n116_), .B(men_men_n58_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n35_), .B(x02), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n102_), .B(men_men_n36_), .Y(men_men_n119_));
  NA3        u097(.A(men_men_n119_), .B(men_men_n118_), .C(x06), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n120_), .B(men_men_n117_), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n85_), .B(x13), .Y(men_men_n122_));
  NA2        u100(.A(x09), .B(men_men_n35_), .Y(men_men_n123_));
  NA2        u101(.A(x13), .B(men_men_n35_), .Y(men_men_n124_));
  NO2        u102(.A(men_men_n124_), .B(x05), .Y(men_men_n125_));
  NA2        u103(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n126_));
  NO2        u104(.A(x00), .B(men_men_n73_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n128_));
  NA2        u106(.A(x10), .B(men_men_n57_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n129_), .B(men_men_n128_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n51_), .B(x05), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n131_), .B(x13), .Y(men_men_n132_));
  NO3        u110(.A(men_men_n126_), .B(men_men_n80_), .C(men_men_n36_), .Y(men_men_n133_));
  NO2        u111(.A(men_men_n60_), .B(x05), .Y(men_men_n134_));
  NOi41      u112(.An(men_men_n132_), .B(men_men_n134_), .C(men_men_n133_), .D(men_men_n130_), .Y(men_men_n135_));
  NO3        u113(.A(men_men_n135_), .B(x06), .C(x03), .Y(men_men_n136_));
  NO4        u114(.A(men_men_n136_), .B(men_men_n127_), .C(men_men_n121_), .D(men_men_n115_), .Y(men_men_n137_));
  NA2        u115(.A(x13), .B(men_men_n36_), .Y(men_men_n138_));
  OAI210     u116(.A0(men_men_n85_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  NO2        u118(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n141_));
  OA210      u119(.A0(x00), .A1(men_men_n78_), .B0(men_men_n141_), .Y(men_men_n142_));
  NO2        u120(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n29_), .B(x06), .Y(men_men_n144_));
  AOI210     u122(.A0(men_men_n144_), .A1(men_men_n49_), .B0(men_men_n143_), .Y(men_men_n145_));
  OA210      u123(.A0(men_men_n145_), .A1(men_men_n142_), .B0(men_men_n140_), .Y(men_men_n146_));
  NO2        u124(.A(x09), .B(x05), .Y(men_men_n147_));
  NA2        u125(.A(men_men_n147_), .B(men_men_n47_), .Y(men_men_n148_));
  AOI210     u126(.A0(men_men_n148_), .A1(men_men_n111_), .B0(men_men_n49_), .Y(men_men_n149_));
  NA2        u127(.A(x09), .B(x00), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n116_), .B(men_men_n150_), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n77_), .B(men_men_n51_), .Y(men_men_n152_));
  AOI210     u130(.A0(men_men_n152_), .A1(men_men_n151_), .B0(men_men_n144_), .Y(men_men_n153_));
  NO3        u131(.A(men_men_n153_), .B(men_men_n149_), .C(men_men_n146_), .Y(men_men_n154_));
  NO2        u132(.A(x03), .B(x02), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n86_), .B(men_men_n102_), .Y(men_men_n156_));
  OAI210     u134(.A0(men_men_n156_), .A1(men_men_n117_), .B0(men_men_n155_), .Y(men_men_n157_));
  OA210      u135(.A0(men_men_n154_), .A1(x11), .B0(men_men_n157_), .Y(men_men_n158_));
  OAI210     u136(.A0(men_men_n137_), .A1(men_men_n23_), .B0(men_men_n158_), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n111_), .B(men_men_n40_), .Y(men_men_n160_));
  NAi21      u138(.An(x06), .B(x10), .Y(men_men_n161_));
  NOi21      u139(.An(x01), .B(x13), .Y(men_men_n162_));
  NA2        u140(.A(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  OR2        u141(.A(men_men_n163_), .B(x08), .Y(men_men_n164_));
  AOI210     u142(.A0(men_men_n164_), .A1(men_men_n160_), .B0(men_men_n41_), .Y(men_men_n165_));
  NO2        u143(.A(men_men_n29_), .B(x03), .Y(men_men_n166_));
  NA2        u144(.A(men_men_n102_), .B(x01), .Y(men_men_n167_));
  NO2        u145(.A(men_men_n167_), .B(x08), .Y(men_men_n168_));
  OAI210     u146(.A0(x05), .A1(men_men_n168_), .B0(men_men_n51_), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n169_), .A1(men_men_n166_), .B0(men_men_n48_), .Y(men_men_n170_));
  AOI210     u148(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n171_));
  OAI210     u149(.A0(men_men_n170_), .A1(men_men_n165_), .B0(men_men_n171_), .Y(men_men_n172_));
  NA2        u150(.A(x04), .B(x02), .Y(men_men_n173_));
  NA2        u151(.A(x10), .B(x05), .Y(men_men_n174_));
  NO2        u152(.A(x09), .B(x01), .Y(men_men_n175_));
  NO2        u153(.A(men_men_n109_), .B(men_men_n31_), .Y(men_men_n176_));
  NA2        u154(.A(men_men_n176_), .B(x00), .Y(men_men_n177_));
  NO2        u155(.A(men_men_n116_), .B(x08), .Y(men_men_n178_));
  NA3        u156(.A(men_men_n162_), .B(men_men_n161_), .C(men_men_n51_), .Y(men_men_n179_));
  NA2        u157(.A(men_men_n95_), .B(x05), .Y(men_men_n180_));
  OAI210     u158(.A0(men_men_n180_), .A1(men_men_n119_), .B0(men_men_n179_), .Y(men_men_n181_));
  AOI210     u159(.A0(men_men_n178_), .A1(x06), .B0(men_men_n181_), .Y(men_men_n182_));
  OAI210     u160(.A0(men_men_n182_), .A1(x11), .B0(men_men_n177_), .Y(men_men_n183_));
  NAi21      u161(.An(men_men_n173_), .B(men_men_n183_), .Y(men_men_n184_));
  INV        u162(.A(men_men_n25_), .Y(men_men_n185_));
  NAi21      u163(.An(x13), .B(x00), .Y(men_men_n186_));
  AOI210     u164(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n186_), .Y(men_men_n187_));
  BUFFER     u165(.A(men_men_n187_), .Y(men_men_n188_));
  BUFFER     u166(.A(men_men_n72_), .Y(men_men_n189_));
  NO2        u167(.A(men_men_n96_), .B(x06), .Y(men_men_n190_));
  NO2        u168(.A(men_men_n186_), .B(men_men_n36_), .Y(men_men_n191_));
  INV        u169(.A(men_men_n191_), .Y(men_men_n192_));
  NO2        u170(.A(men_men_n190_), .B(men_men_n189_), .Y(men_men_n193_));
  OAI210     u171(.A0(men_men_n193_), .A1(men_men_n188_), .B0(men_men_n185_), .Y(men_men_n194_));
  NOi21      u172(.An(x09), .B(x00), .Y(men_men_n195_));
  NO3        u173(.A(men_men_n84_), .B(men_men_n195_), .C(men_men_n47_), .Y(men_men_n196_));
  NA2        u174(.A(men_men_n196_), .B(men_men_n129_), .Y(men_men_n197_));
  NA2        u175(.A(x06), .B(x05), .Y(men_men_n198_));
  OAI210     u176(.A0(men_men_n198_), .A1(men_men_n35_), .B0(men_men_n101_), .Y(men_men_n199_));
  NA2        u177(.A(men_men_n101_), .B(men_men_n197_), .Y(men_men_n200_));
  NO2        u178(.A(men_men_n102_), .B(x12), .Y(men_men_n201_));
  AOI210     u179(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n201_), .Y(men_men_n202_));
  NA2        u180(.A(men_men_n95_), .B(men_men_n51_), .Y(men_men_n203_));
  NO2        u181(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n204_));
  NA2        u182(.A(men_men_n204_), .B(x02), .Y(men_men_n205_));
  NO2        u183(.A(men_men_n205_), .B(men_men_n203_), .Y(men_men_n206_));
  AOI210     u184(.A0(men_men_n202_), .A1(men_men_n200_), .B0(men_men_n206_), .Y(men_men_n207_));
  NA4        u185(.A(men_men_n207_), .B(men_men_n194_), .C(men_men_n184_), .D(men_men_n172_), .Y(men_men_n208_));
  AOI210     u186(.A0(men_men_n159_), .A1(men_men_n101_), .B0(men_men_n208_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n210_));
  NA2        u188(.A(men_men_n210_), .B(men_men_n139_), .Y(men_men_n211_));
  AOI210     u189(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n212_));
  NO2        u190(.A(men_men_n128_), .B(x06), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n212_), .A1(men_men_n211_), .B0(men_men_n213_), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n214_), .B(x12), .Y(men_men_n215_));
  INV        u193(.A(men_men_n77_), .Y(men_men_n216_));
  NA2        u194(.A(men_men_n163_), .B(men_men_n57_), .Y(men_men_n217_));
  NA2        u195(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n218_));
  NO2        u196(.A(men_men_n95_), .B(x06), .Y(men_men_n219_));
  AOI210     u197(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n220_));
  NA4        u198(.A(men_men_n161_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n221_));
  NA2        u199(.A(men_men_n221_), .B(men_men_n144_), .Y(men_men_n222_));
  NA2        u200(.A(men_men_n222_), .B(x02), .Y(men_men_n223_));
  AOI210     u201(.A0(men_men_n223_), .A1(men_men_n218_), .B0(men_men_n23_), .Y(men_men_n224_));
  OAI210     u202(.A0(men_men_n215_), .A1(men_men_n57_), .B0(men_men_n224_), .Y(men_men_n225_));
  INV        u203(.A(men_men_n144_), .Y(men_men_n226_));
  NO2        u204(.A(men_men_n51_), .B(x03), .Y(men_men_n227_));
  OAI210     u205(.A0(men_men_n80_), .A1(men_men_n36_), .B0(men_men_n123_), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n102_), .B(x03), .Y(men_men_n229_));
  AOI220     u207(.A0(men_men_n229_), .A1(men_men_n228_), .B0(men_men_n77_), .B1(men_men_n227_), .Y(men_men_n230_));
  INV        u208(.A(men_men_n161_), .Y(men_men_n231_));
  NOi21      u209(.An(x13), .B(x04), .Y(men_men_n232_));
  NO3        u210(.A(men_men_n232_), .B(men_men_n77_), .C(men_men_n195_), .Y(men_men_n233_));
  NO2        u211(.A(men_men_n233_), .B(x05), .Y(men_men_n234_));
  AOI220     u212(.A0(men_men_n234_), .A1(men_men_n445_), .B0(men_men_n231_), .B1(men_men_n57_), .Y(men_men_n235_));
  OAI210     u213(.A0(men_men_n230_), .A1(men_men_n226_), .B0(men_men_n235_), .Y(men_men_n236_));
  INV        u214(.A(men_men_n93_), .Y(men_men_n237_));
  NO2        u215(.A(men_men_n237_), .B(x12), .Y(men_men_n238_));
  NA2        u216(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n239_));
  NO2        u217(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n240_));
  INV        u218(.A(men_men_n187_), .Y(men_men_n241_));
  NA2        u219(.A(men_men_n150_), .B(men_men_n73_), .Y(men_men_n242_));
  INV        u220(.A(men_men_n242_), .Y(men_men_n243_));
  NA2        u221(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n244_));
  NA2        u222(.A(men_men_n244_), .B(x03), .Y(men_men_n245_));
  OA210      u223(.A0(men_men_n245_), .A1(men_men_n243_), .B0(men_men_n241_), .Y(men_men_n246_));
  NA2        u224(.A(x13), .B(men_men_n101_), .Y(men_men_n247_));
  NA3        u225(.A(men_men_n247_), .B(men_men_n199_), .C(men_men_n94_), .Y(men_men_n248_));
  OAI210     u226(.A0(men_men_n246_), .A1(men_men_n239_), .B0(men_men_n248_), .Y(men_men_n249_));
  AOI210     u227(.A0(men_men_n238_), .A1(men_men_n236_), .B0(men_men_n249_), .Y(men_men_n250_));
  AOI210     u228(.A0(men_men_n250_), .A1(men_men_n225_), .B0(x07), .Y(men_men_n251_));
  NA2        u229(.A(men_men_n72_), .B(men_men_n29_), .Y(men_men_n252_));
  BUFFER     u230(.A(men_men_n138_), .Y(men_men_n253_));
  AOI210     u231(.A0(men_men_n253_), .A1(men_men_n152_), .B0(men_men_n252_), .Y(men_men_n254_));
  NO2        u232(.A(x08), .B(x05), .Y(men_men_n255_));
  OAI210     u233(.A0(men_men_n77_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n256_));
  INV        u234(.A(men_men_n256_), .Y(men_men_n257_));
  NO2        u235(.A(x12), .B(x02), .Y(men_men_n258_));
  INV        u236(.A(men_men_n258_), .Y(men_men_n259_));
  NO2        u237(.A(men_men_n259_), .B(men_men_n237_), .Y(men_men_n260_));
  OA210      u238(.A0(men_men_n257_), .A1(men_men_n254_), .B0(men_men_n260_), .Y(men_men_n261_));
  NA2        u239(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n262_));
  NO2        u240(.A(men_men_n262_), .B(x01), .Y(men_men_n263_));
  NOi21      u241(.An(men_men_n85_), .B(men_men_n123_), .Y(men_men_n264_));
  NO2        u242(.A(men_men_n264_), .B(men_men_n263_), .Y(men_men_n265_));
  AOI210     u243(.A0(men_men_n265_), .A1(men_men_n132_), .B0(men_men_n29_), .Y(men_men_n266_));
  NA2        u244(.A(men_men_n102_), .B(x04), .Y(men_men_n267_));
  NA2        u245(.A(men_men_n267_), .B(men_men_n28_), .Y(men_men_n268_));
  NO2        u246(.A(men_men_n268_), .B(men_men_n122_), .Y(men_men_n269_));
  NO3        u247(.A(men_men_n92_), .B(x12), .C(x03), .Y(men_men_n270_));
  OAI210     u248(.A0(men_men_n269_), .A1(men_men_n266_), .B0(men_men_n270_), .Y(men_men_n271_));
  AOI210     u249(.A0(men_men_n203_), .A1(men_men_n198_), .B0(men_men_n104_), .Y(men_men_n272_));
  NOi21      u250(.An(men_men_n252_), .B(men_men_n219_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n25_), .B(x00), .Y(men_men_n274_));
  OAI210     u252(.A0(men_men_n273_), .A1(men_men_n272_), .B0(men_men_n274_), .Y(men_men_n275_));
  NO2        u253(.A(men_men_n58_), .B(x05), .Y(men_men_n276_));
  NO3        u254(.A(men_men_n276_), .B(men_men_n220_), .C(men_men_n190_), .Y(men_men_n277_));
  NO2        u255(.A(men_men_n239_), .B(men_men_n28_), .Y(men_men_n278_));
  OAI210     u256(.A0(men_men_n277_), .A1(men_men_n226_), .B0(men_men_n278_), .Y(men_men_n279_));
  NA3        u257(.A(men_men_n279_), .B(men_men_n275_), .C(men_men_n271_), .Y(men_men_n280_));
  NO3        u258(.A(men_men_n280_), .B(men_men_n261_), .C(men_men_n251_), .Y(men_men_n281_));
  OAI210     u259(.A0(men_men_n209_), .A1(men_men_n61_), .B0(men_men_n281_), .Y(men02));
  NOi21      u260(.An(men_men_n233_), .B(men_men_n175_), .Y(men_men_n283_));
  NO2        u261(.A(men_men_n283_), .B(men_men_n32_), .Y(men_men_n284_));
  NA2        u262(.A(men_men_n284_), .B(men_men_n174_), .Y(men_men_n285_));
  INV        u263(.A(men_men_n174_), .Y(men_men_n286_));
  AOI210     u264(.A0(men_men_n118_), .A1(men_men_n87_), .B0(men_men_n220_), .Y(men_men_n287_));
  OAI220     u265(.A0(men_men_n287_), .A1(men_men_n102_), .B0(men_men_n86_), .B1(men_men_n51_), .Y(men_men_n288_));
  AOI220     u266(.A0(men_men_n288_), .A1(men_men_n286_), .B0(men_men_n156_), .B1(men_men_n155_), .Y(men_men_n289_));
  AOI210     u267(.A0(men_men_n289_), .A1(men_men_n285_), .B0(men_men_n48_), .Y(men_men_n290_));
  NO2        u268(.A(x05), .B(x02), .Y(men_men_n291_));
  OAI210     u269(.A0(men_men_n211_), .A1(men_men_n195_), .B0(men_men_n291_), .Y(men_men_n292_));
  AOI220     u270(.A0(men_men_n255_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n293_));
  NA2        u271(.A(men_men_n232_), .B(men_men_n80_), .Y(men_men_n294_));
  AOI210     u272(.A0(men_men_n294_), .A1(men_men_n292_), .B0(men_men_n144_), .Y(men_men_n295_));
  NAi21      u273(.An(men_men_n234_), .B(men_men_n230_), .Y(men_men_n296_));
  NO2        u274(.A(men_men_n244_), .B(men_men_n47_), .Y(men_men_n297_));
  NA2        u275(.A(men_men_n297_), .B(men_men_n296_), .Y(men_men_n298_));
  AN2        u276(.A(men_men_n229_), .B(men_men_n228_), .Y(men_men_n299_));
  OAI210     u277(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n300_));
  NA2        u278(.A(x13), .B(men_men_n28_), .Y(men_men_n301_));
  BUFFER     u279(.A(men_men_n148_), .Y(men_men_n302_));
  AOI210     u280(.A0(men_men_n302_), .A1(men_men_n139_), .B0(men_men_n300_), .Y(men_men_n303_));
  OAI210     u281(.A0(men_men_n303_), .A1(men_men_n299_), .B0(men_men_n96_), .Y(men_men_n304_));
  NA3        u282(.A(men_men_n96_), .B(men_men_n85_), .C(men_men_n227_), .Y(men_men_n305_));
  NA3        u283(.A(men_men_n95_), .B(men_men_n84_), .C(men_men_n42_), .Y(men_men_n306_));
  AOI210     u284(.A0(men_men_n306_), .A1(men_men_n305_), .B0(x04), .Y(men_men_n307_));
  INV        u285(.A(men_men_n155_), .Y(men_men_n308_));
  NO2        u286(.A(men_men_n308_), .B(men_men_n130_), .Y(men_men_n309_));
  AOI210     u287(.A0(men_men_n309_), .A1(x13), .B0(men_men_n307_), .Y(men_men_n310_));
  NA3        u288(.A(men_men_n310_), .B(men_men_n304_), .C(men_men_n298_), .Y(men_men_n311_));
  NO3        u289(.A(men_men_n311_), .B(men_men_n295_), .C(men_men_n290_), .Y(men_men_n312_));
  NA2        u290(.A(men_men_n143_), .B(x03), .Y(men_men_n313_));
  INV        u291(.A(men_men_n186_), .Y(men_men_n314_));
  AOI220     u292(.A0(x08), .A1(men_men_n314_), .B0(men_men_n204_), .B1(x08), .Y(men_men_n315_));
  OAI210     u293(.A0(men_men_n315_), .A1(men_men_n276_), .B0(men_men_n313_), .Y(men_men_n316_));
  NA2        u294(.A(men_men_n316_), .B(men_men_n109_), .Y(men_men_n317_));
  NA2        u295(.A(men_men_n173_), .B(men_men_n167_), .Y(men_men_n318_));
  AN2        u296(.A(men_men_n318_), .B(men_men_n178_), .Y(men_men_n319_));
  NO2        u297(.A(men_men_n131_), .B(men_men_n28_), .Y(men_men_n320_));
  OAI210     u298(.A0(men_men_n320_), .A1(men_men_n319_), .B0(men_men_n110_), .Y(men_men_n321_));
  NA2        u299(.A(men_men_n267_), .B(men_men_n101_), .Y(men_men_n322_));
  NA2        u300(.A(men_men_n101_), .B(men_men_n41_), .Y(men_men_n323_));
  NA3        u301(.A(men_men_n323_), .B(men_men_n322_), .C(men_men_n130_), .Y(men_men_n324_));
  NA4        u302(.A(men_men_n324_), .B(men_men_n321_), .C(men_men_n317_), .D(men_men_n48_), .Y(men_men_n325_));
  INV        u303(.A(men_men_n204_), .Y(men_men_n326_));
  NO2        u304(.A(men_men_n168_), .B(men_men_n40_), .Y(men_men_n327_));
  NA2        u305(.A(men_men_n32_), .B(x05), .Y(men_men_n328_));
  OAI220     u306(.A0(men_men_n328_), .A1(men_men_n327_), .B0(men_men_n326_), .B1(men_men_n59_), .Y(men_men_n329_));
  NA2        u307(.A(men_men_n329_), .B(x02), .Y(men_men_n330_));
  INV        u308(.A(men_men_n240_), .Y(men_men_n331_));
  NA2        u309(.A(men_men_n201_), .B(x04), .Y(men_men_n332_));
  NO3        u310(.A(men_men_n201_), .B(men_men_n166_), .C(men_men_n52_), .Y(men_men_n333_));
  OAI210     u311(.A0(men_men_n150_), .A1(men_men_n36_), .B0(men_men_n101_), .Y(men_men_n334_));
  OAI210     u312(.A0(men_men_n334_), .A1(men_men_n196_), .B0(men_men_n333_), .Y(men_men_n335_));
  NA3        u313(.A(men_men_n335_), .B(men_men_n330_), .C(x06), .Y(men_men_n336_));
  NA2        u314(.A(x09), .B(x03), .Y(men_men_n337_));
  OAI220     u315(.A0(men_men_n337_), .A1(men_men_n129_), .B0(men_men_n210_), .B1(men_men_n63_), .Y(men_men_n338_));
  NO3        u316(.A(men_men_n276_), .B(men_men_n128_), .C(x08), .Y(men_men_n339_));
  INV        u317(.A(men_men_n339_), .Y(men_men_n340_));
  NO2        u318(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n341_));
  NO3        u319(.A(men_men_n116_), .B(men_men_n129_), .C(men_men_n38_), .Y(men_men_n342_));
  AOI210     u320(.A0(men_men_n333_), .A1(men_men_n341_), .B0(men_men_n342_), .Y(men_men_n343_));
  OAI210     u321(.A0(men_men_n340_), .A1(men_men_n28_), .B0(men_men_n343_), .Y(men_men_n344_));
  AO220      u322(.A0(men_men_n344_), .A1(x04), .B0(men_men_n338_), .B1(x05), .Y(men_men_n345_));
  AOI210     u323(.A0(men_men_n336_), .A1(men_men_n325_), .B0(men_men_n345_), .Y(men_men_n346_));
  OAI210     u324(.A0(men_men_n312_), .A1(x12), .B0(men_men_n346_), .Y(men03));
  OR2        u325(.A(men_men_n42_), .B(men_men_n227_), .Y(men_men_n348_));
  AOI210     u326(.A0(men_men_n156_), .A1(men_men_n101_), .B0(men_men_n348_), .Y(men_men_n349_));
  AO210      u327(.A0(men_men_n331_), .A1(men_men_n87_), .B0(men_men_n332_), .Y(men_men_n350_));
  NA2        u328(.A(men_men_n201_), .B(men_men_n155_), .Y(men_men_n351_));
  NA3        u329(.A(men_men_n351_), .B(men_men_n350_), .C(men_men_n205_), .Y(men_men_n352_));
  OAI210     u330(.A0(men_men_n352_), .A1(men_men_n349_), .B0(x05), .Y(men_men_n353_));
  NA2        u331(.A(men_men_n348_), .B(x05), .Y(men_men_n354_));
  AOI210     u332(.A0(men_men_n139_), .A1(men_men_n216_), .B0(men_men_n354_), .Y(men_men_n355_));
  AOI210     u333(.A0(men_men_n229_), .A1(men_men_n81_), .B0(men_men_n125_), .Y(men_men_n356_));
  OAI220     u334(.A0(men_men_n356_), .A1(men_men_n59_), .B0(men_men_n301_), .B1(men_men_n293_), .Y(men_men_n357_));
  OAI210     u335(.A0(men_men_n357_), .A1(men_men_n355_), .B0(men_men_n101_), .Y(men_men_n358_));
  AOI210     u336(.A0(men_men_n148_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n359_));
  NO2        u337(.A(men_men_n175_), .B(men_men_n134_), .Y(men_men_n360_));
  OAI220     u338(.A0(men_men_n360_), .A1(men_men_n37_), .B0(men_men_n151_), .B1(x13), .Y(men_men_n361_));
  OAI210     u339(.A0(men_men_n361_), .A1(men_men_n359_), .B0(x04), .Y(men_men_n362_));
  NO3        u340(.A(men_men_n323_), .B(men_men_n86_), .C(men_men_n59_), .Y(men_men_n363_));
  AOI210     u341(.A0(men_men_n192_), .A1(men_men_n101_), .B0(men_men_n148_), .Y(men_men_n364_));
  OA210      u342(.A0(men_men_n168_), .A1(x12), .B0(men_men_n134_), .Y(men_men_n365_));
  NO3        u343(.A(men_men_n365_), .B(men_men_n364_), .C(men_men_n363_), .Y(men_men_n366_));
  NA4        u344(.A(men_men_n366_), .B(men_men_n362_), .C(men_men_n358_), .D(men_men_n353_), .Y(men04));
  NO2        u345(.A(men_men_n90_), .B(men_men_n39_), .Y(men_men_n368_));
  XO2        u346(.A(men_men_n368_), .B(men_men_n247_), .Y(men05));
  NO2        u347(.A(men_men_n300_), .B(men_men_n25_), .Y(men_men_n370_));
  NA3        u348(.A(men_men_n144_), .B(men_men_n131_), .C(men_men_n31_), .Y(men_men_n371_));
  AOI210     u349(.A0(men_men_n443_), .A1(men_men_n371_), .B0(men_men_n24_), .Y(men_men_n372_));
  OAI210     u350(.A0(men_men_n372_), .A1(men_men_n370_), .B0(men_men_n101_), .Y(men_men_n373_));
  NA2        u351(.A(x11), .B(men_men_n31_), .Y(men_men_n374_));
  NA2        u352(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n375_));
  NA2        u353(.A(men_men_n252_), .B(x03), .Y(men_men_n376_));
  OAI220     u354(.A0(men_men_n376_), .A1(men_men_n375_), .B0(men_men_n374_), .B1(men_men_n82_), .Y(men_men_n377_));
  OAI210     u355(.A0(men_men_n26_), .A1(men_men_n101_), .B0(x07), .Y(men_men_n378_));
  AOI210     u356(.A0(men_men_n377_), .A1(x06), .B0(men_men_n378_), .Y(men_men_n379_));
  AOI220     u357(.A0(men_men_n82_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n380_));
  NO3        u358(.A(men_men_n380_), .B(men_men_n23_), .C(x00), .Y(men_men_n381_));
  NA2        u359(.A(men_men_n70_), .B(x02), .Y(men_men_n382_));
  NA2        u360(.A(men_men_n382_), .B(men_men_n376_), .Y(men_men_n383_));
  OR2        u361(.A(men_men_n383_), .B(men_men_n239_), .Y(men_men_n384_));
  NO2        u362(.A(men_men_n23_), .B(x10), .Y(men_men_n385_));
  OAI210     u363(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n386_));
  OR3        u364(.A(men_men_n386_), .B(men_men_n385_), .C(men_men_n44_), .Y(men_men_n387_));
  NA2        u365(.A(men_men_n387_), .B(men_men_n384_), .Y(men_men_n388_));
  OAI210     u366(.A0(men_men_n388_), .A1(men_men_n381_), .B0(men_men_n101_), .Y(men_men_n389_));
  NA2        u367(.A(men_men_n33_), .B(men_men_n101_), .Y(men_men_n390_));
  AOI210     u368(.A0(men_men_n390_), .A1(men_men_n93_), .B0(x07), .Y(men_men_n391_));
  AOI220     u369(.A0(men_men_n391_), .A1(men_men_n389_), .B0(men_men_n379_), .B1(men_men_n373_), .Y(men_men_n392_));
  NA3        u370(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n393_));
  AO210      u371(.A0(men_men_n393_), .A1(men_men_n262_), .B0(men_men_n259_), .Y(men_men_n394_));
  AOI210     u372(.A0(men_men_n385_), .A1(men_men_n75_), .B0(men_men_n143_), .Y(men_men_n395_));
  OR2        u373(.A(men_men_n395_), .B(x03), .Y(men_men_n396_));
  NA2        u374(.A(men_men_n341_), .B(men_men_n61_), .Y(men_men_n397_));
  NO2        u375(.A(men_men_n397_), .B(x11), .Y(men_men_n398_));
  NO3        u376(.A(men_men_n398_), .B(men_men_n147_), .C(men_men_n28_), .Y(men_men_n399_));
  AOI220     u377(.A0(men_men_n399_), .A1(men_men_n396_), .B0(men_men_n394_), .B1(men_men_n47_), .Y(men_men_n400_));
  NO4        u378(.A(men_men_n323_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n401_));
  OAI210     u379(.A0(men_men_n401_), .A1(men_men_n400_), .B0(men_men_n102_), .Y(men_men_n402_));
  AOI210     u380(.A0(men_men_n332_), .A1(men_men_n112_), .B0(men_men_n258_), .Y(men_men_n403_));
  NOi21      u381(.An(men_men_n313_), .B(men_men_n134_), .Y(men_men_n404_));
  NO2        u382(.A(men_men_n404_), .B(men_men_n259_), .Y(men_men_n405_));
  OAI210     u383(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n406_));
  AOI210     u384(.A0(men_men_n247_), .A1(men_men_n47_), .B0(men_men_n406_), .Y(men_men_n407_));
  NO4        u385(.A(men_men_n407_), .B(men_men_n405_), .C(men_men_n403_), .D(x08), .Y(men_men_n408_));
  NO2        u386(.A(men_men_n385_), .B(men_men_n31_), .Y(men_men_n409_));
  NA2        u387(.A(x09), .B(men_men_n41_), .Y(men_men_n410_));
  OAI220     u388(.A0(men_men_n410_), .A1(men_men_n409_), .B0(men_men_n374_), .B1(men_men_n66_), .Y(men_men_n411_));
  NO2        u389(.A(x13), .B(x12), .Y(men_men_n412_));
  NO2        u390(.A(men_men_n131_), .B(men_men_n28_), .Y(men_men_n413_));
  NO2        u391(.A(men_men_n413_), .B(men_men_n263_), .Y(men_men_n414_));
  OR3        u392(.A(men_men_n414_), .B(x12), .C(x03), .Y(men_men_n415_));
  NA3        u393(.A(men_men_n326_), .B(men_men_n126_), .C(x12), .Y(men_men_n416_));
  AO210      u394(.A0(men_men_n326_), .A1(men_men_n126_), .B0(men_men_n247_), .Y(men_men_n417_));
  NA4        u395(.A(men_men_n417_), .B(men_men_n416_), .C(men_men_n415_), .D(x08), .Y(men_men_n418_));
  AOI210     u396(.A0(men_men_n412_), .A1(men_men_n411_), .B0(men_men_n418_), .Y(men_men_n419_));
  AOI210     u397(.A0(men_men_n408_), .A1(men_men_n402_), .B0(men_men_n419_), .Y(men_men_n420_));
  OAI210     u398(.A0(men_men_n397_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n421_));
  NO2        u399(.A(men_men_n442_), .B(men_men_n375_), .Y(men_men_n422_));
  OAI210     u400(.A0(men_men_n422_), .A1(men_men_n421_), .B0(men_men_n191_), .Y(men_men_n423_));
  NA3        u401(.A(men_men_n414_), .B(men_men_n404_), .C(men_men_n322_), .Y(men_men_n424_));
  INV        u402(.A(x14), .Y(men_men_n425_));
  NO3        u403(.A(men_men_n313_), .B(men_men_n107_), .C(x11), .Y(men_men_n426_));
  NO3        u404(.A(men_men_n167_), .B(men_men_n75_), .C(men_men_n57_), .Y(men_men_n427_));
  NO3        u405(.A(men_men_n393_), .B(men_men_n323_), .C(men_men_n186_), .Y(men_men_n428_));
  NO4        u406(.A(men_men_n428_), .B(men_men_n427_), .C(men_men_n426_), .D(men_men_n425_), .Y(men_men_n429_));
  NA3        u407(.A(men_men_n429_), .B(men_men_n424_), .C(men_men_n423_), .Y(men_men_n430_));
  AOI220     u408(.A0(men_men_n390_), .A1(men_men_n61_), .B0(men_men_n413_), .B1(men_men_n166_), .Y(men_men_n431_));
  NOi21      u409(.An(men_men_n267_), .B(men_men_n151_), .Y(men_men_n432_));
  NO3        u410(.A(men_men_n128_), .B(men_men_n24_), .C(x06), .Y(men_men_n433_));
  AOI210     u411(.A0(men_men_n274_), .A1(men_men_n231_), .B0(men_men_n433_), .Y(men_men_n434_));
  OAI210     u412(.A0(men_men_n44_), .A1(x04), .B0(men_men_n434_), .Y(men_men_n435_));
  OAI210     u413(.A0(men_men_n435_), .A1(men_men_n432_), .B0(men_men_n101_), .Y(men_men_n436_));
  OAI210     u414(.A0(men_men_n431_), .A1(men_men_n92_), .B0(men_men_n436_), .Y(men_men_n437_));
  NO4        u415(.A(men_men_n437_), .B(men_men_n430_), .C(men_men_n420_), .D(men_men_n392_), .Y(men06));
  INV        u416(.A(x07), .Y(men_men_n441_));
  INV        u417(.A(x07), .Y(men_men_n442_));
  INV        u418(.A(men_men_n91_), .Y(men_men_n443_));
  INV        u419(.A(men_men_n94_), .Y(men_men_n444_));
  INV        u420(.A(x06), .Y(men_men_n445_));
  INV        u421(.A(x01), .Y(men_men_n446_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule