// Benchmark "top" written by ABC on Thu Jun 20 14:00:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n137_, new_new_n138_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n338_, new_new_n339_, new_new_n340_, new_new_n341_,
    new_new_n342_, new_new_n343_, new_new_n344_, new_new_n345_,
    new_new_n346_, new_new_n347_, new_new_n348_, new_new_n349_,
    new_new_n350_, new_new_n351_, new_new_n352_, new_new_n353_,
    new_new_n354_, new_new_n355_, new_new_n356_, new_new_n357_,
    new_new_n358_, new_new_n359_, new_new_n360_, new_new_n361_,
    new_new_n362_, new_new_n363_, new_new_n364_, new_new_n365_,
    new_new_n366_, new_new_n367_, new_new_n368_, new_new_n369_,
    new_new_n370_, new_new_n371_, new_new_n372_, new_new_n373_,
    new_new_n374_, new_new_n375_, new_new_n376_, new_new_n377_,
    new_new_n378_, new_new_n379_, new_new_n380_, new_new_n381_,
    new_new_n382_, new_new_n383_, new_new_n384_, new_new_n385_,
    new_new_n386_, new_new_n387_, new_new_n388_, new_new_n389_,
    new_new_n390_, new_new_n391_, new_new_n392_, new_new_n393_,
    new_new_n394_, new_new_n395_, new_new_n396_, new_new_n397_,
    new_new_n398_, new_new_n399_, new_new_n400_, new_new_n401_,
    new_new_n402_, new_new_n403_, new_new_n404_, new_new_n405_,
    new_new_n406_, new_new_n407_, new_new_n408_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n455_, new_new_n456_, new_new_n457_, new_new_n458_,
    new_new_n459_, new_new_n460_, new_new_n461_, new_new_n462_,
    new_new_n463_, new_new_n464_, new_new_n465_, new_new_n466_,
    new_new_n467_, new_new_n468_, new_new_n469_, new_new_n470_,
    new_new_n471_, new_new_n472_, new_new_n473_, new_new_n474_,
    new_new_n475_, new_new_n476_, new_new_n477_, new_new_n478_,
    new_new_n479_, new_new_n480_, new_new_n481_, new_new_n482_,
    new_new_n483_, new_new_n484_, new_new_n485_, new_new_n486_,
    new_new_n487_, new_new_n488_, new_new_n489_, new_new_n490_,
    new_new_n491_, new_new_n492_, new_new_n493_, new_new_n494_,
    new_new_n495_, new_new_n496_, new_new_n497_, new_new_n498_,
    new_new_n499_, new_new_n500_, new_new_n501_, new_new_n503_,
    new_new_n504_, new_new_n505_, new_new_n506_, new_new_n507_,
    new_new_n508_, new_new_n509_, new_new_n510_, new_new_n511_,
    new_new_n512_, new_new_n513_, new_new_n514_, new_new_n515_,
    new_new_n516_, new_new_n517_, new_new_n518_, new_new_n519_,
    new_new_n520_, new_new_n521_, new_new_n522_, new_new_n523_,
    new_new_n524_, new_new_n525_, new_new_n526_, new_new_n527_,
    new_new_n528_, new_new_n529_, new_new_n530_, new_new_n531_,
    new_new_n532_, new_new_n533_, new_new_n534_, new_new_n535_,
    new_new_n536_, new_new_n537_, new_new_n538_, new_new_n539_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n640_, new_new_n641_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(zz01));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  NO2        g036(.A(new_new_n58_), .B(new_new_n57_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g039(.A(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NA3        g041(.A(new_new_n63_), .B(new_new_n61_), .C(new_new_n31_), .Y(new_new_n64_));
  NA2        g042(.A(i_1_), .B(i_10_), .Y(new_new_n65_));
  NO2        g043(.A(new_new_n65_), .B(i_6_), .Y(new_new_n66_));
  NAi31      g044(.An(new_new_n66_), .B(new_new_n64_), .C(new_new_n60_), .Y(new_new_n67_));
  NA2        g045(.A(new_new_n50_), .B(i_2_), .Y(new_new_n68_));
  AOI210     g046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n69_));
  NA2        g047(.A(i_1_), .B(i_6_), .Y(new_new_n70_));
  NO2        g048(.A(new_new_n70_), .B(new_new_n25_), .Y(new_new_n71_));
  INV        g049(.A(i_0_), .Y(new_new_n72_));
  NAi21      g050(.An(i_5_), .B(i_10_), .Y(new_new_n73_));
  NA2        g051(.A(i_5_), .B(i_9_), .Y(new_new_n74_));
  AOI210     g052(.A0(new_new_n74_), .A1(new_new_n73_), .B0(new_new_n72_), .Y(new_new_n75_));
  NO2        g053(.A(new_new_n75_), .B(new_new_n71_), .Y(new_new_n76_));
  OAI210     g054(.A0(new_new_n69_), .A1(new_new_n68_), .B0(new_new_n76_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n77_), .A1(new_new_n67_), .B0(i_0_), .Y(new_new_n78_));
  NA2        g056(.A(i_12_), .B(i_5_), .Y(new_new_n79_));
  NA2        g057(.A(i_2_), .B(i_8_), .Y(new_new_n80_));
  NO2        g058(.A(new_new_n80_), .B(new_new_n57_), .Y(new_new_n81_));
  NO2        g059(.A(i_3_), .B(i_9_), .Y(new_new_n82_));
  NO2        g060(.A(i_3_), .B(i_7_), .Y(new_new_n83_));
  NO2        g061(.A(new_new_n82_), .B(new_new_n62_), .Y(new_new_n84_));
  INV        g062(.A(i_6_), .Y(new_new_n85_));
  NO2        g063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  INV        g064(.A(new_new_n86_), .Y(new_new_n87_));
  OAI210     g065(.A0(new_new_n84_), .A1(new_new_n81_), .B0(new_new_n87_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n62_), .Y(new_new_n91_));
  NA2        g069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  NO3        g070(.A(new_new_n92_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n93_));
  NO2        g071(.A(new_new_n93_), .B(new_new_n91_), .Y(new_new_n94_));
  AOI210     g072(.A0(new_new_n94_), .A1(new_new_n88_), .B0(new_new_n79_), .Y(new_new_n95_));
  AN3        g073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NO2        g075(.A(i_5_), .B(i_8_), .Y(new_new_n98_));
  NOi21      g076(.An(new_new_n98_), .B(new_new_n97_), .Y(new_new_n99_));
  AOI220     g077(.A0(new_new_n99_), .A1(new_new_n61_), .B0(new_new_n96_), .B1(new_new_n32_), .Y(new_new_n100_));
  INV        g078(.A(i_7_), .Y(new_new_n101_));
  NA2        g079(.A(new_new_n46_), .B(new_new_n101_), .Y(new_new_n102_));
  NO2        g080(.A(i_0_), .B(i_5_), .Y(new_new_n103_));
  NO2        g081(.A(new_new_n103_), .B(new_new_n85_), .Y(new_new_n104_));
  NA2        g082(.A(i_12_), .B(i_3_), .Y(new_new_n105_));
  INV        g083(.A(new_new_n105_), .Y(new_new_n106_));
  NA3        g084(.A(new_new_n106_), .B(new_new_n104_), .C(new_new_n102_), .Y(new_new_n107_));
  NAi21      g085(.An(i_7_), .B(i_11_), .Y(new_new_n108_));
  AN2        g086(.A(i_2_), .B(i_10_), .Y(new_new_n109_));
  NO2        g087(.A(new_new_n109_), .B(i_7_), .Y(new_new_n110_));
  OR2        g088(.A(new_new_n79_), .B(new_new_n57_), .Y(new_new_n111_));
  NO2        g089(.A(i_8_), .B(new_new_n101_), .Y(new_new_n112_));
  NO3        g090(.A(new_new_n112_), .B(new_new_n111_), .C(new_new_n110_), .Y(new_new_n113_));
  NA2        g091(.A(i_12_), .B(i_7_), .Y(new_new_n114_));
  NO2        g092(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n115_));
  NA2        g093(.A(i_11_), .B(i_12_), .Y(new_new_n116_));
  INV        g094(.A(new_new_n116_), .Y(new_new_n117_));
  NO2        g095(.A(new_new_n117_), .B(new_new_n113_), .Y(new_new_n118_));
  NA3        g096(.A(new_new_n118_), .B(new_new_n107_), .C(new_new_n100_), .Y(new_new_n119_));
  NOi21      g097(.An(i_1_), .B(i_5_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(i_11_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n122_));
  NA2        g100(.A(i_7_), .B(new_new_n25_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n122_), .Y(new_new_n124_));
  NO2        g102(.A(new_new_n124_), .B(new_new_n46_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n126_));
  NAi21      g104(.An(i_3_), .B(i_8_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(new_new_n61_), .Y(new_new_n128_));
  NOi31      g106(.An(new_new_n128_), .B(new_new_n126_), .C(new_new_n125_), .Y(new_new_n129_));
  NO2        g107(.A(i_1_), .B(new_new_n85_), .Y(new_new_n130_));
  NO2        g108(.A(i_6_), .B(i_5_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(i_3_), .Y(new_new_n132_));
  AO210      g110(.A0(new_new_n132_), .A1(new_new_n47_), .B0(new_new_n130_), .Y(new_new_n133_));
  OAI220     g111(.A0(new_new_n133_), .A1(new_new_n108_), .B0(new_new_n129_), .B1(new_new_n121_), .Y(new_new_n134_));
  NO3        g112(.A(new_new_n134_), .B(new_new_n119_), .C(new_new_n95_), .Y(new_new_n135_));
  NA3        g113(.A(new_new_n135_), .B(new_new_n78_), .C(new_new_n56_), .Y(zz02));
  NO2        g114(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n137_));
  NA2        g115(.A(new_new_n641_), .B(new_new_n137_), .Y(new_new_n138_));
  NA4        g116(.A(new_new_n138_), .B(new_new_n76_), .C(new_new_n68_), .D(new_new_n30_), .Y(zz00));
  AN2        g117(.A(i_8_), .B(i_7_), .Y(new_new_n140_));
  NA2        g118(.A(new_new_n140_), .B(i_6_), .Y(new_new_n141_));
  NO2        g119(.A(i_12_), .B(i_13_), .Y(new_new_n142_));
  NAi21      g120(.An(i_5_), .B(i_11_), .Y(new_new_n143_));
  NO2        g121(.A(i_0_), .B(i_1_), .Y(new_new_n144_));
  NA2        g122(.A(i_2_), .B(i_3_), .Y(new_new_n145_));
  NO2        g123(.A(new_new_n145_), .B(i_4_), .Y(new_new_n146_));
  AN2        g124(.A(new_new_n142_), .B(new_new_n82_), .Y(new_new_n147_));
  NA2        g125(.A(i_1_), .B(i_5_), .Y(new_new_n148_));
  OR2        g126(.A(i_0_), .B(i_1_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n149_), .B(new_new_n79_), .C(i_13_), .Y(new_new_n150_));
  NAi32      g128(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n151_));
  NAi21      g129(.An(new_new_n151_), .B(new_new_n150_), .Y(new_new_n152_));
  NOi21      g130(.An(i_4_), .B(i_10_), .Y(new_new_n153_));
  NOi21      g131(.An(i_4_), .B(i_9_), .Y(new_new_n154_));
  NOi21      g132(.An(i_11_), .B(i_13_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n154_), .Y(new_new_n156_));
  NO2        g134(.A(new_new_n72_), .B(new_new_n62_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n72_), .B(i_5_), .Y(new_new_n158_));
  NO2        g136(.A(i_2_), .B(i_1_), .Y(new_new_n159_));
  NAi21      g137(.An(i_4_), .B(i_12_), .Y(new_new_n160_));
  INV        g138(.A(i_8_), .Y(new_new_n161_));
  NO2        g139(.A(i_3_), .B(i_8_), .Y(new_new_n162_));
  NO3        g140(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n103_), .B(new_new_n57_), .Y(new_new_n164_));
  NO2        g142(.A(i_13_), .B(i_9_), .Y(new_new_n165_));
  NAi21      g143(.An(i_12_), .B(i_3_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n44_), .B(i_5_), .Y(new_new_n167_));
  NAi21      g145(.An(i_12_), .B(i_7_), .Y(new_new_n168_));
  NA3        g146(.A(i_13_), .B(new_new_n161_), .C(i_10_), .Y(new_new_n169_));
  NA2        g147(.A(i_0_), .B(i_5_), .Y(new_new_n170_));
  NAi31      g148(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n171_));
  NO2        g149(.A(new_new_n36_), .B(i_13_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n72_), .B(new_new_n26_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n46_), .B(new_new_n62_), .Y(new_new_n174_));
  INV        g152(.A(i_13_), .Y(new_new_n175_));
  NO2        g153(.A(i_12_), .B(new_new_n175_), .Y(new_new_n176_));
  NO2        g154(.A(i_12_), .B(new_new_n37_), .Y(new_new_n177_));
  OR2        g155(.A(i_8_), .B(i_7_), .Y(new_new_n178_));
  INV        g156(.A(i_12_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n44_), .B(new_new_n179_), .Y(new_new_n180_));
  NO3        g158(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n181_));
  NA2        g159(.A(i_2_), .B(i_1_), .Y(new_new_n182_));
  NO3        g160(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n183_));
  NAi21      g161(.An(i_4_), .B(i_3_), .Y(new_new_n184_));
  NO2        g162(.A(i_0_), .B(i_6_), .Y(new_new_n185_));
  NOi41      g163(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n186_));
  NO2        g164(.A(i_11_), .B(new_new_n175_), .Y(new_new_n187_));
  NOi21      g165(.An(i_1_), .B(i_6_), .Y(new_new_n188_));
  NAi21      g166(.An(i_3_), .B(i_7_), .Y(new_new_n189_));
  NA2        g167(.A(new_new_n179_), .B(i_9_), .Y(new_new_n190_));
  OR4        g168(.A(new_new_n190_), .B(new_new_n189_), .C(new_new_n188_), .D(new_new_n158_), .Y(new_new_n191_));
  NA2        g169(.A(new_new_n72_), .B(i_5_), .Y(new_new_n192_));
  NA2        g170(.A(i_3_), .B(i_9_), .Y(new_new_n193_));
  NAi21      g171(.An(i_7_), .B(i_10_), .Y(new_new_n194_));
  NO2        g172(.A(new_new_n194_), .B(new_new_n193_), .Y(new_new_n195_));
  NA3        g173(.A(new_new_n195_), .B(new_new_n192_), .C(new_new_n63_), .Y(new_new_n196_));
  NA2        g174(.A(new_new_n196_), .B(new_new_n191_), .Y(new_new_n197_));
  INV        g175(.A(new_new_n141_), .Y(new_new_n198_));
  NA2        g176(.A(new_new_n179_), .B(i_13_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n199_), .B(new_new_n74_), .Y(new_new_n200_));
  AOI220     g178(.A0(new_new_n200_), .A1(new_new_n198_), .B0(new_new_n197_), .B1(new_new_n187_), .Y(new_new_n201_));
  NA2        g179(.A(i_12_), .B(i_6_), .Y(new_new_n202_));
  OR2        g180(.A(i_13_), .B(i_9_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n184_), .B(i_2_), .Y(new_new_n204_));
  NA2        g182(.A(new_new_n187_), .B(i_9_), .Y(new_new_n205_));
  NO3        g183(.A(i_11_), .B(new_new_n175_), .C(new_new_n25_), .Y(new_new_n206_));
  NO2        g184(.A(new_new_n189_), .B(i_8_), .Y(new_new_n207_));
  NO3        g185(.A(i_12_), .B(new_new_n175_), .C(new_new_n37_), .Y(new_new_n208_));
  NO2        g186(.A(i_2_), .B(new_new_n101_), .Y(new_new_n209_));
  AN2        g187(.A(i_3_), .B(i_10_), .Y(new_new_n210_));
  NO2        g188(.A(i_5_), .B(new_new_n37_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n212_));
  NO3        g190(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n213_));
  NO2        g191(.A(i_2_), .B(i_3_), .Y(new_new_n214_));
  OR2        g192(.A(i_0_), .B(i_5_), .Y(new_new_n215_));
  NO2        g193(.A(i_12_), .B(i_10_), .Y(new_new_n216_));
  NOi21      g194(.An(i_5_), .B(i_0_), .Y(new_new_n217_));
  NO2        g195(.A(i_1_), .B(i_7_), .Y(new_new_n218_));
  NOi21      g196(.An(new_new_n148_), .B(new_new_n104_), .Y(new_new_n219_));
  NOi32      g197(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n220_));
  INV        g198(.A(new_new_n220_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n151_), .B(new_new_n149_), .Y(new_new_n222_));
  NOi32      g200(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n223_));
  NAi21      g201(.An(i_6_), .B(i_1_), .Y(new_new_n224_));
  NO2        g202(.A(i_1_), .B(new_new_n101_), .Y(new_new_n225_));
  NAi21      g203(.An(i_3_), .B(i_4_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n226_), .B(i_9_), .Y(new_new_n227_));
  AN2        g205(.A(i_6_), .B(i_7_), .Y(new_new_n228_));
  OAI210     g206(.A0(new_new_n228_), .A1(new_new_n225_), .B0(new_new_n227_), .Y(new_new_n229_));
  NA2        g207(.A(i_2_), .B(i_7_), .Y(new_new_n230_));
  NO2        g208(.A(new_new_n226_), .B(i_10_), .Y(new_new_n231_));
  NA3        g209(.A(new_new_n231_), .B(new_new_n230_), .C(new_new_n185_), .Y(new_new_n232_));
  AOI210     g210(.A0(new_new_n232_), .A1(new_new_n229_), .B0(new_new_n158_), .Y(new_new_n233_));
  AOI210     g211(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n234_));
  OAI210     g212(.A0(new_new_n234_), .A1(new_new_n159_), .B0(new_new_n231_), .Y(new_new_n235_));
  AOI220     g213(.A0(new_new_n231_), .A1(new_new_n218_), .B0(new_new_n181_), .B1(new_new_n159_), .Y(new_new_n236_));
  AOI210     g214(.A0(new_new_n236_), .A1(new_new_n235_), .B0(i_5_), .Y(new_new_n237_));
  NO3        g215(.A(new_new_n237_), .B(new_new_n233_), .C(new_new_n222_), .Y(new_new_n238_));
  NO2        g216(.A(new_new_n238_), .B(new_new_n221_), .Y(new_new_n239_));
  AN2        g217(.A(i_12_), .B(i_5_), .Y(new_new_n240_));
  NO2        g218(.A(i_11_), .B(i_6_), .Y(new_new_n241_));
  NO2        g219(.A(i_5_), .B(i_10_), .Y(new_new_n242_));
  NO2        g220(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n243_));
  NO3        g221(.A(new_new_n85_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n244_));
  NO2        g222(.A(i_11_), .B(i_12_), .Y(new_new_n245_));
  NAi21      g223(.An(i_13_), .B(i_0_), .Y(new_new_n246_));
  NO3        g224(.A(i_1_), .B(i_12_), .C(new_new_n85_), .Y(new_new_n247_));
  NO2        g225(.A(i_0_), .B(i_11_), .Y(new_new_n248_));
  AN2        g226(.A(i_1_), .B(i_6_), .Y(new_new_n249_));
  NOi21      g227(.An(i_2_), .B(i_12_), .Y(new_new_n250_));
  NAi21      g228(.An(i_9_), .B(i_4_), .Y(new_new_n251_));
  OR2        g229(.A(i_13_), .B(i_10_), .Y(new_new_n252_));
  NO3        g230(.A(new_new_n252_), .B(new_new_n116_), .C(new_new_n251_), .Y(new_new_n253_));
  NO2        g231(.A(new_new_n101_), .B(new_new_n25_), .Y(new_new_n254_));
  NA2        g232(.A(new_new_n208_), .B(new_new_n254_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n255_), .B(new_new_n219_), .Y(new_new_n256_));
  INV        g234(.A(new_new_n256_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n257_), .B(new_new_n26_), .Y(new_new_n258_));
  NA2        g236(.A(new_new_n161_), .B(i_10_), .Y(new_new_n259_));
  NA3        g237(.A(new_new_n192_), .B(new_new_n63_), .C(i_2_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n260_), .B(new_new_n259_), .Y(new_new_n261_));
  INV        g239(.A(new_new_n261_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n262_), .B(new_new_n205_), .Y(new_new_n263_));
  NO3        g241(.A(new_new_n263_), .B(new_new_n258_), .C(new_new_n239_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n72_), .B(i_13_), .Y(new_new_n265_));
  NO2        g243(.A(i_10_), .B(i_9_), .Y(new_new_n266_));
  NAi21      g244(.An(i_12_), .B(i_8_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n267_), .B(i_3_), .Y(new_new_n268_));
  NO3        g246(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n269_));
  NA2        g247(.A(new_new_n202_), .B(new_new_n97_), .Y(new_new_n270_));
  NA2        g248(.A(new_new_n270_), .B(new_new_n269_), .Y(new_new_n271_));
  NA2        g249(.A(i_8_), .B(i_9_), .Y(new_new_n272_));
  AOI210     g250(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n273_));
  OR2        g251(.A(new_new_n273_), .B(new_new_n272_), .Y(new_new_n274_));
  NA2        g252(.A(new_new_n208_), .B(new_new_n164_), .Y(new_new_n275_));
  NO2        g253(.A(new_new_n275_), .B(new_new_n274_), .Y(new_new_n276_));
  NA2        g254(.A(new_new_n187_), .B(new_new_n211_), .Y(new_new_n277_));
  NO3        g255(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n278_));
  INV        g256(.A(new_new_n278_), .Y(new_new_n279_));
  NA3        g257(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n280_));
  NA4        g258(.A(new_new_n143_), .B(new_new_n115_), .C(new_new_n79_), .D(new_new_n23_), .Y(new_new_n281_));
  OAI220     g259(.A0(new_new_n281_), .A1(new_new_n280_), .B0(new_new_n279_), .B1(new_new_n277_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n282_), .B(new_new_n276_), .Y(new_new_n283_));
  NA2        g261(.A(new_new_n96_), .B(i_13_), .Y(new_new_n284_));
  NO2        g262(.A(i_11_), .B(i_1_), .Y(new_new_n285_));
  NOi21      g263(.An(i_2_), .B(i_7_), .Y(new_new_n286_));
  NO2        g264(.A(i_6_), .B(i_10_), .Y(new_new_n287_));
  NA3        g265(.A(new_new_n186_), .B(new_new_n155_), .C(new_new_n131_), .Y(new_new_n288_));
  NA2        g266(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n289_));
  NO2        g267(.A(new_new_n149_), .B(i_3_), .Y(new_new_n290_));
  NAi31      g268(.An(new_new_n289_), .B(new_new_n290_), .C(new_new_n176_), .Y(new_new_n291_));
  NA3        g269(.A(new_new_n243_), .B(new_new_n157_), .C(new_new_n146_), .Y(new_new_n292_));
  NA3        g270(.A(new_new_n292_), .B(new_new_n291_), .C(new_new_n288_), .Y(new_new_n293_));
  INV        g271(.A(new_new_n293_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n278_), .B(new_new_n242_), .Y(new_new_n295_));
  NAi21      g273(.An(new_new_n169_), .B(new_new_n245_), .Y(new_new_n296_));
  NA2        g274(.A(new_new_n27_), .B(i_10_), .Y(new_new_n297_));
  NA2        g275(.A(new_new_n213_), .B(new_new_n181_), .Y(new_new_n298_));
  OAI220     g276(.A0(new_new_n298_), .A1(new_new_n260_), .B0(new_new_n297_), .B1(new_new_n284_), .Y(new_new_n299_));
  INV        g277(.A(new_new_n299_), .Y(new_new_n300_));
  NA3        g278(.A(new_new_n300_), .B(new_new_n294_), .C(new_new_n283_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n240_), .B(new_new_n175_), .Y(new_new_n302_));
  NA2        g280(.A(new_new_n228_), .B(new_new_n223_), .Y(new_new_n303_));
  OR2        g281(.A(new_new_n302_), .B(new_new_n303_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n36_), .B(i_8_), .Y(new_new_n305_));
  AOI210     g283(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n253_), .Y(new_new_n306_));
  NA2        g284(.A(new_new_n306_), .B(new_new_n304_), .Y(new_new_n307_));
  NO2        g285(.A(i_12_), .B(new_new_n161_), .Y(new_new_n308_));
  NA2        g286(.A(new_new_n44_), .B(i_10_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n309_), .B(i_6_), .Y(new_new_n310_));
  NO2        g288(.A(new_new_n149_), .B(i_5_), .Y(new_new_n311_));
  NA3        g289(.A(new_new_n170_), .B(new_new_n70_), .C(new_new_n44_), .Y(new_new_n312_));
  NA2        g290(.A(new_new_n208_), .B(new_new_n83_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n312_), .B(new_new_n313_), .Y(new_new_n314_));
  NA2        g292(.A(new_new_n174_), .B(new_new_n173_), .Y(new_new_n315_));
  NA2        g293(.A(new_new_n266_), .B(new_new_n172_), .Y(new_new_n316_));
  NO2        g294(.A(new_new_n315_), .B(new_new_n316_), .Y(new_new_n317_));
  AOI210     g295(.A0(new_new_n224_), .A1(new_new_n46_), .B0(new_new_n225_), .Y(new_new_n318_));
  NA2        g296(.A(i_0_), .B(new_new_n48_), .Y(new_new_n319_));
  NA3        g297(.A(new_new_n308_), .B(new_new_n206_), .C(new_new_n319_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n318_), .B(new_new_n320_), .Y(new_new_n321_));
  NO3        g299(.A(new_new_n321_), .B(new_new_n317_), .C(new_new_n314_), .Y(new_new_n322_));
  NO3        g300(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n252_), .B(i_1_), .Y(new_new_n324_));
  NOi31      g302(.An(new_new_n324_), .B(new_new_n270_), .C(new_new_n72_), .Y(new_new_n325_));
  NOi21      g303(.An(i_10_), .B(i_6_), .Y(new_new_n326_));
  NO2        g304(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n114_), .B(new_new_n23_), .Y(new_new_n328_));
  NO2        g306(.A(i_12_), .B(new_new_n85_), .Y(new_new_n329_));
  OR2        g307(.A(i_2_), .B(i_5_), .Y(new_new_n330_));
  OR2        g308(.A(new_new_n330_), .B(new_new_n249_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n230_), .B(new_new_n185_), .Y(new_new_n332_));
  AOI210     g310(.A0(new_new_n332_), .A1(new_new_n331_), .B0(new_new_n296_), .Y(new_new_n333_));
  INV        g311(.A(new_new_n333_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n334_), .B(new_new_n322_), .Y(new_new_n335_));
  NO3        g313(.A(new_new_n335_), .B(new_new_n307_), .C(new_new_n301_), .Y(new_new_n336_));
  NA3        g314(.A(new_new_n336_), .B(new_new_n264_), .C(new_new_n201_), .Y(zz07));
  NO2        g315(.A(new_new_n92_), .B(new_new_n54_), .Y(new_new_n338_));
  NA2        g316(.A(new_new_n287_), .B(new_new_n83_), .Y(new_new_n339_));
  NA2        g317(.A(i_11_), .B(new_new_n161_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n142_), .B(new_new_n340_), .Y(new_new_n341_));
  NO2        g319(.A(new_new_n341_), .B(new_new_n339_), .Y(new_new_n342_));
  NA3        g320(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n343_));
  NO2        g321(.A(new_new_n179_), .B(i_4_), .Y(new_new_n344_));
  NA2        g322(.A(new_new_n344_), .B(i_8_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n105_), .B(new_new_n343_), .Y(new_new_n346_));
  NA2        g324(.A(i_2_), .B(new_new_n85_), .Y(new_new_n347_));
  OAI210     g325(.A0(new_new_n86_), .A1(new_new_n162_), .B0(new_new_n163_), .Y(new_new_n348_));
  NO2        g326(.A(i_7_), .B(new_new_n37_), .Y(new_new_n349_));
  NA2        g327(.A(i_4_), .B(i_8_), .Y(new_new_n350_));
  AOI210     g328(.A0(new_new_n350_), .A1(new_new_n210_), .B0(new_new_n349_), .Y(new_new_n351_));
  OAI220     g329(.A0(new_new_n351_), .A1(new_new_n347_), .B0(new_new_n348_), .B1(i_13_), .Y(new_new_n352_));
  NO4        g330(.A(new_new_n352_), .B(new_new_n346_), .C(new_new_n342_), .D(new_new_n338_), .Y(new_new_n353_));
  AOI210     g331(.A0(new_new_n127_), .A1(new_new_n61_), .B0(i_10_), .Y(new_new_n354_));
  AOI210     g332(.A0(new_new_n354_), .A1(new_new_n179_), .B0(new_new_n153_), .Y(new_new_n355_));
  OR2        g333(.A(i_6_), .B(i_10_), .Y(new_new_n356_));
  OR3        g334(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n357_));
  OR2        g335(.A(new_new_n355_), .B(new_new_n203_), .Y(new_new_n358_));
  AOI210     g336(.A0(new_new_n358_), .A1(new_new_n353_), .B0(new_new_n62_), .Y(new_new_n359_));
  NOi21      g337(.An(i_11_), .B(i_7_), .Y(new_new_n360_));
  AO210      g338(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n361_), .B(new_new_n360_), .Y(new_new_n362_));
  NA2        g340(.A(new_new_n362_), .B(new_new_n165_), .Y(new_new_n363_));
  NA3        g341(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n363_), .B(new_new_n62_), .Y(new_new_n365_));
  OR2        g343(.A(new_new_n236_), .B(new_new_n41_), .Y(new_new_n366_));
  NO3        g344(.A(new_new_n194_), .B(new_new_n166_), .C(new_new_n340_), .Y(new_new_n367_));
  OAI210     g345(.A0(new_new_n367_), .A1(new_new_n176_), .B0(new_new_n62_), .Y(new_new_n368_));
  OR2        g346(.A(new_new_n166_), .B(new_new_n108_), .Y(new_new_n369_));
  NO2        g347(.A(i_1_), .B(i_12_), .Y(new_new_n370_));
  NA3        g348(.A(new_new_n370_), .B(new_new_n109_), .C(new_new_n24_), .Y(new_new_n371_));
  BUFFER     g349(.A(new_new_n371_), .Y(new_new_n372_));
  NA3        g350(.A(new_new_n372_), .B(new_new_n368_), .C(new_new_n366_), .Y(new_new_n373_));
  OAI210     g351(.A0(new_new_n373_), .A1(new_new_n365_), .B0(i_6_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n364_), .B(new_new_n108_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n375_), .B(new_new_n329_), .Y(new_new_n376_));
  NO2        g354(.A(i_6_), .B(i_11_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n376_), .B(new_new_n271_), .Y(new_new_n378_));
  NO3        g356(.A(new_new_n356_), .B(new_new_n178_), .C(new_new_n23_), .Y(new_new_n379_));
  AOI210     g357(.A0(i_1_), .A1(new_new_n195_), .B0(new_new_n379_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n380_), .B(new_new_n44_), .Y(new_new_n381_));
  INV        g359(.A(i_2_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n137_), .B(i_9_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n46_), .B(i_1_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n383_), .B(new_new_n382_), .Y(new_new_n385_));
  AOI210     g363(.A0(new_new_n285_), .A1(new_new_n254_), .B0(new_new_n183_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n386_), .B(new_new_n347_), .Y(new_new_n387_));
  NO2        g365(.A(i_11_), .B(new_new_n37_), .Y(new_new_n388_));
  OR2        g366(.A(new_new_n387_), .B(new_new_n385_), .Y(new_new_n389_));
  NO3        g367(.A(new_new_n389_), .B(new_new_n381_), .C(new_new_n378_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n179_), .B(new_new_n101_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n391_), .B(new_new_n360_), .Y(new_new_n392_));
  NA2        g370(.A(new_new_n392_), .B(i_1_), .Y(new_new_n393_));
  NO2        g371(.A(new_new_n393_), .B(new_new_n357_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n251_), .B(new_new_n85_), .Y(new_new_n395_));
  NA2        g373(.A(new_new_n394_), .B(new_new_n46_), .Y(new_new_n396_));
  NA2        g374(.A(i_3_), .B(new_new_n161_), .Y(new_new_n397_));
  NO2        g375(.A(new_new_n397_), .B(new_new_n114_), .Y(new_new_n398_));
  AN2        g376(.A(new_new_n398_), .B(new_new_n310_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n178_), .B(new_new_n44_), .Y(new_new_n400_));
  NO3        g378(.A(new_new_n400_), .B(new_new_n212_), .C(new_new_n180_), .Y(new_new_n401_));
  NO2        g379(.A(new_new_n116_), .B(new_new_n37_), .Y(new_new_n402_));
  NO2        g380(.A(new_new_n402_), .B(i_6_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n85_), .B(i_9_), .Y(new_new_n404_));
  NO2        g382(.A(new_new_n404_), .B(new_new_n62_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n405_), .B(new_new_n370_), .Y(new_new_n406_));
  NO4        g384(.A(new_new_n406_), .B(new_new_n403_), .C(new_new_n401_), .D(i_4_), .Y(new_new_n407_));
  NA2        g385(.A(i_1_), .B(i_3_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n272_), .B(new_new_n92_), .Y(new_new_n409_));
  AOI210     g387(.A0(new_new_n400_), .A1(new_new_n326_), .B0(new_new_n409_), .Y(new_new_n410_));
  NO2        g388(.A(new_new_n410_), .B(new_new_n408_), .Y(new_new_n411_));
  NO3        g389(.A(new_new_n411_), .B(new_new_n407_), .C(new_new_n399_), .Y(new_new_n412_));
  NA4        g390(.A(new_new_n412_), .B(new_new_n396_), .C(new_new_n390_), .D(new_new_n374_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n414_));
  INV        g392(.A(new_new_n414_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n415_), .B(i_1_), .Y(new_new_n416_));
  AOI210     g394(.A0(new_new_n202_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n417_));
  NO2        g395(.A(new_new_n226_), .B(i_2_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n418_), .B(new_new_n417_), .Y(new_new_n419_));
  AOI210     g397(.A0(new_new_n419_), .A1(new_new_n416_), .B0(i_13_), .Y(new_new_n420_));
  OR2        g398(.A(i_11_), .B(i_7_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n54_), .B(i_12_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n286_), .B(new_new_n24_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n423_), .B(new_new_n395_), .Y(new_new_n424_));
  OAI220     g402(.A0(new_new_n424_), .A1(new_new_n41_), .B0(new_new_n640_), .B1(new_new_n92_), .Y(new_new_n425_));
  INV        g403(.A(new_new_n425_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n241_), .B(new_new_n384_), .Y(new_new_n427_));
  NO2        g405(.A(new_new_n427_), .B(new_new_n184_), .Y(new_new_n428_));
  AOI210     g406(.A0(new_new_n267_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n429_));
  NOi31      g407(.An(new_new_n429_), .B(new_new_n339_), .C(new_new_n44_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n126_), .B(i_13_), .Y(new_new_n431_));
  NO2        g409(.A(new_new_n431_), .B(new_new_n417_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n26_), .B(new_new_n161_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n433_), .B(i_7_), .Y(new_new_n434_));
  AOI220     g412(.A0(new_new_n241_), .A1(new_new_n384_), .B0(new_new_n91_), .B1(new_new_n102_), .Y(new_new_n435_));
  NO2        g413(.A(new_new_n435_), .B(new_new_n345_), .Y(new_new_n436_));
  NO4        g414(.A(new_new_n436_), .B(new_new_n432_), .C(new_new_n430_), .D(new_new_n428_), .Y(new_new_n437_));
  OR2        g415(.A(i_11_), .B(i_6_), .Y(new_new_n438_));
  NA3        g416(.A(new_new_n344_), .B(new_new_n433_), .C(i_7_), .Y(new_new_n439_));
  NO2        g417(.A(new_new_n439_), .B(new_new_n438_), .Y(new_new_n440_));
  NA3        g418(.A(new_new_n250_), .B(new_new_n349_), .C(new_new_n97_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n377_), .B(i_13_), .Y(new_new_n442_));
  NAi21      g420(.An(i_11_), .B(i_12_), .Y(new_new_n443_));
  NOi41      g421(.An(new_new_n110_), .B(new_new_n443_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n444_), .B(new_new_n46_), .Y(new_new_n445_));
  NA3        g423(.A(new_new_n445_), .B(new_new_n442_), .C(new_new_n441_), .Y(new_new_n446_));
  OAI210     g424(.A0(new_new_n446_), .A1(new_new_n440_), .B0(new_new_n62_), .Y(new_new_n447_));
  NO2        g425(.A(i_2_), .B(i_12_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n225_), .B(new_new_n448_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n227_), .B(new_new_n225_), .Y(new_new_n450_));
  NA2        g428(.A(new_new_n450_), .B(new_new_n449_), .Y(new_new_n451_));
  NA3        g429(.A(new_new_n451_), .B(new_new_n45_), .C(new_new_n175_), .Y(new_new_n452_));
  NA4        g430(.A(new_new_n452_), .B(new_new_n447_), .C(new_new_n437_), .D(new_new_n426_), .Y(new_new_n453_));
  OR4        g431(.A(new_new_n453_), .B(new_new_n420_), .C(new_new_n413_), .D(new_new_n359_), .Y(zz05));
  NA2        g432(.A(new_new_n392_), .B(new_new_n204_), .Y(new_new_n455_));
  AN2        g433(.A(new_new_n24_), .B(i_10_), .Y(new_new_n456_));
  NA3        g434(.A(new_new_n456_), .B(new_new_n448_), .C(new_new_n108_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n345_), .B(i_11_), .Y(new_new_n458_));
  NA2        g436(.A(new_new_n86_), .B(new_new_n458_), .Y(new_new_n459_));
  NA3        g437(.A(new_new_n459_), .B(new_new_n457_), .C(new_new_n455_), .Y(new_new_n460_));
  NO3        g438(.A(i_11_), .B(new_new_n179_), .C(i_13_), .Y(new_new_n461_));
  NO2        g439(.A(new_new_n123_), .B(new_new_n23_), .Y(new_new_n462_));
  NA2        g440(.A(i_12_), .B(i_8_), .Y(new_new_n463_));
  OAI210     g441(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n463_), .Y(new_new_n464_));
  INV        g442(.A(new_new_n266_), .Y(new_new_n465_));
  AOI220     g443(.A0(new_new_n214_), .A1(new_new_n328_), .B0(new_new_n464_), .B1(new_new_n462_), .Y(new_new_n466_));
  INV        g444(.A(new_new_n466_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n467_), .B(new_new_n460_), .Y(new_new_n468_));
  INV        g446(.A(new_new_n155_), .Y(new_new_n469_));
  INV        g447(.A(new_new_n186_), .Y(new_new_n470_));
  OAI210     g448(.A0(new_new_n418_), .A1(new_new_n268_), .B0(new_new_n110_), .Y(new_new_n471_));
  AOI210     g449(.A0(new_new_n471_), .A1(new_new_n470_), .B0(new_new_n469_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n272_), .B(new_new_n26_), .Y(new_new_n473_));
  NO2        g451(.A(new_new_n473_), .B(new_new_n254_), .Y(new_new_n474_));
  NA2        g452(.A(new_new_n474_), .B(i_2_), .Y(new_new_n475_));
  INV        g453(.A(new_new_n475_), .Y(new_new_n476_));
  AOI210     g454(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n252_), .Y(new_new_n477_));
  AOI210     g455(.A0(new_new_n477_), .A1(new_new_n476_), .B0(new_new_n472_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n160_), .B(new_new_n124_), .Y(new_new_n479_));
  OAI210     g457(.A0(new_new_n479_), .A1(new_new_n462_), .B0(i_2_), .Y(new_new_n480_));
  INV        g458(.A(new_new_n156_), .Y(new_new_n481_));
  NO3        g459(.A(new_new_n361_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n482_));
  AOI210     g460(.A0(new_new_n481_), .A1(new_new_n86_), .B0(new_new_n482_), .Y(new_new_n483_));
  AOI210     g461(.A0(new_new_n483_), .A1(new_new_n480_), .B0(new_new_n161_), .Y(new_new_n484_));
  OA210      g462(.A0(new_new_n362_), .A1(new_new_n125_), .B0(i_13_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n147_), .B(new_new_n340_), .Y(new_new_n486_));
  NO2        g464(.A(new_new_n486_), .B(new_new_n230_), .Y(new_new_n487_));
  AOI210     g465(.A0(new_new_n166_), .A1(new_new_n145_), .B0(new_new_n305_), .Y(new_new_n488_));
  OAI210     g466(.A0(new_new_n488_), .A1(new_new_n176_), .B0(new_new_n254_), .Y(new_new_n489_));
  NO2        g467(.A(new_new_n102_), .B(new_new_n44_), .Y(new_new_n490_));
  INV        g468(.A(new_new_n209_), .Y(new_new_n491_));
  NA4        g469(.A(new_new_n491_), .B(new_new_n210_), .C(new_new_n123_), .D(new_new_n42_), .Y(new_new_n492_));
  OAI210     g470(.A0(new_new_n492_), .A1(new_new_n490_), .B0(new_new_n489_), .Y(new_new_n493_));
  NO4        g471(.A(new_new_n493_), .B(new_new_n487_), .C(new_new_n485_), .D(new_new_n484_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n328_), .B(new_new_n28_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n461_), .B(new_new_n207_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n496_), .B(new_new_n495_), .Y(new_new_n497_));
  NO2        g475(.A(new_new_n61_), .B(i_12_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n498_), .B(new_new_n125_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n499_), .B(new_new_n340_), .Y(new_new_n500_));
  AOI220     g478(.A0(new_new_n500_), .A1(new_new_n36_), .B0(new_new_n497_), .B1(new_new_n46_), .Y(new_new_n501_));
  NA4        g479(.A(new_new_n501_), .B(new_new_n494_), .C(new_new_n478_), .D(new_new_n468_), .Y(zz06));
  NO2        g480(.A(new_new_n171_), .B(new_new_n289_), .Y(new_new_n503_));
  INV        g481(.A(new_new_n217_), .Y(new_new_n504_));
  OR2        g482(.A(new_new_n504_), .B(i_12_), .Y(new_new_n505_));
  NA2        g483(.A(new_new_n329_), .B(new_new_n62_), .Y(new_new_n506_));
  INV        g484(.A(new_new_n506_), .Y(new_new_n507_));
  NA2        g485(.A(new_new_n507_), .B(new_new_n72_), .Y(new_new_n508_));
  INV        g486(.A(new_new_n216_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n74_), .B(new_new_n130_), .Y(new_new_n510_));
  INV        g488(.A(new_new_n123_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n511_), .B(new_new_n46_), .Y(new_new_n512_));
  AOI210     g490(.A0(new_new_n512_), .A1(new_new_n510_), .B0(new_new_n509_), .Y(new_new_n513_));
  NO2        g491(.A(new_new_n188_), .B(i_9_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n514_), .B(new_new_n498_), .Y(new_new_n515_));
  AOI210     g493(.A0(new_new_n515_), .A1(new_new_n303_), .B0(new_new_n158_), .Y(new_new_n516_));
  NAi32      g494(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n438_), .B(new_new_n517_), .Y(new_new_n518_));
  OR3        g496(.A(new_new_n518_), .B(new_new_n516_), .C(new_new_n513_), .Y(new_new_n519_));
  NO2        g497(.A(new_new_n421_), .B(i_2_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n521_));
  NO2        g499(.A(new_new_n521_), .B(new_new_n249_), .Y(new_new_n522_));
  NA2        g500(.A(new_new_n522_), .B(new_new_n520_), .Y(new_new_n523_));
  BUFFER     g501(.A(new_new_n362_), .Y(new_new_n524_));
  NA3        g502(.A(new_new_n524_), .B(new_new_n144_), .C(new_new_n68_), .Y(new_new_n525_));
  AO210      g503(.A0(new_new_n295_), .A1(new_new_n465_), .B0(new_new_n36_), .Y(new_new_n526_));
  NA3        g504(.A(new_new_n526_), .B(new_new_n525_), .C(new_new_n523_), .Y(new_new_n527_));
  NO2        g505(.A(i_6_), .B(i_11_), .Y(new_new_n528_));
  AOI220     g506(.A0(new_new_n528_), .A1(new_new_n323_), .B0(new_new_n503_), .B1(new_new_n434_), .Y(new_new_n529_));
  NA3        g507(.A(new_new_n230_), .B(new_new_n181_), .C(new_new_n144_), .Y(new_new_n530_));
  NA2        g508(.A(new_new_n244_), .B(new_new_n69_), .Y(new_new_n531_));
  NA4        g509(.A(new_new_n531_), .B(new_new_n530_), .C(new_new_n529_), .D(new_new_n348_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n268_), .B(new_new_n266_), .Y(new_new_n533_));
  NO2        g511(.A(new_new_n356_), .B(new_new_n102_), .Y(new_new_n534_));
  OAI210     g512(.A0(new_new_n534_), .A1(new_new_n111_), .B0(new_new_n248_), .Y(new_new_n535_));
  INV        g513(.A(new_new_n331_), .Y(new_new_n536_));
  NA3        g514(.A(new_new_n536_), .B(new_new_n216_), .C(i_7_), .Y(new_new_n537_));
  NA3        g515(.A(new_new_n537_), .B(new_new_n535_), .C(new_new_n533_), .Y(new_new_n538_));
  NO4        g516(.A(new_new_n538_), .B(new_new_n532_), .C(new_new_n527_), .D(new_new_n519_), .Y(new_new_n539_));
  NA4        g517(.A(new_new_n539_), .B(new_new_n508_), .C(new_new_n505_), .D(new_new_n238_), .Y(zz03));
  NA2        g518(.A(i_12_), .B(i_10_), .Y(new_new_n541_));
  NO2        g519(.A(i_11_), .B(new_new_n179_), .Y(new_new_n542_));
  NA3        g520(.A(new_new_n530_), .B(new_new_n348_), .C(new_new_n229_), .Y(new_new_n543_));
  NA2        g521(.A(new_new_n543_), .B(new_new_n40_), .Y(new_new_n544_));
  NOi21      g522(.An(new_new_n96_), .B(new_new_n474_), .Y(new_new_n545_));
  NO3        g523(.A(new_new_n369_), .B(new_new_n272_), .C(new_new_n130_), .Y(new_new_n546_));
  AN2        g524(.A(new_new_n270_), .B(new_new_n55_), .Y(new_new_n547_));
  NO3        g525(.A(new_new_n547_), .B(new_new_n546_), .C(new_new_n545_), .Y(new_new_n548_));
  AOI210     g526(.A0(new_new_n548_), .A1(new_new_n544_), .B0(new_new_n48_), .Y(new_new_n549_));
  NO4        g527(.A(new_new_n234_), .B(new_new_n240_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n550_));
  NA2        g528(.A(new_new_n158_), .B(new_new_n326_), .Y(new_new_n551_));
  NOi31      g529(.An(new_new_n551_), .B(new_new_n550_), .C(new_new_n39_), .Y(new_new_n552_));
  NO2        g530(.A(new_new_n552_), .B(new_new_n62_), .Y(new_new_n553_));
  NOi21      g531(.An(i_5_), .B(i_9_), .Y(new_new_n554_));
  NA2        g532(.A(new_new_n554_), .B(new_new_n265_), .Y(new_new_n555_));
  BUFFER     g533(.A(new_new_n202_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n556_), .B(new_new_n285_), .Y(new_new_n557_));
  NO2        g535(.A(new_new_n557_), .B(new_new_n555_), .Y(new_new_n558_));
  NO3        g536(.A(new_new_n558_), .B(new_new_n553_), .C(new_new_n549_), .Y(new_new_n559_));
  NA2        g537(.A(new_new_n327_), .B(i_0_), .Y(new_new_n560_));
  NO4        g538(.A(new_new_n330_), .B(new_new_n168_), .C(new_new_n252_), .D(new_new_n249_), .Y(new_new_n561_));
  NA2        g539(.A(new_new_n561_), .B(i_11_), .Y(new_new_n562_));
  NA2        g540(.A(new_new_n461_), .B(new_new_n217_), .Y(new_new_n563_));
  AOI210     g541(.A0(new_new_n287_), .A1(new_new_n86_), .B0(new_new_n57_), .Y(new_new_n564_));
  NO2        g542(.A(new_new_n564_), .B(new_new_n563_), .Y(new_new_n565_));
  NO2        g543(.A(new_new_n190_), .B(new_new_n148_), .Y(new_new_n566_));
  NA2        g544(.A(i_0_), .B(i_10_), .Y(new_new_n567_));
  INV        g545(.A(new_new_n309_), .Y(new_new_n568_));
  NO4        g546(.A(new_new_n114_), .B(new_new_n57_), .C(new_new_n397_), .D(i_5_), .Y(new_new_n569_));
  AO220      g547(.A0(new_new_n569_), .A1(new_new_n568_), .B0(new_new_n566_), .B1(i_6_), .Y(new_new_n570_));
  NO2        g548(.A(new_new_n570_), .B(new_new_n565_), .Y(new_new_n571_));
  NA2        g549(.A(new_new_n571_), .B(new_new_n562_), .Y(new_new_n572_));
  NO2        g550(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n573_));
  NA2        g551(.A(i_11_), .B(i_9_), .Y(new_new_n574_));
  NO3        g552(.A(i_12_), .B(new_new_n574_), .C(new_new_n347_), .Y(new_new_n575_));
  AN2        g553(.A(new_new_n575_), .B(new_new_n573_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n243_), .B(new_new_n157_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n577_), .B(new_new_n152_), .Y(new_new_n578_));
  NO2        g556(.A(new_new_n574_), .B(new_new_n72_), .Y(new_new_n579_));
  INV        g557(.A(new_new_n247_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n580_), .B(new_new_n555_), .Y(new_new_n581_));
  NO3        g559(.A(new_new_n581_), .B(new_new_n578_), .C(new_new_n576_), .Y(new_new_n582_));
  NA2        g560(.A(new_new_n388_), .B(new_new_n120_), .Y(new_new_n583_));
  NO2        g561(.A(i_6_), .B(new_new_n583_), .Y(new_new_n584_));
  NA2        g562(.A(new_new_n155_), .B(new_new_n103_), .Y(new_new_n585_));
  INV        g563(.A(new_new_n584_), .Y(new_new_n586_));
  INV        g564(.A(new_new_n215_), .Y(new_new_n587_));
  NA2        g565(.A(new_new_n586_), .B(new_new_n582_), .Y(new_new_n588_));
  NO2        g566(.A(new_new_n541_), .B(new_new_n214_), .Y(new_new_n589_));
  NA2        g567(.A(new_new_n589_), .B(new_new_n579_), .Y(new_new_n590_));
  NA2        g568(.A(new_new_n423_), .B(new_new_n311_), .Y(new_new_n591_));
  NAi21      g569(.An(i_9_), .B(i_5_), .Y(new_new_n592_));
  NO2        g570(.A(new_new_n592_), .B(new_new_n246_), .Y(new_new_n593_));
  NA2        g571(.A(new_new_n593_), .B(new_new_n362_), .Y(new_new_n594_));
  OAI220     g572(.A0(new_new_n594_), .A1(new_new_n85_), .B0(new_new_n591_), .B1(new_new_n156_), .Y(new_new_n595_));
  NO2        g573(.A(new_new_n595_), .B(new_new_n307_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n596_), .B(new_new_n590_), .Y(new_new_n597_));
  NO3        g575(.A(new_new_n597_), .B(new_new_n588_), .C(new_new_n572_), .Y(new_new_n598_));
  AOI210     g576(.A0(new_new_n506_), .A1(new_new_n414_), .B0(new_new_n585_), .Y(new_new_n599_));
  INV        g577(.A(new_new_n599_), .Y(new_new_n600_));
  OAI210     g578(.A0(new_new_n185_), .A1(i_9_), .B0(new_new_n177_), .Y(new_new_n601_));
  AOI210     g579(.A0(new_new_n601_), .A1(new_new_n560_), .B0(new_new_n148_), .Y(new_new_n602_));
  INV        g580(.A(new_new_n602_), .Y(new_new_n603_));
  NA2        g581(.A(new_new_n603_), .B(new_new_n600_), .Y(new_new_n604_));
  NO3        g582(.A(new_new_n567_), .B(new_new_n554_), .C(new_new_n160_), .Y(new_new_n605_));
  AOI220     g583(.A0(new_new_n605_), .A1(i_11_), .B0(new_new_n325_), .B1(new_new_n74_), .Y(new_new_n606_));
  NO3        g584(.A(new_new_n167_), .B(new_new_n240_), .C(i_0_), .Y(new_new_n607_));
  OAI210     g585(.A0(new_new_n607_), .A1(new_new_n75_), .B0(i_13_), .Y(new_new_n608_));
  NA2        g586(.A(new_new_n608_), .B(new_new_n606_), .Y(new_new_n609_));
  NA3        g587(.A(new_new_n242_), .B(new_new_n155_), .C(new_new_n154_), .Y(new_new_n610_));
  INV        g588(.A(new_new_n610_), .Y(new_new_n611_));
  NO3        g589(.A(new_new_n574_), .B(new_new_n170_), .C(new_new_n160_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n612_), .B(new_new_n611_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n613_), .B(new_new_n288_), .Y(new_new_n614_));
  NO2        g592(.A(new_new_n85_), .B(i_5_), .Y(new_new_n615_));
  NA3        g593(.A(new_new_n542_), .B(new_new_n109_), .C(new_new_n123_), .Y(new_new_n616_));
  INV        g594(.A(new_new_n616_), .Y(new_new_n617_));
  NA2        g595(.A(new_new_n617_), .B(new_new_n615_), .Y(new_new_n618_));
  NAi21      g596(.An(new_new_n183_), .B(new_new_n184_), .Y(new_new_n619_));
  NO4        g597(.A(new_new_n182_), .B(new_new_n167_), .C(i_0_), .D(i_12_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n620_), .B(new_new_n619_), .Y(new_new_n621_));
  NA2        g599(.A(new_new_n621_), .B(new_new_n618_), .Y(new_new_n622_));
  NO4        g600(.A(new_new_n622_), .B(new_new_n614_), .C(new_new_n609_), .D(new_new_n604_), .Y(new_new_n623_));
  NA2        g601(.A(new_new_n520_), .B(new_new_n37_), .Y(new_new_n624_));
  NA2        g602(.A(new_new_n624_), .B(new_new_n355_), .Y(new_new_n625_));
  NA2        g603(.A(new_new_n625_), .B(new_new_n165_), .Y(new_new_n626_));
  NAi31      g604(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n627_));
  AOI210     g605(.A0(new_new_n116_), .A1(new_new_n69_), .B0(new_new_n627_), .Y(new_new_n628_));
  AOI210     g606(.A0(new_new_n628_), .A1(new_new_n48_), .B0(new_new_n561_), .Y(new_new_n629_));
  AOI210     g607(.A0(new_new_n629_), .A1(new_new_n626_), .B0(new_new_n72_), .Y(new_new_n630_));
  INV        g608(.A(new_new_n237_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n631_), .B(new_new_n469_), .Y(new_new_n632_));
  NO3        g610(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n633_));
  OAI210     g611(.A0(new_new_n587_), .A1(new_new_n211_), .B0(new_new_n633_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n634_), .B(new_new_n443_), .Y(new_new_n635_));
  NO3        g613(.A(new_new_n635_), .B(new_new_n632_), .C(new_new_n630_), .Y(new_new_n636_));
  NA4        g614(.A(new_new_n636_), .B(new_new_n623_), .C(new_new_n598_), .D(new_new_n559_), .Y(zz04));
  INV        g615(.A(new_new_n422_), .Y(new_new_n640_));
  INV        g616(.A(i_6_), .Y(new_new_n641_));
endmodule


