// Benchmark "top" written by ABC on Fri Jun 21 17:49:22 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n133_, new_new_n134_, new_new_n135_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n1002_, new_new_n1003_,
    new_new_n1004_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NO2        g028(.A(new_new_n47_), .B(new_new_n46_), .Y(new_new_n51_));
  NA2        g029(.A(i_0_), .B(i_2_), .Y(new_new_n52_));
  NA2        g030(.A(i_7_), .B(i_9_), .Y(new_new_n53_));
  NO2        g031(.A(new_new_n53_), .B(new_new_n52_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n51_), .B(new_new_n45_), .Y(new_new_n55_));
  NA3        g033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  OAI210     g036(.A0(new_new_n58_), .A1(new_new_n57_), .B0(new_new_n56_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g039(.A(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NA3        g041(.A(new_new_n63_), .B(new_new_n61_), .C(new_new_n31_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n64_), .B(new_new_n60_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n50_), .B(i_2_), .Y(new_new_n66_));
  AOI210     g044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n67_));
  NA2        g045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n74_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n75_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  NO2        g055(.A(i_3_), .B(i_9_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_7_), .Y(new_new_n79_));
  INV        g057(.A(i_6_), .Y(new_new_n80_));
  OR4        g058(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n81_));
  INV        g059(.A(new_new_n81_), .Y(new_new_n82_));
  NO2        g060(.A(i_2_), .B(i_7_), .Y(new_new_n83_));
  NAi21      g061(.An(i_6_), .B(i_10_), .Y(new_new_n84_));
  NA2        g062(.A(i_6_), .B(i_9_), .Y(new_new_n85_));
  AOI210     g063(.A0(new_new_n85_), .A1(new_new_n84_), .B0(new_new_n62_), .Y(new_new_n86_));
  NA2        g064(.A(i_2_), .B(i_6_), .Y(new_new_n87_));
  INV        g065(.A(new_new_n86_), .Y(new_new_n88_));
  NO2        g066(.A(new_new_n88_), .B(new_new_n77_), .Y(new_new_n89_));
  AN3        g067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n90_));
  NAi21      g068(.An(i_6_), .B(i_11_), .Y(new_new_n91_));
  NO2        g069(.A(i_5_), .B(i_8_), .Y(new_new_n92_));
  NOi21      g070(.An(new_new_n92_), .B(new_new_n91_), .Y(new_new_n93_));
  AOI220     g071(.A0(new_new_n93_), .A1(new_new_n61_), .B0(new_new_n90_), .B1(new_new_n32_), .Y(new_new_n94_));
  INV        g072(.A(i_7_), .Y(new_new_n95_));
  NA2        g073(.A(new_new_n46_), .B(new_new_n95_), .Y(new_new_n96_));
  NO2        g074(.A(i_0_), .B(i_5_), .Y(new_new_n97_));
  NO2        g075(.A(new_new_n97_), .B(new_new_n80_), .Y(new_new_n98_));
  NA2        g076(.A(i_12_), .B(i_3_), .Y(new_new_n99_));
  INV        g077(.A(new_new_n99_), .Y(new_new_n100_));
  NA3        g078(.A(new_new_n100_), .B(new_new_n98_), .C(new_new_n96_), .Y(new_new_n101_));
  NAi21      g079(.An(i_7_), .B(i_11_), .Y(new_new_n102_));
  NO3        g080(.A(new_new_n102_), .B(new_new_n84_), .C(new_new_n52_), .Y(new_new_n103_));
  AN2        g081(.A(i_2_), .B(i_10_), .Y(new_new_n104_));
  NO2        g082(.A(new_new_n104_), .B(i_7_), .Y(new_new_n105_));
  OR2        g083(.A(new_new_n77_), .B(new_new_n57_), .Y(new_new_n106_));
  NO2        g084(.A(i_8_), .B(new_new_n95_), .Y(new_new_n107_));
  NO3        g085(.A(new_new_n107_), .B(new_new_n106_), .C(new_new_n105_), .Y(new_new_n108_));
  NA2        g086(.A(i_12_), .B(i_7_), .Y(new_new_n109_));
  NO2        g087(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n110_));
  NA2        g088(.A(new_new_n110_), .B(i_0_), .Y(new_new_n111_));
  NA2        g089(.A(i_11_), .B(i_12_), .Y(new_new_n112_));
  OAI210     g090(.A0(new_new_n111_), .A1(new_new_n109_), .B0(new_new_n112_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n113_), .B(new_new_n108_), .Y(new_new_n114_));
  NAi41      g092(.An(new_new_n103_), .B(new_new_n114_), .C(new_new_n101_), .D(new_new_n94_), .Y(new_new_n115_));
  NOi21      g093(.An(i_1_), .B(i_5_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(i_11_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n95_), .B(new_new_n37_), .Y(new_new_n118_));
  NA2        g096(.A(i_7_), .B(new_new_n25_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(new_new_n118_), .Y(new_new_n120_));
  NO2        g098(.A(new_new_n120_), .B(new_new_n46_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n85_), .B(new_new_n84_), .Y(new_new_n122_));
  NAi21      g100(.An(i_3_), .B(i_8_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n61_), .Y(new_new_n124_));
  NOi21      g102(.An(new_new_n124_), .B(new_new_n122_), .Y(new_new_n125_));
  NO2        g103(.A(i_1_), .B(new_new_n80_), .Y(new_new_n126_));
  NO2        g104(.A(i_6_), .B(i_5_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(i_3_), .Y(new_new_n128_));
  AO210      g106(.A0(new_new_n128_), .A1(new_new_n47_), .B0(new_new_n126_), .Y(new_new_n129_));
  OAI220     g107(.A0(new_new_n129_), .A1(new_new_n102_), .B0(new_new_n125_), .B1(new_new_n117_), .Y(new_new_n130_));
  NO3        g108(.A(new_new_n130_), .B(new_new_n115_), .C(new_new_n89_), .Y(new_new_n131_));
  NA3        g109(.A(new_new_n131_), .B(new_new_n76_), .C(new_new_n55_), .Y(mai2));
  NO2        g110(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n133_));
  NA2        g111(.A(i_6_), .B(new_new_n25_), .Y(new_new_n134_));
  NA2        g112(.A(new_new_n134_), .B(new_new_n133_), .Y(new_new_n135_));
  NA4        g113(.A(new_new_n135_), .B(new_new_n74_), .C(new_new_n66_), .D(new_new_n30_), .Y(mai0));
  AN2        g114(.A(i_8_), .B(i_7_), .Y(new_new_n137_));
  NA2        g115(.A(new_new_n137_), .B(i_6_), .Y(new_new_n138_));
  NO2        g116(.A(i_12_), .B(i_13_), .Y(new_new_n139_));
  NAi21      g117(.An(i_5_), .B(i_11_), .Y(new_new_n140_));
  NOi21      g118(.An(new_new_n139_), .B(new_new_n140_), .Y(new_new_n141_));
  NO2        g119(.A(i_0_), .B(i_1_), .Y(new_new_n142_));
  NA2        g120(.A(i_2_), .B(i_3_), .Y(new_new_n143_));
  NO2        g121(.A(new_new_n143_), .B(i_4_), .Y(new_new_n144_));
  NA2        g122(.A(new_new_n144_), .B(new_new_n141_), .Y(new_new_n145_));
  AN2        g123(.A(new_new_n139_), .B(new_new_n78_), .Y(new_new_n146_));
  NA2        g124(.A(i_1_), .B(i_5_), .Y(new_new_n147_));
  NO2        g125(.A(new_new_n70_), .B(new_new_n46_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n36_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n149_), .B(new_new_n147_), .C(i_13_), .Y(new_new_n150_));
  OR2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NO3        g129(.A(new_new_n151_), .B(new_new_n77_), .C(i_13_), .Y(new_new_n152_));
  NAi32      g130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n153_));
  NAi21      g131(.An(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  NOi21      g132(.An(i_4_), .B(i_10_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n40_), .Y(new_new_n156_));
  NO2        g134(.A(i_3_), .B(i_5_), .Y(new_new_n157_));
  NO3        g135(.A(new_new_n70_), .B(i_2_), .C(i_1_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n157_), .Y(new_new_n159_));
  OAI210     g137(.A0(new_new_n159_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n160_), .B(new_new_n150_), .Y(new_new_n161_));
  AOI210     g139(.A0(new_new_n161_), .A1(new_new_n145_), .B0(new_new_n138_), .Y(new_new_n162_));
  NA3        g140(.A(new_new_n70_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n163_));
  NOi21      g141(.An(i_4_), .B(i_9_), .Y(new_new_n164_));
  NOi21      g142(.An(i_11_), .B(i_13_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  BUFFER     g144(.A(new_new_n166_), .Y(new_new_n167_));
  NO2        g145(.A(i_4_), .B(i_5_), .Y(new_new_n168_));
  NAi21      g146(.An(i_12_), .B(i_11_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n169_), .B(i_13_), .Y(new_new_n170_));
  NA2        g148(.A(new_new_n170_), .B(new_new_n78_), .Y(new_new_n171_));
  AOI210     g149(.A0(new_new_n171_), .A1(new_new_n167_), .B0(new_new_n163_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n70_), .B(new_new_n62_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(new_new_n46_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n36_), .B(i_5_), .Y(new_new_n175_));
  NAi31      g153(.An(new_new_n175_), .B(new_new_n146_), .C(i_11_), .Y(new_new_n176_));
  NA2        g154(.A(i_3_), .B(i_5_), .Y(new_new_n177_));
  BUFFER     g155(.A(new_new_n166_), .Y(new_new_n178_));
  AOI210     g156(.A0(new_new_n178_), .A1(new_new_n176_), .B0(new_new_n174_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n70_), .B(i_5_), .Y(new_new_n180_));
  NO2        g158(.A(i_13_), .B(i_10_), .Y(new_new_n181_));
  NA3        g159(.A(new_new_n181_), .B(new_new_n180_), .C(new_new_n44_), .Y(new_new_n182_));
  NO2        g160(.A(i_2_), .B(i_1_), .Y(new_new_n183_));
  NA2        g161(.A(new_new_n183_), .B(i_3_), .Y(new_new_n184_));
  NAi21      g162(.An(i_4_), .B(i_12_), .Y(new_new_n185_));
  NO3        g163(.A(new_new_n185_), .B(new_new_n184_), .C(new_new_n182_), .Y(new_new_n186_));
  NO3        g164(.A(new_new_n186_), .B(new_new_n179_), .C(new_new_n172_), .Y(new_new_n187_));
  INV        g165(.A(i_8_), .Y(new_new_n188_));
  NA2        g166(.A(i_8_), .B(i_6_), .Y(new_new_n189_));
  NO3        g167(.A(i_3_), .B(new_new_n80_), .C(new_new_n48_), .Y(new_new_n190_));
  NA2        g168(.A(new_new_n190_), .B(new_new_n107_), .Y(new_new_n191_));
  NO3        g169(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n192_));
  NA3        g170(.A(new_new_n192_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n193_));
  NO3        g171(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n194_));
  OAI210     g172(.A0(new_new_n90_), .A1(i_12_), .B0(new_new_n194_), .Y(new_new_n195_));
  AOI210     g173(.A0(new_new_n195_), .A1(new_new_n193_), .B0(new_new_n191_), .Y(new_new_n196_));
  NO2        g174(.A(i_3_), .B(i_8_), .Y(new_new_n197_));
  NO3        g175(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n198_));
  NA3        g176(.A(new_new_n198_), .B(new_new_n197_), .C(new_new_n40_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n97_), .B(new_new_n57_), .Y(new_new_n200_));
  NO2        g178(.A(i_13_), .B(i_9_), .Y(new_new_n201_));
  NA3        g179(.A(new_new_n201_), .B(i_6_), .C(new_new_n188_), .Y(new_new_n202_));
  NAi21      g180(.An(i_12_), .B(i_3_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n44_), .B(i_5_), .Y(new_new_n204_));
  NO3        g182(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n205_));
  NA2        g183(.A(new_new_n205_), .B(i_10_), .Y(new_new_n206_));
  OAI220     g184(.A0(new_new_n206_), .A1(new_new_n202_), .B0(new_new_n57_), .B1(new_new_n199_), .Y(new_new_n207_));
  AOI210     g185(.A0(new_new_n207_), .A1(i_7_), .B0(new_new_n196_), .Y(new_new_n208_));
  OAI220     g186(.A0(new_new_n208_), .A1(i_4_), .B0(new_new_n189_), .B1(new_new_n187_), .Y(new_new_n209_));
  NAi21      g187(.An(i_12_), .B(i_7_), .Y(new_new_n210_));
  NA3        g188(.A(i_13_), .B(new_new_n188_), .C(i_10_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n211_), .B(new_new_n210_), .Y(new_new_n212_));
  NA2        g190(.A(i_0_), .B(i_5_), .Y(new_new_n213_));
  OAI220     g191(.A0(new_new_n80_), .A1(new_new_n184_), .B0(new_new_n174_), .B1(new_new_n128_), .Y(new_new_n214_));
  NAi31      g192(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n36_), .B(i_13_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n46_), .B(new_new_n62_), .Y(new_new_n217_));
  NA2        g195(.A(new_new_n217_), .B(new_new_n216_), .Y(new_new_n218_));
  INV        g196(.A(i_13_), .Y(new_new_n219_));
  NO2        g197(.A(i_12_), .B(new_new_n219_), .Y(new_new_n220_));
  NA3        g198(.A(new_new_n220_), .B(new_new_n192_), .C(new_new_n190_), .Y(new_new_n221_));
  OAI210     g199(.A0(new_new_n218_), .A1(new_new_n215_), .B0(new_new_n221_), .Y(new_new_n222_));
  AOI220     g200(.A0(new_new_n222_), .A1(new_new_n137_), .B0(new_new_n214_), .B1(new_new_n212_), .Y(new_new_n223_));
  NO2        g201(.A(i_12_), .B(new_new_n37_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n177_), .B(i_4_), .Y(new_new_n225_));
  NA2        g203(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n226_));
  OR2        g204(.A(i_8_), .B(i_7_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(new_new_n80_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n52_), .B(i_1_), .Y(new_new_n229_));
  INV        g207(.A(i_12_), .Y(new_new_n230_));
  NO3        g208(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n231_));
  NA2        g209(.A(i_2_), .B(i_1_), .Y(new_new_n232_));
  NO3        g210(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n233_));
  NAi21      g211(.An(i_4_), .B(i_3_), .Y(new_new_n234_));
  NO2        g212(.A(new_new_n234_), .B(new_new_n72_), .Y(new_new_n235_));
  NO2        g213(.A(i_0_), .B(i_6_), .Y(new_new_n236_));
  NOi41      g214(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n238_));
  NO2        g216(.A(new_new_n232_), .B(new_new_n177_), .Y(new_new_n239_));
  NAi21      g217(.An(new_new_n238_), .B(new_new_n239_), .Y(new_new_n240_));
  NO2        g218(.A(i_11_), .B(new_new_n219_), .Y(new_new_n241_));
  NOi21      g219(.An(i_1_), .B(i_6_), .Y(new_new_n242_));
  NAi21      g220(.An(i_3_), .B(i_7_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n244_));
  NO2        g222(.A(i_12_), .B(i_3_), .Y(new_new_n245_));
  NA3        g223(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n246_));
  INV        g224(.A(new_new_n138_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n230_), .B(i_13_), .Y(new_new_n248_));
  NO2        g226(.A(new_new_n248_), .B(new_new_n72_), .Y(new_new_n249_));
  NA2        g227(.A(new_new_n249_), .B(new_new_n247_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n227_), .B(new_new_n37_), .Y(new_new_n251_));
  NA2        g229(.A(i_12_), .B(i_6_), .Y(new_new_n252_));
  OR2        g230(.A(i_13_), .B(i_9_), .Y(new_new_n253_));
  NO3        g231(.A(new_new_n253_), .B(new_new_n252_), .C(new_new_n48_), .Y(new_new_n254_));
  NO2        g232(.A(new_new_n234_), .B(i_2_), .Y(new_new_n255_));
  NA3        g233(.A(new_new_n255_), .B(new_new_n254_), .C(new_new_n44_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n241_), .B(i_9_), .Y(new_new_n257_));
  OAI210     g235(.A0(new_new_n62_), .A1(new_new_n257_), .B0(new_new_n256_), .Y(new_new_n258_));
  NO3        g236(.A(i_11_), .B(new_new_n219_), .C(new_new_n25_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n243_), .B(i_8_), .Y(new_new_n260_));
  NO2        g238(.A(i_6_), .B(new_new_n48_), .Y(new_new_n261_));
  NA3        g239(.A(new_new_n261_), .B(new_new_n260_), .C(new_new_n259_), .Y(new_new_n262_));
  NO3        g240(.A(new_new_n26_), .B(new_new_n80_), .C(i_5_), .Y(new_new_n263_));
  NA3        g241(.A(new_new_n263_), .B(new_new_n251_), .C(new_new_n220_), .Y(new_new_n264_));
  AOI210     g242(.A0(new_new_n264_), .A1(new_new_n262_), .B0(i_1_), .Y(new_new_n265_));
  AOI210     g243(.A0(new_new_n258_), .A1(new_new_n251_), .B0(new_new_n265_), .Y(new_new_n266_));
  NA4        g244(.A(new_new_n266_), .B(new_new_n250_), .C(new_new_n240_), .D(new_new_n223_), .Y(new_new_n267_));
  NO3        g245(.A(i_12_), .B(new_new_n219_), .C(new_new_n37_), .Y(new_new_n268_));
  INV        g246(.A(new_new_n268_), .Y(new_new_n269_));
  NA2        g247(.A(i_8_), .B(new_new_n95_), .Y(new_new_n270_));
  NO3        g248(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n271_));
  AOI220     g249(.A0(new_new_n271_), .A1(new_new_n190_), .B0(new_new_n157_), .B1(new_new_n229_), .Y(new_new_n272_));
  NO2        g250(.A(new_new_n272_), .B(new_new_n270_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n232_), .B(i_0_), .Y(new_new_n274_));
  AOI220     g252(.A0(new_new_n274_), .A1(i_8_), .B0(i_1_), .B1(new_new_n137_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n261_), .B(new_new_n26_), .Y(new_new_n276_));
  NO2        g254(.A(new_new_n276_), .B(new_new_n275_), .Y(new_new_n277_));
  NA2        g255(.A(i_0_), .B(i_1_), .Y(new_new_n278_));
  NO2        g256(.A(new_new_n278_), .B(i_2_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n58_), .B(i_6_), .Y(new_new_n280_));
  NA2        g258(.A(new_new_n280_), .B(new_new_n279_), .Y(new_new_n281_));
  OAI210     g259(.A0(new_new_n159_), .A1(new_new_n138_), .B0(new_new_n281_), .Y(new_new_n282_));
  NO3        g260(.A(new_new_n282_), .B(new_new_n277_), .C(new_new_n273_), .Y(new_new_n283_));
  NO2        g261(.A(i_3_), .B(i_10_), .Y(new_new_n284_));
  NA3        g262(.A(new_new_n284_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n285_));
  NO2        g263(.A(i_2_), .B(new_new_n95_), .Y(new_new_n286_));
  NA2        g264(.A(i_1_), .B(new_new_n36_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n287_), .B(i_8_), .Y(new_new_n288_));
  INV        g266(.A(new_new_n288_), .Y(new_new_n289_));
  AN2        g267(.A(i_3_), .B(i_10_), .Y(new_new_n290_));
  NA3        g268(.A(new_new_n290_), .B(new_new_n192_), .C(new_new_n170_), .Y(new_new_n291_));
  NO2        g269(.A(i_5_), .B(new_new_n37_), .Y(new_new_n292_));
  NO2        g270(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n293_));
  OR2        g271(.A(new_new_n289_), .B(new_new_n285_), .Y(new_new_n294_));
  OAI220     g272(.A0(new_new_n294_), .A1(i_6_), .B0(new_new_n283_), .B1(new_new_n269_), .Y(new_new_n295_));
  NO4        g273(.A(new_new_n295_), .B(new_new_n267_), .C(new_new_n209_), .D(new_new_n162_), .Y(new_new_n296_));
  NO3        g274(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n297_));
  NO2        g275(.A(new_new_n58_), .B(new_new_n80_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n274_), .B(new_new_n298_), .Y(new_new_n299_));
  NO3        g277(.A(i_6_), .B(new_new_n188_), .C(i_7_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n300_), .B(new_new_n192_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n301_), .B(new_new_n299_), .Y(new_new_n302_));
  NO2        g280(.A(i_2_), .B(i_3_), .Y(new_new_n303_));
  OR2        g281(.A(i_0_), .B(i_5_), .Y(new_new_n304_));
  NA3        g282(.A(new_new_n228_), .B(new_new_n303_), .C(i_1_), .Y(new_new_n305_));
  NA3        g283(.A(new_new_n274_), .B(new_new_n157_), .C(new_new_n107_), .Y(new_new_n306_));
  NAi21      g284(.An(i_8_), .B(i_7_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n307_), .B(i_6_), .Y(new_new_n308_));
  NO2        g286(.A(new_new_n151_), .B(new_new_n46_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n309_), .B(new_new_n308_), .Y(new_new_n310_));
  NA3        g288(.A(new_new_n310_), .B(new_new_n306_), .C(new_new_n305_), .Y(new_new_n311_));
  OAI210     g289(.A0(new_new_n311_), .A1(new_new_n302_), .B0(i_4_), .Y(new_new_n312_));
  NO2        g290(.A(i_12_), .B(i_10_), .Y(new_new_n313_));
  NOi21      g291(.An(i_5_), .B(i_0_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n287_), .B(new_new_n123_), .Y(new_new_n315_));
  NA4        g293(.A(new_new_n79_), .B(new_new_n36_), .C(new_new_n80_), .D(i_8_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n315_), .B(new_new_n313_), .Y(new_new_n317_));
  NO2        g295(.A(i_6_), .B(i_8_), .Y(new_new_n318_));
  NOi21      g296(.An(i_0_), .B(i_2_), .Y(new_new_n319_));
  AN2        g297(.A(new_new_n319_), .B(new_new_n318_), .Y(new_new_n320_));
  NO2        g298(.A(i_1_), .B(i_7_), .Y(new_new_n321_));
  AO220      g299(.A0(new_new_n321_), .A1(new_new_n320_), .B0(new_new_n308_), .B1(new_new_n229_), .Y(new_new_n322_));
  NA2        g300(.A(new_new_n322_), .B(i_4_), .Y(new_new_n323_));
  NA3        g301(.A(new_new_n323_), .B(new_new_n317_), .C(new_new_n312_), .Y(new_new_n324_));
  NO3        g302(.A(new_new_n227_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n325_));
  NO3        g303(.A(new_new_n307_), .B(i_2_), .C(i_1_), .Y(new_new_n326_));
  OAI210     g304(.A0(new_new_n326_), .A1(new_new_n325_), .B0(i_6_), .Y(new_new_n327_));
  NA2        g305(.A(new_new_n242_), .B(new_new_n286_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n328_), .B(new_new_n327_), .Y(new_new_n329_));
  NA2        g307(.A(new_new_n329_), .B(i_3_), .Y(new_new_n330_));
  INV        g308(.A(new_new_n79_), .Y(new_new_n331_));
  INV        g309(.A(new_new_n278_), .Y(new_new_n332_));
  NA2        g310(.A(new_new_n332_), .B(new_new_n127_), .Y(new_new_n333_));
  AOI210     g311(.A0(new_new_n87_), .A1(new_new_n333_), .B0(new_new_n331_), .Y(new_new_n334_));
  INV        g312(.A(i_9_), .Y(new_new_n335_));
  NA2        g313(.A(new_new_n335_), .B(new_new_n200_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n336_), .B(new_new_n46_), .Y(new_new_n337_));
  NO3        g315(.A(new_new_n337_), .B(new_new_n334_), .C(new_new_n277_), .Y(new_new_n338_));
  AOI210     g316(.A0(new_new_n338_), .A1(new_new_n330_), .B0(new_new_n156_), .Y(new_new_n339_));
  AOI210     g317(.A0(new_new_n324_), .A1(new_new_n297_), .B0(new_new_n339_), .Y(new_new_n340_));
  NOi32      g318(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n341_));
  INV        g319(.A(new_new_n341_), .Y(new_new_n342_));
  NAi21      g320(.An(i_0_), .B(i_6_), .Y(new_new_n343_));
  NAi21      g321(.An(i_1_), .B(i_5_), .Y(new_new_n344_));
  NA2        g322(.A(new_new_n344_), .B(new_new_n343_), .Y(new_new_n345_));
  NA2        g323(.A(new_new_n345_), .B(new_new_n25_), .Y(new_new_n346_));
  OAI210     g324(.A0(new_new_n346_), .A1(new_new_n153_), .B0(new_new_n238_), .Y(new_new_n347_));
  NAi41      g325(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n348_));
  OAI220     g326(.A0(new_new_n348_), .A1(new_new_n344_), .B0(new_new_n215_), .B1(new_new_n153_), .Y(new_new_n349_));
  AOI210     g327(.A0(new_new_n348_), .A1(new_new_n153_), .B0(new_new_n151_), .Y(new_new_n350_));
  NOi32      g328(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n351_));
  NAi21      g329(.An(i_6_), .B(i_1_), .Y(new_new_n352_));
  NA3        g330(.A(new_new_n352_), .B(new_new_n351_), .C(new_new_n46_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n353_), .B(i_0_), .Y(new_new_n354_));
  OR3        g332(.A(new_new_n354_), .B(new_new_n350_), .C(new_new_n349_), .Y(new_new_n355_));
  NO2        g333(.A(i_1_), .B(new_new_n95_), .Y(new_new_n356_));
  NAi21      g334(.An(i_3_), .B(i_4_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n357_), .B(i_9_), .Y(new_new_n358_));
  AN2        g336(.A(i_6_), .B(i_7_), .Y(new_new_n359_));
  NA2        g337(.A(i_2_), .B(i_7_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n357_), .B(i_10_), .Y(new_new_n361_));
  NA3        g339(.A(new_new_n361_), .B(new_new_n360_), .C(new_new_n236_), .Y(new_new_n362_));
  INV        g340(.A(new_new_n362_), .Y(new_new_n363_));
  AOI210     g341(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n364_));
  AOI220     g342(.A0(new_new_n361_), .A1(new_new_n321_), .B0(new_new_n231_), .B1(new_new_n183_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n365_), .B(i_5_), .Y(new_new_n366_));
  NO4        g344(.A(new_new_n366_), .B(new_new_n363_), .C(new_new_n355_), .D(new_new_n347_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n367_), .B(new_new_n342_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n58_), .B(new_new_n25_), .Y(new_new_n369_));
  AN2        g347(.A(i_12_), .B(i_5_), .Y(new_new_n370_));
  NA2        g348(.A(i_3_), .B(new_new_n370_), .Y(new_new_n371_));
  NO2        g349(.A(i_11_), .B(i_6_), .Y(new_new_n372_));
  NA3        g350(.A(new_new_n372_), .B(new_new_n309_), .C(new_new_n219_), .Y(new_new_n373_));
  NO2        g351(.A(new_new_n373_), .B(new_new_n371_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n234_), .B(i_5_), .Y(new_new_n375_));
  NO2        g353(.A(i_5_), .B(i_10_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n139_), .B(new_new_n45_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n377_), .B(new_new_n234_), .Y(new_new_n378_));
  OAI210     g356(.A0(new_new_n378_), .A1(new_new_n374_), .B0(new_new_n369_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n380_));
  NA2        g358(.A(new_new_n374_), .B(new_new_n380_), .Y(new_new_n381_));
  NO3        g359(.A(new_new_n80_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n382_));
  INV        g360(.A(new_new_n284_), .Y(new_new_n383_));
  NO2        g361(.A(i_11_), .B(i_12_), .Y(new_new_n384_));
  NA2        g362(.A(new_new_n384_), .B(new_new_n36_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n383_), .B(new_new_n385_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n376_), .B(new_new_n230_), .Y(new_new_n387_));
  NA2        g365(.A(i_4_), .B(i_11_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n388_), .B(new_new_n215_), .Y(new_new_n389_));
  NAi21      g367(.An(i_13_), .B(i_0_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n390_), .B(new_new_n232_), .Y(new_new_n391_));
  OAI210     g369(.A0(new_new_n389_), .A1(new_new_n386_), .B0(new_new_n391_), .Y(new_new_n392_));
  NA3        g370(.A(new_new_n392_), .B(new_new_n381_), .C(new_new_n379_), .Y(new_new_n393_));
  NO3        g371(.A(i_1_), .B(i_12_), .C(new_new_n80_), .Y(new_new_n394_));
  NO2        g372(.A(i_0_), .B(i_11_), .Y(new_new_n395_));
  AN2        g373(.A(i_1_), .B(i_6_), .Y(new_new_n396_));
  NOi21      g374(.An(i_2_), .B(i_12_), .Y(new_new_n397_));
  NA2        g375(.A(new_new_n397_), .B(new_new_n396_), .Y(new_new_n398_));
  INV        g376(.A(new_new_n398_), .Y(new_new_n399_));
  NA2        g377(.A(new_new_n137_), .B(i_9_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n400_), .B(i_4_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n399_), .B(new_new_n401_), .Y(new_new_n402_));
  OR2        g380(.A(i_13_), .B(i_10_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n166_), .B(new_new_n118_), .Y(new_new_n404_));
  BUFFER     g382(.A(new_new_n211_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n95_), .B(new_new_n25_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n268_), .B(new_new_n406_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n261_), .B(new_new_n205_), .Y(new_new_n408_));
  OAI220     g386(.A0(new_new_n408_), .A1(new_new_n405_), .B0(new_new_n407_), .B1(new_new_n97_), .Y(new_new_n409_));
  INV        g387(.A(new_new_n409_), .Y(new_new_n410_));
  AOI210     g388(.A0(new_new_n410_), .A1(new_new_n402_), .B0(new_new_n26_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n306_), .B(new_new_n305_), .Y(new_new_n412_));
  AOI220     g390(.A0(new_new_n280_), .A1(new_new_n271_), .B0(new_new_n274_), .B1(new_new_n298_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n413_), .B(i_5_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n177_), .B(new_new_n80_), .Y(new_new_n415_));
  AOI220     g393(.A0(new_new_n415_), .A1(new_new_n279_), .B0(new_new_n263_), .B1(new_new_n205_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n416_), .B(new_new_n270_), .Y(new_new_n417_));
  NO3        g395(.A(new_new_n417_), .B(new_new_n414_), .C(new_new_n412_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n190_), .B(new_new_n90_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n309_), .B(new_new_n80_), .Y(new_new_n420_));
  AOI210     g398(.A0(new_new_n420_), .A1(new_new_n419_), .B0(new_new_n307_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n188_), .B(i_10_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n63_), .B(i_2_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n280_), .B(new_new_n229_), .Y(new_new_n424_));
  OAI220     g402(.A0(new_new_n424_), .A1(new_new_n177_), .B0(new_new_n423_), .B1(new_new_n422_), .Y(new_new_n425_));
  NA3        g403(.A(new_new_n321_), .B(new_new_n320_), .C(i_5_), .Y(new_new_n426_));
  INV        g404(.A(new_new_n300_), .Y(new_new_n427_));
  OAI210     g405(.A0(new_new_n427_), .A1(new_new_n184_), .B0(new_new_n426_), .Y(new_new_n428_));
  NO3        g406(.A(new_new_n428_), .B(new_new_n425_), .C(new_new_n421_), .Y(new_new_n429_));
  AOI210     g407(.A0(new_new_n429_), .A1(new_new_n418_), .B0(new_new_n257_), .Y(new_new_n430_));
  NO4        g408(.A(new_new_n430_), .B(new_new_n411_), .C(new_new_n393_), .D(new_new_n368_), .Y(new_new_n431_));
  NO2        g409(.A(new_new_n70_), .B(i_13_), .Y(new_new_n432_));
  NO2        g410(.A(i_10_), .B(i_9_), .Y(new_new_n433_));
  NAi21      g411(.An(i_12_), .B(i_8_), .Y(new_new_n434_));
  NO2        g412(.A(new_new_n434_), .B(i_3_), .Y(new_new_n435_));
  NA2        g413(.A(i_2_), .B(new_new_n98_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n436_), .B(new_new_n199_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n293_), .B(i_0_), .Y(new_new_n438_));
  NO3        g416(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n252_), .B(new_new_n91_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n440_), .B(new_new_n439_), .Y(new_new_n441_));
  NA2        g419(.A(i_8_), .B(i_9_), .Y(new_new_n442_));
  NO3        g420(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n443_));
  NA3        g421(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n444_));
  NA4        g422(.A(new_new_n140_), .B(new_new_n110_), .C(new_new_n77_), .D(new_new_n23_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n445_), .B(new_new_n444_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n446_), .B(new_new_n437_), .Y(new_new_n447_));
  OA210      g425(.A0(new_new_n336_), .A1(new_new_n95_), .B0(new_new_n281_), .Y(new_new_n448_));
  OA220      g426(.A0(new_new_n448_), .A1(new_new_n156_), .B0(new_new_n202_), .B1(new_new_n226_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n90_), .B(i_13_), .Y(new_new_n450_));
  NA2        g428(.A(new_new_n415_), .B(new_new_n369_), .Y(new_new_n451_));
  NO2        g429(.A(i_2_), .B(i_13_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n451_), .B(new_new_n450_), .Y(new_new_n453_));
  NO3        g431(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n454_));
  NO2        g432(.A(i_6_), .B(i_7_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n455_), .B(new_new_n454_), .Y(new_new_n456_));
  NO2        g434(.A(i_11_), .B(i_1_), .Y(new_new_n457_));
  OR2        g435(.A(i_11_), .B(i_8_), .Y(new_new_n458_));
  NOi21      g436(.An(i_2_), .B(i_7_), .Y(new_new_n459_));
  NAi31      g437(.An(new_new_n458_), .B(new_new_n459_), .C(i_0_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n403_), .B(i_6_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n461_), .B(i_1_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n462_), .B(new_new_n460_), .Y(new_new_n463_));
  NO2        g441(.A(i_3_), .B(new_new_n188_), .Y(new_new_n464_));
  NO2        g442(.A(i_6_), .B(i_10_), .Y(new_new_n465_));
  NA3        g443(.A(new_new_n465_), .B(new_new_n297_), .C(new_new_n464_), .Y(new_new_n466_));
  NO2        g444(.A(new_new_n466_), .B(new_new_n149_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n151_), .B(i_3_), .Y(new_new_n469_));
  NO3        g447(.A(new_new_n467_), .B(new_new_n463_), .C(new_new_n453_), .Y(new_new_n470_));
  NAi21      g448(.An(new_new_n211_), .B(new_new_n384_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n321_), .B(new_new_n213_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n26_), .B(i_5_), .Y(new_new_n473_));
  NA3        g451(.A(i_6_), .B(new_new_n473_), .C(new_new_n137_), .Y(new_new_n474_));
  OR3        g452(.A(new_new_n287_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n475_));
  OAI220     g453(.A0(new_new_n475_), .A1(new_new_n474_), .B0(new_new_n472_), .B1(new_new_n471_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n27_), .B(i_10_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n297_), .B(new_new_n231_), .Y(new_new_n478_));
  OAI220     g456(.A0(new_new_n478_), .A1(new_new_n423_), .B0(new_new_n477_), .B1(new_new_n450_), .Y(new_new_n479_));
  NA3        g457(.A(new_new_n290_), .B(new_new_n217_), .C(new_new_n70_), .Y(new_new_n480_));
  NO2        g458(.A(new_new_n480_), .B(new_new_n456_), .Y(new_new_n481_));
  NO3        g459(.A(new_new_n481_), .B(new_new_n479_), .C(new_new_n476_), .Y(new_new_n482_));
  NA4        g460(.A(new_new_n482_), .B(new_new_n470_), .C(new_new_n449_), .D(new_new_n447_), .Y(new_new_n483_));
  NA3        g461(.A(new_new_n290_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n484_));
  INV        g462(.A(new_new_n484_), .Y(new_new_n485_));
  BUFFER     g463(.A(new_new_n271_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n486_), .B(new_new_n485_), .Y(new_new_n487_));
  AN2        g465(.A(i_11_), .B(new_new_n439_), .Y(new_new_n488_));
  INV        g466(.A(new_new_n158_), .Y(new_new_n489_));
  OAI210     g467(.A0(new_new_n489_), .A1(new_new_n226_), .B0(new_new_n291_), .Y(new_new_n490_));
  AOI220     g468(.A0(new_new_n490_), .A1(new_new_n308_), .B0(new_new_n488_), .B1(new_new_n293_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n341_), .B(new_new_n70_), .Y(new_new_n492_));
  INV        g470(.A(new_new_n351_), .Y(new_new_n493_));
  NO2        g471(.A(new_new_n36_), .B(i_8_), .Y(new_new_n494_));
  NAi41      g472(.An(new_new_n492_), .B(new_new_n465_), .C(new_new_n494_), .D(new_new_n46_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n39_), .B(i_13_), .Y(new_new_n496_));
  INV        g474(.A(new_new_n495_), .Y(new_new_n497_));
  NO2        g475(.A(i_7_), .B(new_new_n193_), .Y(new_new_n498_));
  OR2        g476(.A(new_new_n177_), .B(i_4_), .Y(new_new_n499_));
  INV        g477(.A(new_new_n499_), .Y(new_new_n500_));
  AOI220     g478(.A0(new_new_n500_), .A1(new_new_n498_), .B0(i_1_), .B1(new_new_n404_), .Y(new_new_n501_));
  NA4        g479(.A(new_new_n501_), .B(new_new_n496_), .C(new_new_n491_), .D(new_new_n487_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n375_), .B(new_new_n279_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n371_), .B(new_new_n503_), .Y(new_new_n504_));
  NO2        g482(.A(i_12_), .B(new_new_n188_), .Y(new_new_n505_));
  NA2        g483(.A(new_new_n505_), .B(new_new_n219_), .Y(new_new_n506_));
  NO2        g484(.A(i_10_), .B(new_new_n506_), .Y(new_new_n507_));
  NOi31      g485(.An(new_new_n300_), .B(new_new_n403_), .C(new_new_n38_), .Y(new_new_n508_));
  OAI210     g486(.A0(new_new_n508_), .A1(new_new_n507_), .B0(new_new_n504_), .Y(new_new_n509_));
  NO2        g487(.A(i_8_), .B(i_7_), .Y(new_new_n510_));
  OAI210     g488(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n511_), .B(new_new_n217_), .Y(new_new_n512_));
  OAI220     g490(.A0(new_new_n46_), .A1(new_new_n499_), .B0(new_new_n512_), .B1(new_new_n234_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n44_), .B(i_10_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n514_), .B(i_6_), .Y(new_new_n515_));
  NA3        g493(.A(new_new_n515_), .B(new_new_n513_), .C(new_new_n510_), .Y(new_new_n516_));
  AOI220     g494(.A0(new_new_n415_), .A1(new_new_n309_), .B0(new_new_n239_), .B1(new_new_n236_), .Y(new_new_n517_));
  OAI220     g495(.A0(new_new_n517_), .A1(new_new_n248_), .B0(new_new_n450_), .B1(new_new_n128_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n518_), .B(new_new_n251_), .Y(new_new_n519_));
  NA3        g497(.A(new_new_n290_), .B(new_new_n168_), .C(new_new_n90_), .Y(new_new_n520_));
  NO2        g498(.A(new_new_n151_), .B(i_5_), .Y(new_new_n521_));
  NA2        g499(.A(new_new_n521_), .B(new_new_n303_), .Y(new_new_n522_));
  NA2        g500(.A(new_new_n522_), .B(new_new_n520_), .Y(new_new_n523_));
  NA2        g501(.A(new_new_n523_), .B(new_new_n443_), .Y(new_new_n524_));
  NA4        g502(.A(new_new_n524_), .B(new_new_n519_), .C(new_new_n516_), .D(new_new_n509_), .Y(new_new_n525_));
  NA2        g503(.A(new_new_n268_), .B(new_new_n79_), .Y(new_new_n526_));
  NO2        g504(.A(new_new_n333_), .B(new_new_n526_), .Y(new_new_n527_));
  NA2        g505(.A(new_new_n280_), .B(new_new_n271_), .Y(new_new_n528_));
  NO2        g506(.A(new_new_n528_), .B(new_new_n167_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n217_), .B(i_0_), .Y(new_new_n530_));
  NA2        g508(.A(new_new_n433_), .B(new_new_n216_), .Y(new_new_n531_));
  NO2        g509(.A(new_new_n530_), .B(new_new_n531_), .Y(new_new_n532_));
  AOI210     g510(.A0(new_new_n352_), .A1(new_new_n46_), .B0(new_new_n356_), .Y(new_new_n533_));
  NA2        g511(.A(i_0_), .B(new_new_n48_), .Y(new_new_n534_));
  NA3        g512(.A(new_new_n505_), .B(new_new_n259_), .C(new_new_n534_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n533_), .B(new_new_n535_), .Y(new_new_n536_));
  NO4        g514(.A(new_new_n536_), .B(new_new_n532_), .C(new_new_n529_), .D(new_new_n527_), .Y(new_new_n537_));
  NO4        g515(.A(new_new_n242_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n538_));
  NO3        g516(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n227_), .B(new_new_n36_), .Y(new_new_n540_));
  AN2        g518(.A(new_new_n540_), .B(new_new_n539_), .Y(new_new_n541_));
  OA210      g519(.A0(new_new_n541_), .A1(new_new_n538_), .B0(new_new_n341_), .Y(new_new_n542_));
  NO2        g520(.A(new_new_n403_), .B(i_1_), .Y(new_new_n543_));
  NOi31      g521(.An(new_new_n543_), .B(new_new_n440_), .C(new_new_n70_), .Y(new_new_n544_));
  AN3        g522(.A(new_new_n544_), .B(new_new_n401_), .C(new_new_n473_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n413_), .B(new_new_n171_), .Y(new_new_n546_));
  NO3        g524(.A(new_new_n546_), .B(new_new_n545_), .C(new_new_n542_), .Y(new_new_n547_));
  NOi21      g525(.An(i_10_), .B(i_6_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n80_), .B(new_new_n25_), .Y(new_new_n549_));
  AOI220     g527(.A0(new_new_n268_), .A1(new_new_n549_), .B0(new_new_n259_), .B1(new_new_n548_), .Y(new_new_n550_));
  NO2        g528(.A(new_new_n550_), .B(new_new_n438_), .Y(new_new_n551_));
  NO2        g529(.A(new_new_n109_), .B(new_new_n23_), .Y(new_new_n552_));
  NA2        g530(.A(new_new_n300_), .B(new_new_n158_), .Y(new_new_n553_));
  AOI220     g531(.A0(new_new_n553_), .A1(new_new_n424_), .B0(new_new_n178_), .B1(new_new_n176_), .Y(new_new_n554_));
  NOi21      g532(.An(new_new_n141_), .B(new_new_n316_), .Y(new_new_n555_));
  NO3        g533(.A(new_new_n555_), .B(new_new_n554_), .C(new_new_n551_), .Y(new_new_n556_));
  NO2        g534(.A(new_new_n492_), .B(new_new_n365_), .Y(new_new_n557_));
  INV        g535(.A(new_new_n303_), .Y(new_new_n558_));
  NO2        g536(.A(i_12_), .B(new_new_n80_), .Y(new_new_n559_));
  NA3        g537(.A(new_new_n559_), .B(new_new_n259_), .C(new_new_n534_), .Y(new_new_n560_));
  NA2        g538(.A(new_new_n372_), .B(new_new_n268_), .Y(new_new_n561_));
  AOI210     g539(.A0(new_new_n561_), .A1(new_new_n560_), .B0(new_new_n558_), .Y(new_new_n562_));
  NO3        g540(.A(i_4_), .B(new_new_n327_), .C(new_new_n285_), .Y(new_new_n563_));
  OR2        g541(.A(i_2_), .B(i_5_), .Y(new_new_n564_));
  OR2        g542(.A(new_new_n564_), .B(new_new_n396_), .Y(new_new_n565_));
  NA2        g543(.A(new_new_n360_), .B(new_new_n236_), .Y(new_new_n566_));
  AOI210     g544(.A0(new_new_n566_), .A1(new_new_n565_), .B0(new_new_n471_), .Y(new_new_n567_));
  NO4        g545(.A(new_new_n567_), .B(new_new_n563_), .C(new_new_n562_), .D(new_new_n557_), .Y(new_new_n568_));
  NA4        g546(.A(new_new_n568_), .B(new_new_n556_), .C(new_new_n547_), .D(new_new_n537_), .Y(new_new_n569_));
  NO4        g547(.A(new_new_n569_), .B(new_new_n525_), .C(new_new_n502_), .D(new_new_n483_), .Y(new_new_n570_));
  NA4        g548(.A(new_new_n570_), .B(new_new_n431_), .C(new_new_n340_), .D(new_new_n296_), .Y(mai7));
  NO2        g549(.A(new_new_n87_), .B(new_new_n53_), .Y(new_new_n572_));
  NO2        g550(.A(new_new_n102_), .B(new_new_n84_), .Y(new_new_n573_));
  NA2        g551(.A(i_3_), .B(new_new_n573_), .Y(new_new_n574_));
  NA2        g552(.A(new_new_n465_), .B(new_new_n79_), .Y(new_new_n575_));
  NA2        g553(.A(i_11_), .B(new_new_n188_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n139_), .B(new_new_n576_), .Y(new_new_n577_));
  OAI210     g555(.A0(new_new_n577_), .A1(new_new_n575_), .B0(new_new_n574_), .Y(new_new_n578_));
  NO2        g556(.A(new_new_n230_), .B(i_4_), .Y(new_new_n579_));
  NA2        g557(.A(new_new_n579_), .B(i_8_), .Y(new_new_n580_));
  NA2        g558(.A(i_2_), .B(new_new_n80_), .Y(new_new_n581_));
  OAI210     g559(.A0(new_new_n83_), .A1(new_new_n197_), .B0(new_new_n198_), .Y(new_new_n582_));
  NO2        g560(.A(i_7_), .B(new_new_n37_), .Y(new_new_n583_));
  NA2        g561(.A(i_4_), .B(i_8_), .Y(new_new_n584_));
  NO2        g562(.A(new_new_n578_), .B(new_new_n572_), .Y(new_new_n585_));
  INV        g563(.A(new_new_n155_), .Y(new_new_n586_));
  OR2        g564(.A(i_6_), .B(i_10_), .Y(new_new_n587_));
  NO2        g565(.A(new_new_n587_), .B(new_new_n23_), .Y(new_new_n588_));
  OR3        g566(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n589_));
  NO3        g567(.A(new_new_n589_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n590_));
  INV        g568(.A(new_new_n194_), .Y(new_new_n591_));
  NO2        g569(.A(new_new_n590_), .B(new_new_n588_), .Y(new_new_n592_));
  OA220      g570(.A0(new_new_n592_), .A1(new_new_n558_), .B0(new_new_n586_), .B1(new_new_n253_), .Y(new_new_n593_));
  AOI210     g571(.A0(new_new_n593_), .A1(new_new_n585_), .B0(new_new_n62_), .Y(new_new_n594_));
  NOi21      g572(.An(i_11_), .B(i_7_), .Y(new_new_n595_));
  AO210      g573(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n596_));
  NO2        g574(.A(new_new_n596_), .B(new_new_n595_), .Y(new_new_n597_));
  NA2        g575(.A(new_new_n597_), .B(new_new_n201_), .Y(new_new_n598_));
  NA3        g576(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n599_));
  NAi31      g577(.An(new_new_n599_), .B(new_new_n210_), .C(i_11_), .Y(new_new_n600_));
  AOI210     g578(.A0(new_new_n600_), .A1(new_new_n598_), .B0(new_new_n62_), .Y(new_new_n601_));
  NA2        g579(.A(new_new_n82_), .B(new_new_n62_), .Y(new_new_n602_));
  AO210      g580(.A0(new_new_n602_), .A1(new_new_n365_), .B0(new_new_n41_), .Y(new_new_n603_));
  NO3        g581(.A(i_7_), .B(new_new_n203_), .C(new_new_n576_), .Y(new_new_n604_));
  OAI210     g582(.A0(new_new_n604_), .A1(new_new_n220_), .B0(new_new_n62_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n397_), .B(new_new_n31_), .Y(new_new_n606_));
  OR2        g584(.A(new_new_n203_), .B(new_new_n102_), .Y(new_new_n607_));
  NA2        g585(.A(new_new_n607_), .B(new_new_n606_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n62_), .B(i_9_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n609_), .B(i_4_), .Y(new_new_n610_));
  NA2        g588(.A(new_new_n610_), .B(new_new_n608_), .Y(new_new_n611_));
  NO2        g589(.A(i_1_), .B(i_12_), .Y(new_new_n612_));
  NA3        g590(.A(new_new_n612_), .B(new_new_n104_), .C(new_new_n24_), .Y(new_new_n613_));
  NA4        g591(.A(new_new_n613_), .B(new_new_n611_), .C(new_new_n605_), .D(new_new_n603_), .Y(new_new_n614_));
  OAI210     g592(.A0(new_new_n614_), .A1(new_new_n601_), .B0(i_6_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n599_), .B(new_new_n102_), .Y(new_new_n616_));
  NA2        g594(.A(new_new_n616_), .B(new_new_n559_), .Y(new_new_n617_));
  NO2        g595(.A(i_6_), .B(i_11_), .Y(new_new_n618_));
  NA2        g596(.A(new_new_n617_), .B(new_new_n441_), .Y(new_new_n619_));
  NO4        g597(.A(new_new_n210_), .B(new_new_n123_), .C(i_13_), .D(new_new_n80_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n620_), .B(new_new_n609_), .Y(new_new_n621_));
  INV        g599(.A(new_new_n621_), .Y(new_new_n622_));
  NA3        g600(.A(new_new_n510_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n623_));
  NA2        g601(.A(new_new_n133_), .B(i_9_), .Y(new_new_n624_));
  NA3        g602(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n46_), .B(i_1_), .Y(new_new_n626_));
  NA3        g604(.A(new_new_n626_), .B(new_new_n252_), .C(new_new_n44_), .Y(new_new_n627_));
  OAI220     g605(.A0(new_new_n627_), .A1(new_new_n625_), .B0(new_new_n624_), .B1(new_new_n1003_), .Y(new_new_n628_));
  NA3        g606(.A(new_new_n609_), .B(new_new_n303_), .C(i_6_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n629_), .B(new_new_n23_), .Y(new_new_n630_));
  AOI210     g608(.A0(new_new_n457_), .A1(new_new_n406_), .B0(new_new_n233_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n631_), .B(new_new_n581_), .Y(new_new_n632_));
  NAi21      g610(.An(new_new_n623_), .B(new_new_n86_), .Y(new_new_n633_));
  NA2        g611(.A(new_new_n626_), .B(new_new_n252_), .Y(new_new_n634_));
  NO2        g612(.A(i_11_), .B(new_new_n37_), .Y(new_new_n635_));
  NA2        g613(.A(new_new_n635_), .B(new_new_n24_), .Y(new_new_n636_));
  OAI210     g614(.A0(new_new_n636_), .A1(new_new_n634_), .B0(new_new_n633_), .Y(new_new_n637_));
  OR4        g615(.A(new_new_n637_), .B(new_new_n632_), .C(new_new_n630_), .D(new_new_n628_), .Y(new_new_n638_));
  NO3        g616(.A(new_new_n638_), .B(new_new_n622_), .C(new_new_n619_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n230_), .B(new_new_n95_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n640_), .B(new_new_n595_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n641_), .B(i_1_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n642_), .B(new_new_n589_), .Y(new_new_n643_));
  NA2        g621(.A(new_new_n643_), .B(new_new_n46_), .Y(new_new_n644_));
  NA2        g622(.A(i_3_), .B(new_new_n188_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n645_), .B(new_new_n109_), .Y(new_new_n646_));
  AN2        g624(.A(new_new_n646_), .B(new_new_n515_), .Y(new_new_n647_));
  NO2        g625(.A(new_new_n112_), .B(new_new_n37_), .Y(new_new_n648_));
  NO2        g626(.A(new_new_n80_), .B(i_9_), .Y(new_new_n649_));
  NA2        g627(.A(i_1_), .B(i_3_), .Y(new_new_n650_));
  NO2        g628(.A(new_new_n442_), .B(new_new_n87_), .Y(new_new_n651_));
  INV        g629(.A(new_new_n651_), .Y(new_new_n652_));
  NO2        g630(.A(new_new_n652_), .B(new_new_n650_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n653_), .B(new_new_n647_), .Y(new_new_n654_));
  NA4        g632(.A(new_new_n654_), .B(new_new_n644_), .C(new_new_n639_), .D(new_new_n615_), .Y(new_new_n655_));
  NO3        g633(.A(new_new_n458_), .B(i_3_), .C(i_7_), .Y(new_new_n656_));
  NOi21      g634(.An(new_new_n656_), .B(i_10_), .Y(new_new_n657_));
  OA210      g635(.A0(new_new_n657_), .A1(new_new_n237_), .B0(new_new_n80_), .Y(new_new_n658_));
  NA2        g636(.A(new_new_n359_), .B(new_new_n358_), .Y(new_new_n659_));
  NA3        g637(.A(new_new_n465_), .B(new_new_n494_), .C(new_new_n46_), .Y(new_new_n660_));
  NO3        g638(.A(new_new_n459_), .B(new_new_n584_), .C(new_new_n80_), .Y(new_new_n661_));
  NA2        g639(.A(new_new_n661_), .B(new_new_n25_), .Y(new_new_n662_));
  NA3        g640(.A(new_new_n155_), .B(new_new_n79_), .C(new_new_n80_), .Y(new_new_n663_));
  NA4        g641(.A(new_new_n663_), .B(new_new_n662_), .C(new_new_n660_), .D(new_new_n659_), .Y(new_new_n664_));
  OAI210     g642(.A0(new_new_n664_), .A1(new_new_n658_), .B0(i_1_), .Y(new_new_n665_));
  AOI210     g643(.A0(new_new_n252_), .A1(new_new_n91_), .B0(i_1_), .Y(new_new_n666_));
  NO2        g644(.A(new_new_n357_), .B(i_2_), .Y(new_new_n667_));
  NA2        g645(.A(new_new_n667_), .B(new_new_n666_), .Y(new_new_n668_));
  OAI210     g646(.A0(new_new_n629_), .A1(new_new_n434_), .B0(new_new_n668_), .Y(new_new_n669_));
  INV        g647(.A(new_new_n669_), .Y(new_new_n670_));
  AOI210     g648(.A0(new_new_n670_), .A1(new_new_n665_), .B0(i_13_), .Y(new_new_n671_));
  OR2        g649(.A(i_11_), .B(i_7_), .Y(new_new_n672_));
  NA3        g650(.A(new_new_n672_), .B(new_new_n100_), .C(new_new_n133_), .Y(new_new_n673_));
  AOI220     g651(.A0(new_new_n452_), .A1(new_new_n155_), .B0(i_2_), .B1(new_new_n133_), .Y(new_new_n674_));
  OAI210     g652(.A0(new_new_n674_), .A1(new_new_n44_), .B0(new_new_n673_), .Y(new_new_n675_));
  AOI210     g653(.A0(new_new_n625_), .A1(new_new_n53_), .B0(i_12_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n237_), .B(new_new_n126_), .Y(new_new_n677_));
  OAI220     g655(.A0(new_new_n677_), .A1(new_new_n41_), .B0(new_new_n1002_), .B1(new_new_n87_), .Y(new_new_n678_));
  AOI210     g656(.A0(new_new_n675_), .A1(new_new_n318_), .B0(new_new_n678_), .Y(new_new_n679_));
  AOI220     g657(.A0(i_12_), .A1(new_new_n69_), .B0(new_new_n372_), .B1(new_new_n626_), .Y(new_new_n680_));
  NO2        g658(.A(new_new_n680_), .B(new_new_n234_), .Y(new_new_n681_));
  AOI210     g659(.A0(new_new_n434_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n682_));
  NOi31      g660(.An(new_new_n682_), .B(new_new_n575_), .C(new_new_n44_), .Y(new_new_n683_));
  NA2        g661(.A(new_new_n122_), .B(i_13_), .Y(new_new_n684_));
  NO2        g662(.A(new_new_n625_), .B(new_new_n109_), .Y(new_new_n685_));
  INV        g663(.A(new_new_n685_), .Y(new_new_n686_));
  OAI220     g664(.A0(new_new_n686_), .A1(new_new_n68_), .B0(new_new_n684_), .B1(new_new_n666_), .Y(new_new_n687_));
  NO3        g665(.A(new_new_n68_), .B(new_new_n32_), .C(new_new_n95_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n26_), .B(new_new_n188_), .Y(new_new_n689_));
  NA2        g667(.A(new_new_n689_), .B(i_7_), .Y(new_new_n690_));
  NO3        g668(.A(new_new_n459_), .B(new_new_n230_), .C(new_new_n80_), .Y(new_new_n691_));
  AOI210     g669(.A0(new_new_n691_), .A1(new_new_n690_), .B0(new_new_n688_), .Y(new_new_n692_));
  NA2        g670(.A(new_new_n86_), .B(new_new_n96_), .Y(new_new_n693_));
  OAI220     g671(.A0(new_new_n693_), .A1(new_new_n580_), .B0(new_new_n692_), .B1(new_new_n591_), .Y(new_new_n694_));
  NO4        g672(.A(new_new_n694_), .B(new_new_n687_), .C(new_new_n683_), .D(new_new_n681_), .Y(new_new_n695_));
  OR2        g673(.A(i_11_), .B(i_6_), .Y(new_new_n696_));
  NA3        g674(.A(new_new_n579_), .B(new_new_n689_), .C(i_7_), .Y(new_new_n697_));
  AOI210     g675(.A0(new_new_n697_), .A1(new_new_n686_), .B0(new_new_n696_), .Y(new_new_n698_));
  NA3        g676(.A(new_new_n397_), .B(new_new_n583_), .C(new_new_n91_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n618_), .B(i_13_), .Y(new_new_n700_));
  NAi21      g678(.An(i_11_), .B(i_12_), .Y(new_new_n701_));
  NOi41      g679(.An(new_new_n105_), .B(new_new_n701_), .C(i_13_), .D(new_new_n80_), .Y(new_new_n702_));
  NO3        g680(.A(new_new_n459_), .B(new_new_n559_), .C(new_new_n584_), .Y(new_new_n703_));
  AOI210     g681(.A0(new_new_n703_), .A1(new_new_n297_), .B0(new_new_n702_), .Y(new_new_n704_));
  NA3        g682(.A(new_new_n704_), .B(new_new_n700_), .C(new_new_n699_), .Y(new_new_n705_));
  OAI210     g683(.A0(new_new_n705_), .A1(new_new_n698_), .B0(new_new_n62_), .Y(new_new_n706_));
  OAI210     g684(.A0(new_new_n230_), .A1(new_new_n358_), .B0(new_new_n356_), .Y(new_new_n707_));
  NO2        g685(.A(new_new_n123_), .B(i_2_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n708_), .B(new_new_n612_), .Y(new_new_n709_));
  NA2        g687(.A(new_new_n709_), .B(new_new_n707_), .Y(new_new_n710_));
  NA3        g688(.A(new_new_n710_), .B(new_new_n45_), .C(new_new_n219_), .Y(new_new_n711_));
  NA4        g689(.A(new_new_n711_), .B(new_new_n706_), .C(new_new_n695_), .D(new_new_n679_), .Y(new_new_n712_));
  OR4        g690(.A(new_new_n712_), .B(new_new_n671_), .C(new_new_n655_), .D(new_new_n594_), .Y(mai5));
  AOI210     g691(.A0(new_new_n641_), .A1(new_new_n255_), .B0(new_new_n404_), .Y(new_new_n714_));
  NO2        g692(.A(new_new_n580_), .B(i_11_), .Y(new_new_n715_));
  NA2        g693(.A(new_new_n83_), .B(new_new_n715_), .Y(new_new_n716_));
  NA2        g694(.A(new_new_n716_), .B(new_new_n714_), .Y(new_new_n717_));
  NO3        g695(.A(i_11_), .B(new_new_n230_), .C(i_13_), .Y(new_new_n718_));
  NO2        g696(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n719_));
  NA2        g697(.A(i_12_), .B(i_8_), .Y(new_new_n720_));
  OAI210     g698(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n720_), .Y(new_new_n721_));
  INV        g699(.A(new_new_n433_), .Y(new_new_n722_));
  AOI220     g700(.A0(new_new_n303_), .A1(new_new_n552_), .B0(new_new_n721_), .B1(new_new_n719_), .Y(new_new_n723_));
  INV        g701(.A(new_new_n723_), .Y(new_new_n724_));
  NO2        g702(.A(new_new_n724_), .B(new_new_n717_), .Y(new_new_n725_));
  INV        g703(.A(new_new_n165_), .Y(new_new_n726_));
  INV        g704(.A(new_new_n237_), .Y(new_new_n727_));
  OAI210     g705(.A0(new_new_n667_), .A1(new_new_n435_), .B0(new_new_n105_), .Y(new_new_n728_));
  AOI210     g706(.A0(new_new_n728_), .A1(new_new_n727_), .B0(new_new_n726_), .Y(new_new_n729_));
  NO2        g707(.A(new_new_n442_), .B(new_new_n26_), .Y(new_new_n730_));
  NO2        g708(.A(new_new_n730_), .B(new_new_n406_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n731_), .B(i_2_), .Y(new_new_n732_));
  INV        g710(.A(new_new_n732_), .Y(new_new_n733_));
  AOI210     g711(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n403_), .Y(new_new_n734_));
  AOI210     g712(.A0(new_new_n734_), .A1(new_new_n733_), .B0(new_new_n729_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n185_), .B(new_new_n120_), .Y(new_new_n736_));
  OAI210     g714(.A0(new_new_n736_), .A1(new_new_n719_), .B0(i_2_), .Y(new_new_n737_));
  NO2        g715(.A(new_new_n737_), .B(new_new_n188_), .Y(new_new_n738_));
  OA210      g716(.A0(new_new_n597_), .A1(new_new_n121_), .B0(i_13_), .Y(new_new_n739_));
  NA2        g717(.A(new_new_n194_), .B(new_new_n197_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n146_), .B(new_new_n576_), .Y(new_new_n741_));
  AOI210     g719(.A0(new_new_n741_), .A1(new_new_n740_), .B0(new_new_n360_), .Y(new_new_n742_));
  AOI210     g720(.A0(new_new_n203_), .A1(new_new_n143_), .B0(new_new_n494_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n743_), .B(new_new_n406_), .Y(new_new_n744_));
  NO2        g722(.A(new_new_n96_), .B(new_new_n44_), .Y(new_new_n745_));
  INV        g723(.A(new_new_n286_), .Y(new_new_n746_));
  NA4        g724(.A(new_new_n746_), .B(new_new_n290_), .C(new_new_n119_), .D(new_new_n42_), .Y(new_new_n747_));
  OAI210     g725(.A0(new_new_n747_), .A1(new_new_n745_), .B0(new_new_n744_), .Y(new_new_n748_));
  NO4        g726(.A(new_new_n748_), .B(new_new_n742_), .C(new_new_n739_), .D(new_new_n738_), .Y(new_new_n749_));
  NA2        g727(.A(new_new_n552_), .B(new_new_n28_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n718_), .B(new_new_n260_), .Y(new_new_n751_));
  NA2        g729(.A(new_new_n751_), .B(new_new_n750_), .Y(new_new_n752_));
  NO2        g730(.A(new_new_n61_), .B(i_12_), .Y(new_new_n753_));
  NO2        g731(.A(new_new_n753_), .B(new_new_n121_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n754_), .B(new_new_n576_), .Y(new_new_n755_));
  AOI220     g733(.A0(new_new_n755_), .A1(new_new_n36_), .B0(new_new_n752_), .B1(new_new_n46_), .Y(new_new_n756_));
  NA4        g734(.A(new_new_n756_), .B(new_new_n749_), .C(new_new_n735_), .D(new_new_n725_), .Y(mai6));
  NO3        g735(.A(new_new_n244_), .B(new_new_n292_), .C(i_1_), .Y(new_new_n758_));
  NO2        g736(.A(new_new_n180_), .B(new_new_n134_), .Y(new_new_n759_));
  OAI210     g737(.A0(new_new_n759_), .A1(new_new_n758_), .B0(new_new_n708_), .Y(new_new_n760_));
  NA4        g738(.A(new_new_n376_), .B(new_new_n464_), .C(new_new_n68_), .D(new_new_n95_), .Y(new_new_n761_));
  INV        g739(.A(new_new_n761_), .Y(new_new_n762_));
  NO2        g740(.A(new_new_n215_), .B(new_new_n468_), .Y(new_new_n763_));
  NO2        g741(.A(i_11_), .B(i_9_), .Y(new_new_n764_));
  NO2        g742(.A(new_new_n762_), .B(new_new_n314_), .Y(new_new_n765_));
  AO210      g743(.A0(new_new_n765_), .A1(new_new_n760_), .B0(i_12_), .Y(new_new_n766_));
  NA2        g744(.A(new_new_n361_), .B(new_new_n321_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n559_), .B(new_new_n62_), .Y(new_new_n768_));
  NA2        g746(.A(new_new_n657_), .B(new_new_n68_), .Y(new_new_n769_));
  NA4        g747(.A(new_new_n602_), .B(new_new_n769_), .C(new_new_n768_), .D(new_new_n767_), .Y(new_new_n770_));
  INV        g748(.A(new_new_n191_), .Y(new_new_n771_));
  AOI220     g749(.A0(new_new_n771_), .A1(new_new_n764_), .B0(new_new_n770_), .B1(new_new_n70_), .Y(new_new_n772_));
  INV        g750(.A(new_new_n313_), .Y(new_new_n773_));
  NA2        g751(.A(new_new_n72_), .B(new_new_n126_), .Y(new_new_n774_));
  NO2        g752(.A(new_new_n774_), .B(new_new_n773_), .Y(new_new_n775_));
  NO2        g753(.A(new_new_n32_), .B(i_11_), .Y(new_new_n776_));
  NA3        g754(.A(new_new_n776_), .B(new_new_n455_), .C(new_new_n376_), .Y(new_new_n777_));
  NAi32      g755(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n778_));
  AOI210     g756(.A0(new_new_n696_), .A1(new_new_n81_), .B0(new_new_n778_), .Y(new_new_n779_));
  OAI210     g757(.A0(new_new_n656_), .A1(new_new_n540_), .B0(new_new_n539_), .Y(new_new_n780_));
  NAi31      g758(.An(new_new_n779_), .B(new_new_n780_), .C(new_new_n777_), .Y(new_new_n781_));
  OR2        g759(.A(new_new_n781_), .B(new_new_n775_), .Y(new_new_n782_));
  NO2        g760(.A(new_new_n672_), .B(i_2_), .Y(new_new_n783_));
  NA2        g761(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n784_));
  OAI210     g762(.A0(new_new_n784_), .A1(new_new_n396_), .B0(new_new_n346_), .Y(new_new_n785_));
  NA2        g763(.A(new_new_n785_), .B(new_new_n783_), .Y(new_new_n786_));
  AO220      g764(.A0(new_new_n345_), .A1(new_new_n335_), .B0(new_new_n382_), .B1(new_new_n576_), .Y(new_new_n787_));
  NA3        g765(.A(new_new_n787_), .B(new_new_n245_), .C(i_7_), .Y(new_new_n788_));
  OR2        g766(.A(new_new_n597_), .B(new_new_n435_), .Y(new_new_n789_));
  NA3        g767(.A(new_new_n789_), .B(new_new_n142_), .C(new_new_n66_), .Y(new_new_n790_));
  OR2        g768(.A(new_new_n722_), .B(new_new_n36_), .Y(new_new_n791_));
  NA4        g769(.A(new_new_n791_), .B(new_new_n790_), .C(new_new_n788_), .D(new_new_n786_), .Y(new_new_n792_));
  OAI210     g770(.A0(i_6_), .A1(i_11_), .B0(new_new_n81_), .Y(new_new_n793_));
  AOI220     g771(.A0(new_new_n793_), .A1(new_new_n539_), .B0(new_new_n763_), .B1(new_new_n690_), .Y(new_new_n794_));
  NA3        g772(.A(new_new_n360_), .B(new_new_n231_), .C(new_new_n142_), .Y(new_new_n795_));
  NA2        g773(.A(new_new_n382_), .B(new_new_n67_), .Y(new_new_n796_));
  NA4        g774(.A(new_new_n796_), .B(new_new_n795_), .C(new_new_n794_), .D(new_new_n582_), .Y(new_new_n797_));
  AO210      g775(.A0(new_new_n494_), .A1(new_new_n46_), .B0(new_new_n82_), .Y(new_new_n798_));
  NA3        g776(.A(new_new_n798_), .B(new_new_n465_), .C(new_new_n213_), .Y(new_new_n799_));
  AOI210     g777(.A0(new_new_n435_), .A1(new_new_n433_), .B0(new_new_n538_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n587_), .B(new_new_n96_), .Y(new_new_n801_));
  OAI210     g779(.A0(new_new_n801_), .A1(new_new_n106_), .B0(new_new_n395_), .Y(new_new_n802_));
  INV        g780(.A(new_new_n565_), .Y(new_new_n803_));
  NA3        g781(.A(new_new_n803_), .B(new_new_n313_), .C(i_7_), .Y(new_new_n804_));
  NA4        g782(.A(new_new_n804_), .B(new_new_n802_), .C(new_new_n800_), .D(new_new_n799_), .Y(new_new_n805_));
  NO4        g783(.A(new_new_n805_), .B(new_new_n797_), .C(new_new_n792_), .D(new_new_n782_), .Y(new_new_n806_));
  NA4        g784(.A(new_new_n806_), .B(new_new_n772_), .C(new_new_n766_), .D(new_new_n367_), .Y(mai3));
  NA2        g785(.A(i_6_), .B(i_7_), .Y(new_new_n808_));
  NO2        g786(.A(new_new_n808_), .B(i_0_), .Y(new_new_n809_));
  NO2        g787(.A(i_11_), .B(new_new_n230_), .Y(new_new_n810_));
  OAI210     g788(.A0(new_new_n809_), .A1(new_new_n274_), .B0(new_new_n810_), .Y(new_new_n811_));
  INV        g789(.A(new_new_n811_), .Y(new_new_n812_));
  NO3        g790(.A(new_new_n438_), .B(new_new_n84_), .C(new_new_n44_), .Y(new_new_n813_));
  OA210      g791(.A0(new_new_n813_), .A1(new_new_n812_), .B0(new_new_n168_), .Y(new_new_n814_));
  INV        g792(.A(new_new_n795_), .Y(new_new_n815_));
  NA2        g793(.A(new_new_n815_), .B(new_new_n40_), .Y(new_new_n816_));
  NO3        g794(.A(new_new_n607_), .B(new_new_n442_), .C(new_new_n126_), .Y(new_new_n817_));
  NA2        g795(.A(new_new_n397_), .B(new_new_n45_), .Y(new_new_n818_));
  AN2        g796(.A(new_new_n440_), .B(new_new_n54_), .Y(new_new_n819_));
  NO2        g797(.A(new_new_n819_), .B(new_new_n817_), .Y(new_new_n820_));
  AOI210     g798(.A0(new_new_n820_), .A1(new_new_n816_), .B0(new_new_n48_), .Y(new_new_n821_));
  NO4        g799(.A(new_new_n364_), .B(new_new_n370_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n822_));
  NA2        g800(.A(new_new_n180_), .B(new_new_n548_), .Y(new_new_n823_));
  NOi21      g801(.An(new_new_n823_), .B(new_new_n822_), .Y(new_new_n824_));
  NA2        g802(.A(new_new_n682_), .B(new_new_n649_), .Y(new_new_n825_));
  NA2        g803(.A(new_new_n319_), .B(i_5_), .Y(new_new_n826_));
  OAI220     g804(.A0(new_new_n826_), .A1(new_new_n825_), .B0(new_new_n824_), .B1(new_new_n62_), .Y(new_new_n827_));
  NOi21      g805(.An(i_5_), .B(i_9_), .Y(new_new_n828_));
  NA2        g806(.A(new_new_n828_), .B(new_new_n432_), .Y(new_new_n829_));
  AOI210     g807(.A0(new_new_n252_), .A1(new_new_n457_), .B0(new_new_n661_), .Y(new_new_n830_));
  NO3        g808(.A(new_new_n400_), .B(new_new_n252_), .C(new_new_n70_), .Y(new_new_n831_));
  NO2        g809(.A(new_new_n169_), .B(new_new_n143_), .Y(new_new_n832_));
  AOI210     g810(.A0(new_new_n832_), .A1(new_new_n236_), .B0(new_new_n831_), .Y(new_new_n833_));
  OAI220     g811(.A0(new_new_n833_), .A1(new_new_n175_), .B0(new_new_n830_), .B1(new_new_n829_), .Y(new_new_n834_));
  NO4        g812(.A(new_new_n834_), .B(new_new_n827_), .C(new_new_n821_), .D(new_new_n814_), .Y(new_new_n835_));
  NA2        g813(.A(new_new_n180_), .B(new_new_n24_), .Y(new_new_n836_));
  NO2        g814(.A(new_new_n648_), .B(new_new_n573_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n837_), .B(new_new_n836_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n297_), .B(new_new_n124_), .Y(new_new_n839_));
  NAi21      g817(.An(new_new_n156_), .B(i_5_), .Y(new_new_n840_));
  NO2        g818(.A(new_new_n839_), .B(new_new_n387_), .Y(new_new_n841_));
  NO2        g819(.A(new_new_n841_), .B(new_new_n838_), .Y(new_new_n842_));
  NA2        g820(.A(new_new_n549_), .B(i_0_), .Y(new_new_n843_));
  NO3        g821(.A(new_new_n843_), .B(new_new_n371_), .C(new_new_n83_), .Y(new_new_n844_));
  NO4        g822(.A(new_new_n564_), .B(new_new_n210_), .C(new_new_n403_), .D(new_new_n396_), .Y(new_new_n845_));
  AOI210     g823(.A0(new_new_n845_), .A1(i_11_), .B0(new_new_n844_), .Y(new_new_n846_));
  AN2        g824(.A(new_new_n90_), .B(new_new_n235_), .Y(new_new_n847_));
  NA2        g825(.A(new_new_n718_), .B(new_new_n314_), .Y(new_new_n848_));
  AOI210     g826(.A0(new_new_n465_), .A1(new_new_n83_), .B0(new_new_n57_), .Y(new_new_n849_));
  OAI220     g827(.A0(new_new_n849_), .A1(new_new_n848_), .B0(new_new_n636_), .B1(new_new_n512_), .Y(new_new_n850_));
  INV        g828(.A(new_new_n514_), .Y(new_new_n851_));
  NO4        g829(.A(new_new_n109_), .B(new_new_n57_), .C(new_new_n645_), .D(i_5_), .Y(new_new_n852_));
  AN2        g830(.A(new_new_n852_), .B(new_new_n851_), .Y(new_new_n853_));
  NA2        g831(.A(new_new_n180_), .B(new_new_n79_), .Y(new_new_n854_));
  NA2        g832(.A(new_new_n543_), .B(i_4_), .Y(new_new_n855_));
  NA2        g833(.A(new_new_n183_), .B(new_new_n197_), .Y(new_new_n856_));
  OAI220     g834(.A0(new_new_n856_), .A1(new_new_n848_), .B0(new_new_n855_), .B1(new_new_n854_), .Y(new_new_n857_));
  NO4        g835(.A(new_new_n857_), .B(new_new_n853_), .C(new_new_n850_), .D(new_new_n847_), .Y(new_new_n858_));
  NA3        g836(.A(new_new_n858_), .B(new_new_n846_), .C(new_new_n842_), .Y(new_new_n859_));
  NO2        g837(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n860_));
  NA2        g838(.A(i_11_), .B(i_9_), .Y(new_new_n861_));
  NO3        g839(.A(i_12_), .B(new_new_n861_), .C(new_new_n581_), .Y(new_new_n862_));
  AN2        g840(.A(new_new_n862_), .B(new_new_n860_), .Y(new_new_n863_));
  NA2        g841(.A(new_new_n380_), .B(new_new_n173_), .Y(new_new_n864_));
  NA2        g842(.A(new_new_n864_), .B(new_new_n154_), .Y(new_new_n865_));
  NO2        g843(.A(new_new_n861_), .B(new_new_n70_), .Y(new_new_n866_));
  NO2        g844(.A(new_new_n169_), .B(i_0_), .Y(new_new_n867_));
  INV        g845(.A(new_new_n867_), .Y(new_new_n868_));
  NA2        g846(.A(new_new_n455_), .B(new_new_n225_), .Y(new_new_n869_));
  AOI210     g847(.A0(new_new_n359_), .A1(i_4_), .B0(new_new_n394_), .Y(new_new_n870_));
  OAI220     g848(.A0(new_new_n870_), .A1(new_new_n829_), .B0(new_new_n869_), .B1(new_new_n868_), .Y(new_new_n871_));
  NO3        g849(.A(new_new_n871_), .B(new_new_n865_), .C(new_new_n863_), .Y(new_new_n872_));
  NA2        g850(.A(new_new_n635_), .B(new_new_n116_), .Y(new_new_n873_));
  NO2        g851(.A(i_6_), .B(new_new_n873_), .Y(new_new_n874_));
  AOI210     g852(.A0(new_new_n434_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n875_));
  NA2        g853(.A(new_new_n165_), .B(new_new_n97_), .Y(new_new_n876_));
  NOi32      g854(.An(new_new_n875_), .Bn(new_new_n183_), .C(new_new_n876_), .Y(new_new_n877_));
  NA2        g855(.A(new_new_n583_), .B(new_new_n314_), .Y(new_new_n878_));
  NO2        g856(.A(new_new_n878_), .B(new_new_n818_), .Y(new_new_n879_));
  NO3        g857(.A(new_new_n879_), .B(new_new_n877_), .C(new_new_n874_), .Y(new_new_n880_));
  NOi21      g858(.An(i_7_), .B(i_5_), .Y(new_new_n881_));
  NOi31      g859(.An(new_new_n881_), .B(i_0_), .C(new_new_n701_), .Y(new_new_n882_));
  OR2        g860(.A(new_new_n876_), .B(new_new_n493_), .Y(new_new_n883_));
  NO3        g861(.A(new_new_n390_), .B(new_new_n348_), .C(new_new_n344_), .Y(new_new_n884_));
  NO2        g862(.A(new_new_n246_), .B(new_new_n304_), .Y(new_new_n885_));
  INV        g863(.A(new_new_n701_), .Y(new_new_n886_));
  AOI210     g864(.A0(new_new_n886_), .A1(new_new_n885_), .B0(new_new_n884_), .Y(new_new_n887_));
  NA4        g865(.A(new_new_n887_), .B(new_new_n883_), .C(new_new_n880_), .D(new_new_n872_), .Y(new_new_n888_));
  AN2        g866(.A(new_new_n318_), .B(new_new_n314_), .Y(new_new_n889_));
  AN2        g867(.A(new_new_n889_), .B(new_new_n832_), .Y(new_new_n890_));
  NA2        g868(.A(new_new_n890_), .B(i_10_), .Y(new_new_n891_));
  OA210      g869(.A0(new_new_n455_), .A1(new_new_n217_), .B0(new_new_n454_), .Y(new_new_n892_));
  NA3        g870(.A(new_new_n454_), .B(new_new_n397_), .C(new_new_n45_), .Y(new_new_n893_));
  OAI210     g871(.A0(new_new_n840_), .A1(i_6_), .B0(new_new_n893_), .Y(new_new_n894_));
  NA2        g872(.A(new_new_n866_), .B(new_new_n290_), .Y(new_new_n895_));
  NA2        g873(.A(new_new_n182_), .B(new_new_n895_), .Y(new_new_n896_));
  AOI220     g874(.A0(new_new_n896_), .A1(new_new_n455_), .B0(new_new_n894_), .B1(new_new_n70_), .Y(new_new_n897_));
  NO2        g875(.A(new_new_n72_), .B(new_new_n720_), .Y(new_new_n898_));
  AOI210     g876(.A0(new_new_n168_), .A1(new_new_n573_), .B0(new_new_n898_), .Y(new_new_n899_));
  NO2        g877(.A(new_new_n899_), .B(new_new_n47_), .Y(new_new_n900_));
  NO3        g878(.A(new_new_n564_), .B(new_new_n343_), .C(new_new_n24_), .Y(new_new_n901_));
  NO2        g879(.A(new_new_n521_), .B(new_new_n901_), .Y(new_new_n902_));
  NAi21      g880(.An(i_9_), .B(i_5_), .Y(new_new_n903_));
  NO2        g881(.A(new_new_n903_), .B(new_new_n390_), .Y(new_new_n904_));
  NA2        g882(.A(new_new_n904_), .B(new_new_n597_), .Y(new_new_n905_));
  OAI220     g883(.A0(new_new_n905_), .A1(new_new_n80_), .B0(new_new_n902_), .B1(new_new_n166_), .Y(new_new_n906_));
  NO3        g884(.A(new_new_n906_), .B(new_new_n900_), .C(new_new_n497_), .Y(new_new_n907_));
  NA3        g885(.A(new_new_n907_), .B(new_new_n897_), .C(new_new_n891_), .Y(new_new_n908_));
  NO3        g886(.A(new_new_n908_), .B(new_new_n888_), .C(new_new_n859_), .Y(new_new_n909_));
  NO2        g887(.A(i_0_), .B(new_new_n701_), .Y(new_new_n910_));
  AOI210     g888(.A0(new_new_n768_), .A1(new_new_n659_), .B0(new_new_n876_), .Y(new_new_n911_));
  INV        g889(.A(new_new_n911_), .Y(new_new_n912_));
  NA3        g890(.A(new_new_n141_), .B(new_new_n649_), .C(new_new_n70_), .Y(new_new_n913_));
  NO2        g891(.A(new_new_n780_), .B(new_new_n390_), .Y(new_new_n914_));
  NA2        g892(.A(new_new_n810_), .B(i_9_), .Y(new_new_n915_));
  NO2        g893(.A(new_new_n474_), .B(new_new_n915_), .Y(new_new_n916_));
  NA2        g894(.A(new_new_n236_), .B(new_new_n224_), .Y(new_new_n917_));
  AOI210     g895(.A0(new_new_n917_), .A1(new_new_n843_), .B0(new_new_n147_), .Y(new_new_n918_));
  NO3        g896(.A(new_new_n918_), .B(new_new_n916_), .C(new_new_n914_), .Y(new_new_n919_));
  NA3        g897(.A(new_new_n919_), .B(new_new_n913_), .C(new_new_n912_), .Y(new_new_n920_));
  NA2        g898(.A(new_new_n889_), .B(new_new_n360_), .Y(new_new_n921_));
  AOI210     g899(.A0(new_new_n285_), .A1(new_new_n156_), .B0(new_new_n921_), .Y(new_new_n922_));
  NA3        g900(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n923_));
  NA2        g901(.A(i_5_), .B(new_new_n469_), .Y(new_new_n924_));
  AOI210     g902(.A0(new_new_n923_), .A1(new_new_n156_), .B0(new_new_n924_), .Y(new_new_n925_));
  NO2        g903(.A(new_new_n925_), .B(new_new_n922_), .Y(new_new_n926_));
  NA2        g904(.A(new_new_n544_), .B(new_new_n72_), .Y(new_new_n927_));
  NO3        g905(.A(new_new_n204_), .B(new_new_n370_), .C(i_0_), .Y(new_new_n928_));
  OAI210     g906(.A0(new_new_n928_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n929_));
  INV        g907(.A(new_new_n213_), .Y(new_new_n930_));
  OAI220     g908(.A0(new_new_n506_), .A1(new_new_n134_), .B0(i_12_), .B1(new_new_n591_), .Y(new_new_n931_));
  NA3        g909(.A(new_new_n931_), .B(i_7_), .C(new_new_n930_), .Y(new_new_n932_));
  NA4        g910(.A(new_new_n932_), .B(new_new_n929_), .C(new_new_n927_), .D(new_new_n926_), .Y(new_new_n933_));
  INV        g911(.A(new_new_n87_), .Y(new_new_n934_));
  AOI210     g912(.A0(new_new_n934_), .A1(new_new_n910_), .B0(new_new_n103_), .Y(new_new_n935_));
  NA2        g913(.A(new_new_n881_), .B(new_new_n469_), .Y(new_new_n936_));
  NA2        g914(.A(new_new_n335_), .B(new_new_n170_), .Y(new_new_n937_));
  OA220      g915(.A0(new_new_n937_), .A1(new_new_n936_), .B0(new_new_n935_), .B1(i_5_), .Y(new_new_n938_));
  AOI210     g916(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n169_), .Y(new_new_n939_));
  NA2        g917(.A(new_new_n939_), .B(new_new_n892_), .Y(new_new_n940_));
  NA3        g918(.A(i_5_), .B(new_new_n274_), .C(new_new_n224_), .Y(new_new_n941_));
  INV        g919(.A(new_new_n941_), .Y(new_new_n942_));
  NA3        g920(.A(new_new_n376_), .B(new_new_n320_), .C(new_new_n216_), .Y(new_new_n943_));
  OAI210     g921(.A0(new_new_n823_), .A1(new_new_n623_), .B0(new_new_n943_), .Y(new_new_n944_));
  NO2        g922(.A(new_new_n944_), .B(new_new_n942_), .Y(new_new_n945_));
  NA3        g923(.A(new_new_n945_), .B(new_new_n940_), .C(new_new_n938_), .Y(new_new_n946_));
  NA2        g924(.A(new_new_n290_), .B(i_5_), .Y(new_new_n947_));
  NA2        g925(.A(new_new_n762_), .B(new_new_n170_), .Y(new_new_n948_));
  BUFFER     g926(.A(new_new_n147_), .Y(new_new_n949_));
  NO3        g927(.A(new_new_n949_), .B(i_12_), .C(new_new_n623_), .Y(new_new_n950_));
  NA2        g928(.A(new_new_n950_), .B(new_new_n213_), .Y(new_new_n951_));
  NA3        g929(.A(new_new_n92_), .B(new_new_n548_), .C(i_11_), .Y(new_new_n952_));
  NO2        g930(.A(new_new_n952_), .B(new_new_n149_), .Y(new_new_n953_));
  NA2        g931(.A(new_new_n881_), .B(new_new_n452_), .Y(new_new_n954_));
  OAI220     g932(.A0(i_7_), .A1(new_new_n947_), .B0(new_new_n954_), .B1(i_1_), .Y(new_new_n955_));
  AOI210     g933(.A0(new_new_n955_), .A1(new_new_n867_), .B0(new_new_n953_), .Y(new_new_n956_));
  NA3        g934(.A(new_new_n956_), .B(new_new_n951_), .C(new_new_n948_), .Y(new_new_n957_));
  NO4        g935(.A(new_new_n957_), .B(new_new_n946_), .C(new_new_n933_), .D(new_new_n920_), .Y(new_new_n958_));
  OAI210     g936(.A0(new_new_n783_), .A1(new_new_n776_), .B0(new_new_n37_), .Y(new_new_n959_));
  NA3        g937(.A(new_new_n875_), .B(new_new_n356_), .C(i_5_), .Y(new_new_n960_));
  NA3        g938(.A(new_new_n960_), .B(new_new_n959_), .C(new_new_n586_), .Y(new_new_n961_));
  NA2        g939(.A(new_new_n961_), .B(new_new_n201_), .Y(new_new_n962_));
  NA2        g940(.A(new_new_n181_), .B(new_new_n183_), .Y(new_new_n963_));
  AO210      g941(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n963_), .Y(new_new_n964_));
  OAI210     g942(.A0(new_new_n590_), .A1(new_new_n588_), .B0(new_new_n303_), .Y(new_new_n965_));
  NAi31      g943(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n966_));
  NO2        g944(.A(new_new_n67_), .B(new_new_n966_), .Y(new_new_n967_));
  INV        g945(.A(new_new_n967_), .Y(new_new_n968_));
  NA3        g946(.A(new_new_n968_), .B(new_new_n965_), .C(new_new_n964_), .Y(new_new_n969_));
  NO2        g947(.A(new_new_n444_), .B(new_new_n252_), .Y(new_new_n970_));
  NO2        g948(.A(new_new_n970_), .B(new_new_n845_), .Y(new_new_n971_));
  OAI210     g949(.A0(new_new_n952_), .A1(new_new_n143_), .B0(new_new_n971_), .Y(new_new_n972_));
  AOI210     g950(.A0(new_new_n969_), .A1(new_new_n48_), .B0(new_new_n972_), .Y(new_new_n973_));
  AOI210     g951(.A0(new_new_n973_), .A1(new_new_n962_), .B0(new_new_n70_), .Y(new_new_n974_));
  NO2        g952(.A(new_new_n541_), .B(new_new_n366_), .Y(new_new_n975_));
  NO2        g953(.A(new_new_n975_), .B(new_new_n726_), .Y(new_new_n976_));
  AOI210     g954(.A0(new_new_n939_), .A1(i_5_), .B0(new_new_n882_), .Y(new_new_n977_));
  NO2        g955(.A(new_new_n977_), .B(new_new_n650_), .Y(new_new_n978_));
  INV        g956(.A(new_new_n56_), .Y(new_new_n979_));
  AOI220     g957(.A0(new_new_n979_), .A1(new_new_n73_), .B0(new_new_n332_), .B1(new_new_n244_), .Y(new_new_n980_));
  NO2        g958(.A(new_new_n980_), .B(new_new_n230_), .Y(new_new_n981_));
  NO2        g959(.A(new_new_n981_), .B(new_new_n978_), .Y(new_new_n982_));
  OAI210     g960(.A0(new_new_n254_), .A1(new_new_n152_), .B0(new_new_n83_), .Y(new_new_n983_));
  NA3        g961(.A(new_new_n730_), .B(new_new_n274_), .C(new_new_n77_), .Y(new_new_n984_));
  AOI210     g962(.A0(new_new_n984_), .A1(new_new_n983_), .B0(i_11_), .Y(new_new_n985_));
  OAI210     g963(.A0(new_new_n1004_), .A1(new_new_n875_), .B0(new_new_n201_), .Y(new_new_n986_));
  NA2        g964(.A(new_new_n158_), .B(i_5_), .Y(new_new_n987_));
  AOI210     g965(.A0(new_new_n986_), .A1(new_new_n740_), .B0(new_new_n987_), .Y(new_new_n988_));
  NO3        g966(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n989_));
  NA2        g967(.A(new_new_n292_), .B(new_new_n989_), .Y(new_new_n990_));
  NO2        g968(.A(new_new_n990_), .B(new_new_n701_), .Y(new_new_n991_));
  NO3        g969(.A(new_new_n903_), .B(new_new_n458_), .C(new_new_n243_), .Y(new_new_n992_));
  NO2        g970(.A(new_new_n992_), .B(new_new_n538_), .Y(new_new_n993_));
  INV        g971(.A(new_new_n349_), .Y(new_new_n994_));
  AOI210     g972(.A0(new_new_n994_), .A1(new_new_n993_), .B0(new_new_n41_), .Y(new_new_n995_));
  NO4        g973(.A(new_new_n995_), .B(new_new_n991_), .C(new_new_n988_), .D(new_new_n985_), .Y(new_new_n996_));
  OAI210     g974(.A0(new_new_n982_), .A1(i_4_), .B0(new_new_n996_), .Y(new_new_n997_));
  NO3        g975(.A(new_new_n997_), .B(new_new_n976_), .C(new_new_n974_), .Y(new_new_n998_));
  NA4        g976(.A(new_new_n998_), .B(new_new_n958_), .C(new_new_n909_), .D(new_new_n835_), .Y(mai4));
  INV        g977(.A(new_new_n676_), .Y(new_new_n1002_));
  INV        g978(.A(i_2_), .Y(new_new_n1003_));
  INV        g979(.A(i_12_), .Y(new_new_n1004_));
endmodule


