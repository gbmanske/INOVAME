//Benchmark atmr_max1024_476_0.125

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n393_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n432_, men_men_n433_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO4        o012(.A(ori_ori_n28_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  AN2        o021(.A(x8), .B(x7), .Y(ori_ori_n38_));
  NA3        o022(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o023(.A(x4), .B(x3), .Y(ori_ori_n40_));
  AOI210     o024(.A0(ori_ori_n39_), .A1(ori_ori_n23_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o025(.A(x2), .B(x0), .Y(ori_ori_n42_));
  INV        o026(.A(x3), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  INV        o028(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n42_), .Y(ori_ori_n47_));
  INV        o031(.A(x4), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(x2), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n50_), .A1(ori_ori_n20_), .B0(ori_ori_n47_), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n52_));
  AOI220     o036(.A0(ori_ori_n52_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n53_));
  INV        o037(.A(x2), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  OAI210     o041(.A0(ori_ori_n53_), .A1(ori_ori_n32_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  NO3        o042(.A(ori_ori_n58_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori01));
  NA2        o043(.A(x8), .B(x7), .Y(ori_ori_n60_));
  NA2        o044(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n61_));
  INV        o045(.A(x9), .Y(ori_ori_n62_));
  NO2        o046(.A(x7), .B(x6), .Y(ori_ori_n63_));
  NO2        o047(.A(ori_ori_n61_), .B(x5), .Y(ori_ori_n64_));
  NO2        o048(.A(x8), .B(x2), .Y(ori_ori_n65_));
  INV        o049(.A(ori_ori_n65_), .Y(ori_ori_n66_));
  NO2        o050(.A(ori_ori_n66_), .B(x1), .Y(ori_ori_n67_));
  AN2        o051(.A(ori_ori_n67_), .B(ori_ori_n63_), .Y(ori_ori_n68_));
  OAI210     o052(.A0(ori_ori_n44_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n56_), .A1(ori_ori_n20_), .B0(ori_ori_n69_), .Y(ori_ori_n70_));
  NO2        o054(.A(ori_ori_n70_), .B(ori_ori_n68_), .Y(ori_ori_n71_));
  NA2        o055(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n73_));
  OAI210     o057(.A0(ori_ori_n73_), .A1(ori_ori_n56_), .B0(x0), .Y(ori_ori_n74_));
  NA2        o058(.A(x5), .B(x3), .Y(ori_ori_n75_));
  NO2        o059(.A(x8), .B(x6), .Y(ori_ori_n76_));
  NO4        o060(.A(ori_ori_n76_), .B(ori_ori_n75_), .C(ori_ori_n63_), .D(ori_ori_n54_), .Y(ori_ori_n77_));
  NAi21      o061(.An(x4), .B(x3), .Y(ori_ori_n78_));
  INV        o062(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NO2        o063(.A(ori_ori_n79_), .B(ori_ori_n22_), .Y(ori_ori_n80_));
  NO2        o064(.A(x4), .B(x2), .Y(ori_ori_n81_));
  NO2        o065(.A(ori_ori_n81_), .B(x3), .Y(ori_ori_n82_));
  NO3        o066(.A(ori_ori_n82_), .B(ori_ori_n80_), .C(ori_ori_n18_), .Y(ori_ori_n83_));
  NO3        o067(.A(ori_ori_n83_), .B(ori_ori_n77_), .C(ori_ori_n74_), .Y(ori_ori_n84_));
  NA2        o068(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n85_));
  NO2        o069(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n86_));
  INV        o070(.A(x8), .Y(ori_ori_n87_));
  NA2        o071(.A(x2), .B(x1), .Y(ori_ori_n88_));
  INV        o072(.A(ori_ori_n86_), .Y(ori_ori_n89_));
  NO2        o073(.A(ori_ori_n89_), .B(ori_ori_n26_), .Y(ori_ori_n90_));
  AOI210     o074(.A0(ori_ori_n56_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n91_));
  OAI210     o075(.A0(ori_ori_n45_), .A1(ori_ori_n37_), .B0(ori_ori_n48_), .Y(ori_ori_n92_));
  NO3        o076(.A(ori_ori_n92_), .B(ori_ori_n91_), .C(ori_ori_n90_), .Y(ori_ori_n93_));
  NA2        o077(.A(x4), .B(ori_ori_n43_), .Y(ori_ori_n94_));
  NO2        o078(.A(ori_ori_n48_), .B(ori_ori_n54_), .Y(ori_ori_n95_));
  OAI210     o079(.A0(ori_ori_n95_), .A1(ori_ori_n43_), .B0(ori_ori_n18_), .Y(ori_ori_n96_));
  AOI210     o080(.A0(ori_ori_n94_), .A1(ori_ori_n52_), .B0(ori_ori_n96_), .Y(ori_ori_n97_));
  NO2        o081(.A(x3), .B(x2), .Y(ori_ori_n98_));
  NA3        o082(.A(ori_ori_n98_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n99_));
  INV        o083(.A(ori_ori_n99_), .Y(ori_ori_n100_));
  NA2        o084(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n101_));
  OAI210     o085(.A0(ori_ori_n101_), .A1(ori_ori_n40_), .B0(ori_ori_n17_), .Y(ori_ori_n102_));
  NO4        o086(.A(ori_ori_n102_), .B(ori_ori_n100_), .C(ori_ori_n97_), .D(ori_ori_n93_), .Y(ori_ori_n103_));
  AO210      o087(.A0(ori_ori_n84_), .A1(ori_ori_n72_), .B0(ori_ori_n103_), .Y(ori02));
  NO2        o088(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n105_));
  NO2        o089(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n106_));
  NA2        o090(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n107_));
  OR2        o091(.A(x8), .B(x0), .Y(ori_ori_n108_));
  INV        o092(.A(ori_ori_n108_), .Y(ori_ori_n109_));
  NAi21      o093(.An(x2), .B(x8), .Y(ori_ori_n110_));
  NO2        o094(.A(x4), .B(x1), .Y(ori_ori_n111_));
  NA3        o095(.A(ori_ori_n111_), .B(x2), .C(ori_ori_n60_), .Y(ori_ori_n112_));
  NOi21      o096(.An(x0), .B(x1), .Y(ori_ori_n113_));
  NO3        o097(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n114_));
  NOi21      o098(.An(x0), .B(x4), .Y(ori_ori_n115_));
  NAi21      o099(.An(x8), .B(x7), .Y(ori_ori_n116_));
  NO2        o100(.A(ori_ori_n116_), .B(ori_ori_n62_), .Y(ori_ori_n117_));
  NA2        o101(.A(ori_ori_n117_), .B(ori_ori_n115_), .Y(ori_ori_n118_));
  AOI210     o102(.A0(ori_ori_n118_), .A1(ori_ori_n112_), .B0(ori_ori_n75_), .Y(ori_ori_n119_));
  NO2        o103(.A(x5), .B(ori_ori_n48_), .Y(ori_ori_n120_));
  NA2        o104(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n121_));
  AOI210     o105(.A0(ori_ori_n121_), .A1(ori_ori_n101_), .B0(ori_ori_n107_), .Y(ori_ori_n122_));
  OAI210     o106(.A0(ori_ori_n122_), .A1(ori_ori_n35_), .B0(ori_ori_n120_), .Y(ori_ori_n123_));
  NAi21      o107(.An(x0), .B(x4), .Y(ori_ori_n124_));
  NO2        o108(.A(x7), .B(x0), .Y(ori_ori_n125_));
  NO2        o109(.A(ori_ori_n81_), .B(ori_ori_n95_), .Y(ori_ori_n126_));
  NO2        o110(.A(ori_ori_n126_), .B(x3), .Y(ori_ori_n127_));
  NA2        o111(.A(ori_ori_n125_), .B(ori_ori_n127_), .Y(ori_ori_n128_));
  NO2        o112(.A(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n129_));
  NA2        o113(.A(x5), .B(x0), .Y(ori_ori_n130_));
  NO2        o114(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n131_));
  NA2        o115(.A(ori_ori_n131_), .B(ori_ori_n129_), .Y(ori_ori_n132_));
  NA4        o116(.A(ori_ori_n132_), .B(ori_ori_n128_), .C(ori_ori_n123_), .D(ori_ori_n36_), .Y(ori_ori_n133_));
  NO2        o117(.A(ori_ori_n133_), .B(ori_ori_n119_), .Y(ori_ori_n134_));
  NO3        o118(.A(ori_ori_n75_), .B(ori_ori_n73_), .C(ori_ori_n24_), .Y(ori_ori_n135_));
  NO2        o119(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n136_));
  NA2        o120(.A(x7), .B(x3), .Y(ori_ori_n137_));
  NO2        o121(.A(ori_ori_n94_), .B(x5), .Y(ori_ori_n138_));
  NO2        o122(.A(x9), .B(x7), .Y(ori_ori_n139_));
  NOi21      o123(.An(x8), .B(x0), .Y(ori_ori_n140_));
  NO2        o124(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n141_));
  INV        o125(.A(x7), .Y(ori_ori_n142_));
  NA2        o126(.A(ori_ori_n142_), .B(ori_ori_n18_), .Y(ori_ori_n143_));
  AOI220     o127(.A0(ori_ori_n143_), .A1(ori_ori_n141_), .B0(ori_ori_n105_), .B1(ori_ori_n38_), .Y(ori_ori_n144_));
  NO2        o128(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n145_));
  NO2        o129(.A(ori_ori_n145_), .B(ori_ori_n115_), .Y(ori_ori_n146_));
  NO2        o130(.A(ori_ori_n146_), .B(ori_ori_n144_), .Y(ori_ori_n147_));
  INV        o131(.A(ori_ori_n147_), .Y(ori_ori_n148_));
  OAI210     o132(.A0(ori_ori_n137_), .A1(ori_ori_n50_), .B0(ori_ori_n148_), .Y(ori_ori_n149_));
  NA2        o133(.A(x5), .B(x1), .Y(ori_ori_n150_));
  INV        o134(.A(ori_ori_n150_), .Y(ori_ori_n151_));
  AOI210     o135(.A0(ori_ori_n151_), .A1(ori_ori_n115_), .B0(ori_ori_n36_), .Y(ori_ori_n152_));
  NAi21      o136(.An(x2), .B(x7), .Y(ori_ori_n153_));
  NO2        o137(.A(ori_ori_n153_), .B(ori_ori_n48_), .Y(ori_ori_n154_));
  NA2        o138(.A(ori_ori_n154_), .B(ori_ori_n64_), .Y(ori_ori_n155_));
  NAi31      o139(.An(ori_ori_n75_), .B(ori_ori_n38_), .C(ori_ori_n35_), .Y(ori_ori_n156_));
  NA3        o140(.A(ori_ori_n156_), .B(ori_ori_n155_), .C(ori_ori_n152_), .Y(ori_ori_n157_));
  NO3        o141(.A(ori_ori_n157_), .B(ori_ori_n149_), .C(ori_ori_n135_), .Y(ori_ori_n158_));
  NO2        o142(.A(ori_ori_n158_), .B(ori_ori_n134_), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n130_), .B(ori_ori_n126_), .Y(ori_ori_n160_));
  NA2        o144(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n161_));
  NA2        o145(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n162_));
  NA3        o146(.A(ori_ori_n162_), .B(ori_ori_n161_), .C(ori_ori_n24_), .Y(ori_ori_n163_));
  AN2        o147(.A(ori_ori_n163_), .B(ori_ori_n131_), .Y(ori_ori_n164_));
  NA2        o148(.A(x8), .B(x0), .Y(ori_ori_n165_));
  NO2        o149(.A(ori_ori_n142_), .B(ori_ori_n25_), .Y(ori_ori_n166_));
  NO2        o150(.A(ori_ori_n113_), .B(x4), .Y(ori_ori_n167_));
  NA2        o151(.A(ori_ori_n167_), .B(ori_ori_n166_), .Y(ori_ori_n168_));
  AOI210     o152(.A0(ori_ori_n165_), .A1(ori_ori_n121_), .B0(ori_ori_n168_), .Y(ori_ori_n169_));
  NA2        o153(.A(x2), .B(x0), .Y(ori_ori_n170_));
  NA2        o154(.A(x4), .B(x1), .Y(ori_ori_n171_));
  NAi21      o155(.An(ori_ori_n111_), .B(ori_ori_n171_), .Y(ori_ori_n172_));
  NOi31      o156(.An(ori_ori_n172_), .B(ori_ori_n145_), .C(ori_ori_n170_), .Y(ori_ori_n173_));
  NO4        o157(.A(ori_ori_n173_), .B(ori_ori_n169_), .C(ori_ori_n164_), .D(ori_ori_n160_), .Y(ori_ori_n174_));
  NO2        o158(.A(ori_ori_n174_), .B(ori_ori_n43_), .Y(ori_ori_n175_));
  NO2        o159(.A(ori_ori_n163_), .B(ori_ori_n73_), .Y(ori_ori_n176_));
  INV        o160(.A(ori_ori_n120_), .Y(ori_ori_n177_));
  NO2        o161(.A(ori_ori_n101_), .B(ori_ori_n17_), .Y(ori_ori_n178_));
  AOI210     o162(.A0(ori_ori_n35_), .A1(ori_ori_n87_), .B0(ori_ori_n178_), .Y(ori_ori_n179_));
  NO3        o163(.A(ori_ori_n179_), .B(ori_ori_n177_), .C(x7), .Y(ori_ori_n180_));
  NA3        o164(.A(ori_ori_n172_), .B(ori_ori_n177_), .C(ori_ori_n42_), .Y(ori_ori_n181_));
  OAI210     o165(.A0(ori_ori_n162_), .A1(ori_ori_n126_), .B0(ori_ori_n181_), .Y(ori_ori_n182_));
  NO3        o166(.A(ori_ori_n182_), .B(ori_ori_n180_), .C(ori_ori_n176_), .Y(ori_ori_n183_));
  NO2        o167(.A(ori_ori_n183_), .B(x3), .Y(ori_ori_n184_));
  NO3        o168(.A(ori_ori_n184_), .B(ori_ori_n175_), .C(ori_ori_n159_), .Y(ori03));
  NO2        o169(.A(ori_ori_n48_), .B(x3), .Y(ori_ori_n186_));
  NO2        o170(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n187_));
  NO2        o171(.A(ori_ori_n75_), .B(x6), .Y(ori_ori_n188_));
  NA2        o172(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n189_));
  NO2        o173(.A(ori_ori_n189_), .B(x4), .Y(ori_ori_n190_));
  NO2        o174(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n191_));
  AN2        o175(.A(ori_ori_n188_), .B(ori_ori_n55_), .Y(ori_ori_n192_));
  INV        o176(.A(ori_ori_n192_), .Y(ori_ori_n193_));
  NA2        o177(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n194_));
  NO2        o178(.A(ori_ori_n194_), .B(ori_ori_n189_), .Y(ori_ori_n195_));
  INV        o179(.A(ori_ori_n195_), .Y(ori_ori_n196_));
  NO3        o180(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n197_));
  NO2        o181(.A(x5), .B(x1), .Y(ori_ori_n198_));
  NO2        o182(.A(ori_ori_n194_), .B(ori_ori_n161_), .Y(ori_ori_n199_));
  NO3        o183(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n200_));
  NO2        o184(.A(ori_ori_n200_), .B(ori_ori_n199_), .Y(ori_ori_n201_));
  INV        o185(.A(ori_ori_n201_), .Y(ori_ori_n202_));
  AOI220     o186(.A0(ori_ori_n202_), .A1(ori_ori_n48_), .B0(ori_ori_n197_), .B1(ori_ori_n120_), .Y(ori_ori_n203_));
  NA3        o187(.A(ori_ori_n203_), .B(ori_ori_n196_), .C(ori_ori_n193_), .Y(ori_ori_n204_));
  NO2        o188(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n205_));
  NA2        o189(.A(ori_ori_n205_), .B(ori_ori_n19_), .Y(ori_ori_n206_));
  NO2        o190(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n207_));
  NO2        o191(.A(ori_ori_n207_), .B(x6), .Y(ori_ori_n208_));
  NOi21      o192(.An(ori_ori_n81_), .B(ori_ori_n208_), .Y(ori_ori_n209_));
  NA2        o193(.A(ori_ori_n207_), .B(x6), .Y(ori_ori_n210_));
  AOI210     o194(.A0(ori_ori_n210_), .A1(ori_ori_n209_), .B0(ori_ori_n142_), .Y(ori_ori_n211_));
  AO210      o195(.A0(ori_ori_n211_), .A1(ori_ori_n206_), .B0(ori_ori_n166_), .Y(ori_ori_n212_));
  NA2        o196(.A(ori_ori_n43_), .B(ori_ori_n54_), .Y(ori_ori_n213_));
  NO2        o197(.A(ori_ori_n213_), .B(ori_ori_n25_), .Y(ori_ori_n214_));
  NO2        o198(.A(ori_ori_n171_), .B(x6), .Y(ori_ori_n215_));
  AOI220     o199(.A0(ori_ori_n215_), .A1(ori_ori_n214_), .B0(ori_ori_n131_), .B1(ori_ori_n86_), .Y(ori_ori_n216_));
  NA2        o200(.A(x6), .B(ori_ori_n48_), .Y(ori_ori_n217_));
  OAI210     o201(.A0(ori_ori_n109_), .A1(ori_ori_n76_), .B0(x4), .Y(ori_ori_n218_));
  AOI210     o202(.A0(ori_ori_n218_), .A1(ori_ori_n217_), .B0(ori_ori_n75_), .Y(ori_ori_n219_));
  NO2        o203(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n220_));
  NO2        o204(.A(ori_ori_n150_), .B(ori_ori_n43_), .Y(ori_ori_n221_));
  OAI210     o205(.A0(ori_ori_n221_), .A1(ori_ori_n199_), .B0(ori_ori_n220_), .Y(ori_ori_n222_));
  NA3        o206(.A(ori_ori_n194_), .B(ori_ori_n120_), .C(x6), .Y(ori_ori_n223_));
  INV        o207(.A(ori_ori_n64_), .Y(ori_ori_n224_));
  NA3        o208(.A(ori_ori_n224_), .B(ori_ori_n223_), .C(ori_ori_n222_), .Y(ori_ori_n225_));
  OAI210     o209(.A0(ori_ori_n225_), .A1(ori_ori_n219_), .B0(x2), .Y(ori_ori_n226_));
  NA3        o210(.A(ori_ori_n226_), .B(ori_ori_n216_), .C(ori_ori_n212_), .Y(ori_ori_n227_));
  AOI210     o211(.A0(ori_ori_n204_), .A1(x8), .B0(ori_ori_n227_), .Y(ori_ori_n228_));
  NO2        o212(.A(ori_ori_n87_), .B(x3), .Y(ori_ori_n229_));
  NA2        o213(.A(ori_ori_n229_), .B(ori_ori_n190_), .Y(ori_ori_n230_));
  NO3        o214(.A(ori_ori_n85_), .B(ori_ori_n76_), .C(ori_ori_n25_), .Y(ori_ori_n231_));
  AOI210     o215(.A0(ori_ori_n208_), .A1(ori_ori_n145_), .B0(ori_ori_n231_), .Y(ori_ori_n232_));
  AOI210     o216(.A0(ori_ori_n232_), .A1(ori_ori_n230_), .B0(x2), .Y(ori_ori_n233_));
  AOI220     o217(.A0(ori_ori_n190_), .A1(ori_ori_n178_), .B0(x2), .B1(ori_ori_n64_), .Y(ori_ori_n234_));
  NA2        o218(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n235_));
  NA2        o219(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n236_));
  NA2        o220(.A(ori_ori_n194_), .B(x6), .Y(ori_ori_n237_));
  NO2        o221(.A(ori_ori_n194_), .B(x6), .Y(ori_ori_n238_));
  INV        o222(.A(ori_ori_n238_), .Y(ori_ori_n239_));
  NA3        o223(.A(ori_ori_n239_), .B(ori_ori_n237_), .C(ori_ori_n136_), .Y(ori_ori_n240_));
  NA3        o224(.A(ori_ori_n240_), .B(ori_ori_n234_), .C(ori_ori_n142_), .Y(ori_ori_n241_));
  NO2        o225(.A(ori_ori_n130_), .B(ori_ori_n18_), .Y(ori_ori_n242_));
  NA2        o226(.A(x6), .B(x2), .Y(ori_ori_n243_));
  NA2        o227(.A(x9), .B(ori_ori_n43_), .Y(ori_ori_n244_));
  NO2        o228(.A(ori_ori_n244_), .B(ori_ori_n189_), .Y(ori_ori_n245_));
  OR3        o229(.A(ori_ori_n245_), .B(ori_ori_n188_), .C(ori_ori_n138_), .Y(ori_ori_n246_));
  NA2        o230(.A(x4), .B(x0), .Y(ori_ori_n247_));
  NA2        o231(.A(ori_ori_n246_), .B(ori_ori_n42_), .Y(ori_ori_n248_));
  NO2        o232(.A(ori_ori_n248_), .B(x8), .Y(ori_ori_n249_));
  INV        o233(.A(ori_ori_n235_), .Y(ori_ori_n250_));
  OAI210     o234(.A0(ori_ori_n242_), .A1(ori_ori_n198_), .B0(ori_ori_n250_), .Y(ori_ori_n251_));
  INV        o235(.A(ori_ori_n165_), .Y(ori_ori_n252_));
  OAI210     o236(.A0(ori_ori_n252_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n253_));
  AOI210     o237(.A0(ori_ori_n253_), .A1(ori_ori_n251_), .B0(ori_ori_n213_), .Y(ori_ori_n254_));
  NO4        o238(.A(ori_ori_n254_), .B(ori_ori_n249_), .C(ori_ori_n241_), .D(ori_ori_n233_), .Y(ori_ori_n255_));
  NA2        o239(.A(ori_ori_n238_), .B(x2), .Y(ori_ori_n256_));
  OAI210     o240(.A0(ori_ori_n252_), .A1(x6), .B0(ori_ori_n44_), .Y(ori_ori_n257_));
  AOI210     o241(.A0(ori_ori_n257_), .A1(ori_ori_n256_), .B0(ori_ori_n177_), .Y(ori_ori_n258_));
  NOi21      o242(.An(ori_ori_n243_), .B(ori_ori_n17_), .Y(ori_ori_n259_));
  NA3        o243(.A(ori_ori_n259_), .B(ori_ori_n198_), .C(ori_ori_n40_), .Y(ori_ori_n260_));
  AOI210     o244(.A0(ori_ori_n36_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n261_));
  NA3        o245(.A(ori_ori_n261_), .B(ori_ori_n151_), .C(ori_ori_n32_), .Y(ori_ori_n262_));
  NA2        o246(.A(x3), .B(x2), .Y(ori_ori_n263_));
  AOI220     o247(.A0(ori_ori_n263_), .A1(ori_ori_n213_), .B0(ori_ori_n262_), .B1(ori_ori_n260_), .Y(ori_ori_n264_));
  NAi21      o248(.An(x4), .B(x0), .Y(ori_ori_n265_));
  NO3        o249(.A(ori_ori_n265_), .B(ori_ori_n44_), .C(x2), .Y(ori_ori_n266_));
  OAI210     o250(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n266_), .Y(ori_ori_n267_));
  OAI220     o251(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n268_));
  NO2        o252(.A(ori_ori_n261_), .B(ori_ori_n259_), .Y(ori_ori_n269_));
  AOI220     o253(.A0(ori_ori_n269_), .A1(ori_ori_n79_), .B0(ori_ori_n268_), .B1(ori_ori_n31_), .Y(ori_ori_n270_));
  AOI210     o254(.A0(ori_ori_n270_), .A1(ori_ori_n267_), .B0(ori_ori_n25_), .Y(ori_ori_n271_));
  NO2        o255(.A(ori_ori_n261_), .B(ori_ori_n259_), .Y(ori_ori_n272_));
  INV        o256(.A(ori_ori_n199_), .Y(ori_ori_n273_));
  NA2        o257(.A(ori_ori_n36_), .B(ori_ori_n43_), .Y(ori_ori_n274_));
  OR2        o258(.A(ori_ori_n274_), .B(ori_ori_n247_), .Y(ori_ori_n275_));
  OAI220     o259(.A0(ori_ori_n275_), .A1(ori_ori_n150_), .B0(ori_ori_n217_), .B1(ori_ori_n273_), .Y(ori_ori_n276_));
  AO210      o260(.A0(ori_ori_n272_), .A1(ori_ori_n138_), .B0(ori_ori_n276_), .Y(ori_ori_n277_));
  NO4        o261(.A(ori_ori_n277_), .B(ori_ori_n271_), .C(ori_ori_n264_), .D(ori_ori_n258_), .Y(ori_ori_n278_));
  OAI210     o262(.A0(ori_ori_n255_), .A1(ori_ori_n228_), .B0(ori_ori_n278_), .Y(ori04));
  NO2        o263(.A(x2), .B(x1), .Y(ori_ori_n280_));
  OAI210     o264(.A0(ori_ori_n236_), .A1(ori_ori_n280_), .B0(ori_ori_n36_), .Y(ori_ori_n281_));
  INV        o265(.A(ori_ori_n265_), .Y(ori_ori_n282_));
  OAI210     o266(.A0(ori_ori_n54_), .A1(ori_ori_n282_), .B0(ori_ori_n229_), .Y(ori_ori_n283_));
  NO2        o267(.A(ori_ori_n263_), .B(ori_ori_n191_), .Y(ori_ori_n284_));
  NA2        o268(.A(x9), .B(x0), .Y(ori_ori_n285_));
  AOI210     o269(.A0(ori_ori_n85_), .A1(ori_ori_n73_), .B0(ori_ori_n285_), .Y(ori_ori_n286_));
  OAI210     o270(.A0(ori_ori_n286_), .A1(ori_ori_n284_), .B0(ori_ori_n87_), .Y(ori_ori_n287_));
  NA3        o271(.A(ori_ori_n287_), .B(x6), .C(ori_ori_n283_), .Y(ori_ori_n288_));
  NA2        o272(.A(ori_ori_n288_), .B(ori_ori_n281_), .Y(ori_ori_n289_));
  OAI210     o273(.A0(ori_ori_n108_), .A1(ori_ori_n101_), .B0(ori_ori_n165_), .Y(ori_ori_n290_));
  NA3        o274(.A(ori_ori_n290_), .B(x6), .C(x3), .Y(ori_ori_n291_));
  NOi21      o275(.An(ori_ori_n140_), .B(ori_ori_n121_), .Y(ori_ori_n292_));
  NA2        o276(.A(ori_ori_n292_), .B(x6), .Y(ori_ori_n293_));
  NA2        o277(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n294_));
  OAI210     o278(.A0(ori_ori_n101_), .A1(ori_ori_n17_), .B0(ori_ori_n294_), .Y(ori_ori_n295_));
  NA2        o279(.A(ori_ori_n295_), .B(ori_ori_n76_), .Y(ori_ori_n296_));
  NA3        o280(.A(ori_ori_n296_), .B(ori_ori_n293_), .C(ori_ori_n291_), .Y(ori_ori_n297_));
  OAI210     o281(.A0(ori_ori_n106_), .A1(x3), .B0(ori_ori_n266_), .Y(ori_ori_n298_));
  NA2        o282(.A(ori_ori_n197_), .B(ori_ori_n81_), .Y(ori_ori_n299_));
  NA3        o283(.A(ori_ori_n299_), .B(ori_ori_n298_), .C(ori_ori_n142_), .Y(ori_ori_n300_));
  AOI210     o284(.A0(ori_ori_n297_), .A1(x4), .B0(ori_ori_n300_), .Y(ori_ori_n301_));
  XO2        o285(.A(x4), .B(x0), .Y(ori_ori_n302_));
  NA2        o286(.A(x4), .B(ori_ori_n88_), .Y(ori_ori_n303_));
  NO2        o287(.A(ori_ori_n303_), .B(x3), .Y(ori_ori_n304_));
  INV        o288(.A(ori_ori_n88_), .Y(ori_ori_n305_));
  NO2        o289(.A(ori_ori_n87_), .B(x4), .Y(ori_ori_n306_));
  AOI220     o290(.A0(ori_ori_n306_), .A1(ori_ori_n44_), .B0(ori_ori_n115_), .B1(ori_ori_n305_), .Y(ori_ori_n307_));
  NO2        o291(.A(ori_ori_n302_), .B(x2), .Y(ori_ori_n308_));
  INV        o292(.A(ori_ori_n308_), .Y(ori_ori_n309_));
  NA4        o293(.A(ori_ori_n309_), .B(ori_ori_n307_), .C(ori_ori_n206_), .D(x6), .Y(ori_ori_n310_));
  NO2        o294(.A(ori_ori_n140_), .B(ori_ori_n78_), .Y(ori_ori_n311_));
  NO2        o295(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n312_));
  NOi21      o296(.An(ori_ori_n111_), .B(ori_ori_n27_), .Y(ori_ori_n313_));
  AOI210     o297(.A0(ori_ori_n312_), .A1(ori_ori_n311_), .B0(ori_ori_n313_), .Y(ori_ori_n314_));
  OAI210     o298(.A0(ori_ori_n265_), .A1(ori_ori_n62_), .B0(ori_ori_n314_), .Y(ori_ori_n315_));
  OAI220     o299(.A0(ori_ori_n315_), .A1(x6), .B0(ori_ori_n310_), .B1(ori_ori_n304_), .Y(ori_ori_n316_));
  OAI210     o300(.A0(x6), .A1(ori_ori_n48_), .B0(ori_ori_n42_), .Y(ori_ori_n317_));
  OAI210     o301(.A0(ori_ori_n317_), .A1(ori_ori_n87_), .B0(ori_ori_n275_), .Y(ori_ori_n318_));
  AOI210     o302(.A0(ori_ori_n318_), .A1(ori_ori_n18_), .B0(ori_ori_n142_), .Y(ori_ori_n319_));
  AO220      o303(.A0(ori_ori_n319_), .A1(ori_ori_n316_), .B0(ori_ori_n301_), .B1(ori_ori_n289_), .Y(ori_ori_n320_));
  NA2        o304(.A(ori_ori_n312_), .B(x6), .Y(ori_ori_n321_));
  AOI210     o305(.A0(x6), .A1(x1), .B0(ori_ori_n141_), .Y(ori_ori_n322_));
  NA2        o306(.A(ori_ori_n306_), .B(x0), .Y(ori_ori_n323_));
  NA2        o307(.A(ori_ori_n81_), .B(x6), .Y(ori_ori_n324_));
  OAI210     o308(.A0(ori_ori_n323_), .A1(ori_ori_n322_), .B0(ori_ori_n324_), .Y(ori_ori_n325_));
  AOI220     o309(.A0(ori_ori_n325_), .A1(ori_ori_n321_), .B0(ori_ori_n200_), .B1(ori_ori_n49_), .Y(ori_ori_n326_));
  NA2        o310(.A(ori_ori_n326_), .B(ori_ori_n320_), .Y(ori_ori_n327_));
  AOI210     o311(.A0(ori_ori_n187_), .A1(x8), .B0(ori_ori_n106_), .Y(ori_ori_n328_));
  NA2        o312(.A(ori_ori_n328_), .B(ori_ori_n294_), .Y(ori_ori_n329_));
  NA3        o313(.A(ori_ori_n329_), .B(ori_ori_n186_), .C(ori_ori_n142_), .Y(ori_ori_n330_));
  AO220      o314(.A0(x4), .A1(ori_ori_n139_), .B0(ori_ori_n105_), .B1(x4), .Y(ori_ori_n331_));
  NA3        o315(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n332_));
  NA2        o316(.A(ori_ori_n205_), .B(x0), .Y(ori_ori_n333_));
  OAI220     o317(.A0(ori_ori_n333_), .A1(x2), .B0(ori_ori_n332_), .B1(ori_ori_n305_), .Y(ori_ori_n334_));
  AOI210     o318(.A0(ori_ori_n331_), .A1(ori_ori_n109_), .B0(ori_ori_n334_), .Y(ori_ori_n335_));
  AOI210     o319(.A0(ori_ori_n335_), .A1(ori_ori_n330_), .B0(ori_ori_n25_), .Y(ori_ori_n336_));
  AOI210     o320(.A0(ori_ori_n110_), .A1(ori_ori_n108_), .B0(ori_ori_n42_), .Y(ori_ori_n337_));
  NOi21      o321(.An(ori_ori_n337_), .B(ori_ori_n171_), .Y(ori_ori_n338_));
  NA2        o322(.A(ori_ori_n338_), .B(ori_ori_n139_), .Y(ori_ori_n339_));
  INV        o323(.A(ori_ori_n339_), .Y(ori_ori_n340_));
  OAI210     o324(.A0(ori_ori_n340_), .A1(ori_ori_n336_), .B0(x6), .Y(ori_ori_n341_));
  NA3        o325(.A(ori_ori_n55_), .B(ori_ori_n38_), .C(ori_ori_n31_), .Y(ori_ori_n342_));
  AOI210     o326(.A0(ori_ori_n342_), .A1(x0), .B0(ori_ori_n32_), .Y(ori_ori_n343_));
  AOI210     o327(.A0(ori_ori_n117_), .A1(x2), .B0(x1), .Y(ori_ori_n344_));
  INV        o328(.A(ori_ori_n344_), .Y(ori_ori_n345_));
  NAi31      o329(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n346_));
  OAI210     o330(.A0(ori_ori_n346_), .A1(x4), .B0(ori_ori_n153_), .Y(ori_ori_n347_));
  NA3        o331(.A(ori_ori_n347_), .B(ori_ori_n137_), .C(x9), .Y(ori_ori_n348_));
  NO3        o332(.A(x9), .B(ori_ori_n142_), .C(x0), .Y(ori_ori_n349_));
  AOI220     o333(.A0(ori_ori_n349_), .A1(ori_ori_n229_), .B0(ori_ori_n311_), .B1(ori_ori_n142_), .Y(ori_ori_n350_));
  NA4        o334(.A(ori_ori_n350_), .B(x1), .C(ori_ori_n348_), .D(ori_ori_n50_), .Y(ori_ori_n351_));
  OAI210     o335(.A0(ori_ori_n345_), .A1(ori_ori_n343_), .B0(ori_ori_n351_), .Y(ori_ori_n352_));
  AOI210     o336(.A0(ori_ori_n38_), .A1(x9), .B0(ori_ori_n124_), .Y(ori_ori_n353_));
  NO3        o337(.A(ori_ori_n353_), .B(ori_ori_n114_), .C(ori_ori_n43_), .Y(ori_ori_n354_));
  NOi31      o338(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n355_));
  AOI220     o339(.A0(ori_ori_n355_), .A1(x4), .B0(ori_ori_n115_), .B1(x3), .Y(ori_ori_n356_));
  AOI210     o340(.A0(x1), .A1(ori_ori_n60_), .B0(ori_ori_n113_), .Y(ori_ori_n357_));
  OAI210     o341(.A0(ori_ori_n357_), .A1(x3), .B0(ori_ori_n356_), .Y(ori_ori_n358_));
  NO3        o342(.A(ori_ori_n358_), .B(ori_ori_n354_), .C(x2), .Y(ori_ori_n359_));
  OAI210     o343(.A0(ori_ori_n265_), .A1(ori_ori_n43_), .B0(ori_ori_n302_), .Y(ori_ori_n360_));
  AOI210     o344(.A0(x9), .A1(ori_ori_n48_), .B0(ori_ori_n332_), .Y(ori_ori_n361_));
  AOI220     o345(.A0(ori_ori_n361_), .A1(ori_ori_n87_), .B0(ori_ori_n360_), .B1(ori_ori_n142_), .Y(ori_ori_n362_));
  NO2        o346(.A(ori_ori_n362_), .B(ori_ori_n54_), .Y(ori_ori_n363_));
  NO2        o347(.A(ori_ori_n363_), .B(ori_ori_n359_), .Y(ori_ori_n364_));
  AOI210     o348(.A0(ori_ori_n364_), .A1(ori_ori_n352_), .B0(ori_ori_n25_), .Y(ori_ori_n365_));
  NA4        o349(.A(ori_ori_n31_), .B(ori_ori_n87_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n366_));
  NO3        o350(.A(ori_ori_n62_), .B(x4), .C(x1), .Y(ori_ori_n367_));
  NA2        o351(.A(ori_ori_n367_), .B(ori_ori_n337_), .Y(ori_ori_n368_));
  NO2        o352(.A(ori_ori_n368_), .B(ori_ori_n98_), .Y(ori_ori_n369_));
  NO3        o353(.A(ori_ori_n393_), .B(ori_ori_n165_), .C(ori_ori_n40_), .Y(ori_ori_n370_));
  OAI210     o354(.A0(ori_ori_n370_), .A1(ori_ori_n369_), .B0(x7), .Y(ori_ori_n371_));
  NA2        o355(.A(ori_ori_n371_), .B(ori_ori_n366_), .Y(ori_ori_n372_));
  OAI210     o356(.A0(ori_ori_n372_), .A1(ori_ori_n365_), .B0(ori_ori_n36_), .Y(ori_ori_n373_));
  NO2        o357(.A(ori_ori_n349_), .B(ori_ori_n191_), .Y(ori_ori_n374_));
  NO4        o358(.A(ori_ori_n374_), .B(ori_ori_n75_), .C(x4), .D(ori_ori_n54_), .Y(ori_ori_n375_));
  NA2        o359(.A(ori_ori_n236_), .B(ori_ori_n21_), .Y(ori_ori_n376_));
  NO2        o360(.A(ori_ori_n150_), .B(ori_ori_n125_), .Y(ori_ori_n377_));
  NA2        o361(.A(ori_ori_n377_), .B(ori_ori_n376_), .Y(ori_ori_n378_));
  AOI210     o362(.A0(ori_ori_n378_), .A1(ori_ori_n156_), .B0(ori_ori_n28_), .Y(ori_ori_n379_));
  NA2        o363(.A(ori_ori_n140_), .B(ori_ori_n187_), .Y(ori_ori_n380_));
  NA3        o364(.A(ori_ori_n380_), .B(ori_ori_n346_), .C(ori_ori_n85_), .Y(ori_ori_n381_));
  NA2        o365(.A(ori_ori_n381_), .B(ori_ori_n166_), .Y(ori_ori_n382_));
  OAI220     o366(.A0(ori_ori_n244_), .A1(ori_ori_n66_), .B0(ori_ori_n150_), .B1(ori_ori_n43_), .Y(ori_ori_n383_));
  NA2        o367(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n384_));
  NO2        o368(.A(ori_ori_n143_), .B(ori_ori_n384_), .Y(ori_ori_n385_));
  AOI220     o369(.A0(ori_ori_n385_), .A1(x0), .B0(ori_ori_n383_), .B1(ori_ori_n125_), .Y(ori_ori_n386_));
  AOI210     o370(.A0(ori_ori_n386_), .A1(ori_ori_n382_), .B0(ori_ori_n217_), .Y(ori_ori_n387_));
  NO3        o371(.A(ori_ori_n387_), .B(ori_ori_n379_), .C(ori_ori_n375_), .Y(ori_ori_n388_));
  NA3        o372(.A(ori_ori_n388_), .B(ori_ori_n373_), .C(ori_ori_n341_), .Y(ori_ori_n389_));
  AOI210     o373(.A0(ori_ori_n327_), .A1(ori_ori_n25_), .B0(ori_ori_n389_), .Y(ori05));
  INV        o374(.A(x2), .Y(ori_ori_n393_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  INV        m012(.A(mai_mai_n24_), .Y(mai_mai_n29_));
  NO2        m013(.A(x4), .B(x3), .Y(mai_mai_n30_));
  INV        m014(.A(mai_mai_n30_), .Y(mai_mai_n31_));
  OA210      m015(.A0(mai_mai_n31_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n32_));
  NOi31      m016(.An(mai_mai_n23_), .B(mai_mai_n32_), .C(mai_mai_n29_), .Y(mai00));
  NO2        m017(.A(x1), .B(x0), .Y(mai_mai_n34_));
  INV        m018(.A(x6), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n35_), .B(mai_mai_n25_), .Y(mai_mai_n36_));
  NA2        m020(.A(x4), .B(x3), .Y(mai_mai_n37_));
  NO2        m021(.A(mai_mai_n23_), .B(mai_mai_n37_), .Y(mai_mai_n38_));
  NO2        m022(.A(x2), .B(x0), .Y(mai_mai_n39_));
  INV        m023(.A(x3), .Y(mai_mai_n40_));
  NO2        m024(.A(mai_mai_n40_), .B(mai_mai_n18_), .Y(mai_mai_n41_));
  INV        m025(.A(mai_mai_n41_), .Y(mai_mai_n42_));
  NO2        m026(.A(mai_mai_n36_), .B(x4), .Y(mai_mai_n43_));
  OAI210     m027(.A0(mai_mai_n43_), .A1(mai_mai_n42_), .B0(mai_mai_n39_), .Y(mai_mai_n44_));
  INV        m028(.A(x4), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n45_), .B(mai_mai_n17_), .Y(mai_mai_n46_));
  NA2        m030(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n47_));
  OAI210     m031(.A0(mai_mai_n47_), .A1(mai_mai_n20_), .B0(mai_mai_n44_), .Y(mai_mai_n48_));
  AOI210     m032(.A0(mai_mai_n22_), .A1(mai_mai_n19_), .B0(mai_mai_n34_), .Y(mai_mai_n49_));
  INV        m033(.A(x2), .Y(mai_mai_n50_));
  NO2        m034(.A(mai_mai_n50_), .B(mai_mai_n17_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n40_), .B(mai_mai_n18_), .Y(mai_mai_n52_));
  NA2        m036(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  OAI210     m037(.A0(mai_mai_n49_), .A1(mai_mai_n31_), .B0(mai_mai_n53_), .Y(mai_mai_n54_));
  NO3        m038(.A(mai_mai_n54_), .B(mai_mai_n48_), .C(mai_mai_n38_), .Y(mai01));
  NA2        m039(.A(x8), .B(x7), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n40_), .B(x1), .Y(mai_mai_n57_));
  INV        m041(.A(x9), .Y(mai_mai_n58_));
  NO2        m042(.A(mai_mai_n58_), .B(mai_mai_n35_), .Y(mai_mai_n59_));
  INV        m043(.A(mai_mai_n59_), .Y(mai_mai_n60_));
  NO3        m044(.A(mai_mai_n60_), .B(mai_mai_n57_), .C(mai_mai_n56_), .Y(mai_mai_n61_));
  NO2        m045(.A(x7), .B(x6), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n63_));
  NO2        m047(.A(x8), .B(x2), .Y(mai_mai_n64_));
  AN2        m048(.A(mai_mai_n63_), .B(mai_mai_n62_), .Y(mai_mai_n65_));
  OAI210     m049(.A0(mai_mai_n41_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n66_));
  OAI210     m050(.A0(mai_mai_n52_), .A1(mai_mai_n20_), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  NAi31      m051(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n68_));
  NO2        m052(.A(mai_mai_n67_), .B(mai_mai_n65_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n69_), .A1(mai_mai_n61_), .B0(x4), .Y(mai_mai_n70_));
  NA2        m054(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n71_));
  OAI210     m055(.A0(mai_mai_n71_), .A1(mai_mai_n52_), .B0(x0), .Y(mai_mai_n72_));
  NA2        m056(.A(x5), .B(x3), .Y(mai_mai_n73_));
  NO2        m057(.A(x8), .B(x6), .Y(mai_mai_n74_));
  NO4        m058(.A(mai_mai_n74_), .B(mai_mai_n73_), .C(mai_mai_n62_), .D(mai_mai_n50_), .Y(mai_mai_n75_));
  NAi21      m059(.An(x4), .B(x3), .Y(mai_mai_n76_));
  INV        m060(.A(mai_mai_n76_), .Y(mai_mai_n77_));
  NO2        m061(.A(mai_mai_n77_), .B(mai_mai_n22_), .Y(mai_mai_n78_));
  NO2        m062(.A(x4), .B(x2), .Y(mai_mai_n79_));
  NO2        m063(.A(mai_mai_n79_), .B(x3), .Y(mai_mai_n80_));
  NO3        m064(.A(mai_mai_n80_), .B(mai_mai_n78_), .C(mai_mai_n18_), .Y(mai_mai_n81_));
  NO3        m065(.A(mai_mai_n81_), .B(mai_mai_n75_), .C(mai_mai_n72_), .Y(mai_mai_n82_));
  NO3        m066(.A(x6), .B(mai_mai_n40_), .C(x1), .Y(mai_mai_n83_));
  NA2        m067(.A(mai_mai_n58_), .B(mai_mai_n45_), .Y(mai_mai_n84_));
  INV        m068(.A(mai_mai_n84_), .Y(mai_mai_n85_));
  OAI210     m069(.A0(mai_mai_n83_), .A1(mai_mai_n63_), .B0(mai_mai_n85_), .Y(mai_mai_n86_));
  NA2        m070(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n87_));
  NO2        m071(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n88_));
  INV        m072(.A(x8), .Y(mai_mai_n89_));
  NA2        m073(.A(x2), .B(x1), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n91_));
  NO2        m075(.A(mai_mai_n91_), .B(mai_mai_n88_), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n92_), .B(mai_mai_n26_), .Y(mai_mai_n93_));
  AOI210     m077(.A0(mai_mai_n52_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n94_));
  OAI210     m078(.A0(mai_mai_n42_), .A1(mai_mai_n36_), .B0(mai_mai_n45_), .Y(mai_mai_n95_));
  NO3        m079(.A(mai_mai_n95_), .B(mai_mai_n94_), .C(mai_mai_n93_), .Y(mai_mai_n96_));
  NA2        m080(.A(x4), .B(mai_mai_n40_), .Y(mai_mai_n97_));
  NO2        m081(.A(mai_mai_n45_), .B(mai_mai_n50_), .Y(mai_mai_n98_));
  NO2        m082(.A(mai_mai_n97_), .B(x1), .Y(mai_mai_n99_));
  NO2        m083(.A(x3), .B(x2), .Y(mai_mai_n100_));
  NA3        m084(.A(mai_mai_n100_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n101_));
  AOI210     m085(.A0(x8), .A1(x6), .B0(mai_mai_n101_), .Y(mai_mai_n102_));
  NA2        m086(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n103_));
  OAI210     m087(.A0(mai_mai_n103_), .A1(mai_mai_n37_), .B0(mai_mai_n17_), .Y(mai_mai_n104_));
  NO4        m088(.A(mai_mai_n104_), .B(mai_mai_n102_), .C(mai_mai_n99_), .D(mai_mai_n96_), .Y(mai_mai_n105_));
  AO220      m089(.A0(mai_mai_n105_), .A1(mai_mai_n86_), .B0(mai_mai_n82_), .B1(mai_mai_n70_), .Y(mai02));
  NO2        m090(.A(x3), .B(mai_mai_n50_), .Y(mai_mai_n107_));
  NO2        m091(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n108_));
  NA2        m092(.A(mai_mai_n40_), .B(x0), .Y(mai_mai_n109_));
  OAI210     m093(.A0(mai_mai_n84_), .A1(x2), .B0(mai_mai_n109_), .Y(mai_mai_n110_));
  AOI220     m094(.A0(mai_mai_n110_), .A1(mai_mai_n108_), .B0(mai_mai_n107_), .B1(x4), .Y(mai_mai_n111_));
  NO3        m095(.A(mai_mai_n111_), .B(x7), .C(x5), .Y(mai_mai_n112_));
  NA2        m096(.A(x9), .B(x2), .Y(mai_mai_n113_));
  OR2        m097(.A(x8), .B(x0), .Y(mai_mai_n114_));
  INV        m098(.A(mai_mai_n114_), .Y(mai_mai_n115_));
  NAi21      m099(.An(x2), .B(x8), .Y(mai_mai_n116_));
  INV        m100(.A(mai_mai_n116_), .Y(mai_mai_n117_));
  OAI220     m101(.A0(mai_mai_n117_), .A1(mai_mai_n115_), .B0(mai_mai_n113_), .B1(x7), .Y(mai_mai_n118_));
  NO2        m102(.A(x4), .B(x1), .Y(mai_mai_n119_));
  NA2        m103(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n120_));
  NO3        m104(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n121_));
  NOi21      m105(.An(x0), .B(x4), .Y(mai_mai_n122_));
  NO2        m106(.A(mai_mai_n120_), .B(mai_mai_n73_), .Y(mai_mai_n123_));
  NO2        m107(.A(x5), .B(mai_mai_n45_), .Y(mai_mai_n124_));
  NA2        m108(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n125_));
  AOI210     m109(.A0(mai_mai_n125_), .A1(mai_mai_n103_), .B0(mai_mai_n109_), .Y(mai_mai_n126_));
  OAI210     m110(.A0(mai_mai_n126_), .A1(mai_mai_n34_), .B0(mai_mai_n124_), .Y(mai_mai_n127_));
  NAi21      m111(.An(x0), .B(x4), .Y(mai_mai_n128_));
  NO2        m112(.A(mai_mai_n128_), .B(x1), .Y(mai_mai_n129_));
  NO2        m113(.A(x7), .B(x0), .Y(mai_mai_n130_));
  NO2        m114(.A(mai_mai_n79_), .B(mai_mai_n98_), .Y(mai_mai_n131_));
  NO2        m115(.A(mai_mai_n131_), .B(x3), .Y(mai_mai_n132_));
  OAI210     m116(.A0(mai_mai_n130_), .A1(mai_mai_n129_), .B0(mai_mai_n132_), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n21_), .B(mai_mai_n40_), .Y(mai_mai_n134_));
  NA2        m118(.A(x5), .B(x0), .Y(mai_mai_n135_));
  NO2        m119(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n136_));
  NA3        m120(.A(mai_mai_n136_), .B(mai_mai_n135_), .C(mai_mai_n134_), .Y(mai_mai_n137_));
  NA4        m121(.A(mai_mai_n137_), .B(mai_mai_n133_), .C(mai_mai_n127_), .D(mai_mai_n35_), .Y(mai_mai_n138_));
  NO3        m122(.A(mai_mai_n138_), .B(mai_mai_n123_), .C(mai_mai_n112_), .Y(mai_mai_n139_));
  NO3        m123(.A(mai_mai_n73_), .B(mai_mai_n71_), .C(mai_mai_n24_), .Y(mai_mai_n140_));
  NO2        m124(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n141_));
  AOI220     m125(.A0(x0), .A1(mai_mai_n141_), .B0(mai_mai_n63_), .B1(mai_mai_n17_), .Y(mai_mai_n142_));
  NO3        m126(.A(mai_mai_n142_), .B(mai_mai_n56_), .C(mai_mai_n58_), .Y(mai_mai_n143_));
  NO2        m127(.A(mai_mai_n97_), .B(x5), .Y(mai_mai_n144_));
  NO2        m128(.A(x9), .B(x7), .Y(mai_mai_n145_));
  NOi21      m129(.An(x8), .B(x0), .Y(mai_mai_n146_));
  NO2        m130(.A(mai_mai_n40_), .B(x2), .Y(mai_mai_n147_));
  INV        m131(.A(x7), .Y(mai_mai_n148_));
  NA2        m132(.A(mai_mai_n148_), .B(mai_mai_n18_), .Y(mai_mai_n149_));
  NA2        m133(.A(mai_mai_n149_), .B(mai_mai_n147_), .Y(mai_mai_n150_));
  NO2        m134(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n151_), .B(mai_mai_n122_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n152_), .B(mai_mai_n150_), .Y(mai_mai_n153_));
  AOI210     m137(.A0(mai_mai_n146_), .A1(mai_mai_n144_), .B0(mai_mai_n153_), .Y(mai_mai_n154_));
  INV        m138(.A(mai_mai_n154_), .Y(mai_mai_n155_));
  NA2        m139(.A(x5), .B(x1), .Y(mai_mai_n156_));
  INV        m140(.A(mai_mai_n156_), .Y(mai_mai_n157_));
  AOI210     m141(.A0(mai_mai_n157_), .A1(mai_mai_n122_), .B0(mai_mai_n35_), .Y(mai_mai_n158_));
  NO2        m142(.A(mai_mai_n58_), .B(mai_mai_n89_), .Y(mai_mai_n159_));
  NO3        m143(.A(x2), .B(mai_mai_n159_), .C(mai_mai_n45_), .Y(mai_mai_n160_));
  NA2        m144(.A(mai_mai_n160_), .B(mai_mai_n63_), .Y(mai_mai_n161_));
  NA2        m145(.A(mai_mai_n161_), .B(mai_mai_n158_), .Y(mai_mai_n162_));
  NO4        m146(.A(mai_mai_n162_), .B(mai_mai_n155_), .C(mai_mai_n143_), .D(mai_mai_n140_), .Y(mai_mai_n163_));
  NO2        m147(.A(mai_mai_n163_), .B(mai_mai_n139_), .Y(mai_mai_n164_));
  NO2        m148(.A(mai_mai_n135_), .B(mai_mai_n131_), .Y(mai_mai_n165_));
  NA2        m149(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n166_));
  NA2        m150(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n167_));
  NA3        m151(.A(mai_mai_n167_), .B(mai_mai_n166_), .C(mai_mai_n24_), .Y(mai_mai_n168_));
  AN2        m152(.A(mai_mai_n168_), .B(mai_mai_n136_), .Y(mai_mai_n169_));
  NA2        m153(.A(x8), .B(x0), .Y(mai_mai_n170_));
  NO2        m154(.A(mai_mai_n148_), .B(mai_mai_n25_), .Y(mai_mai_n171_));
  NA2        m155(.A(x2), .B(x0), .Y(mai_mai_n172_));
  NA2        m156(.A(x4), .B(x1), .Y(mai_mai_n173_));
  NAi21      m157(.An(mai_mai_n119_), .B(mai_mai_n173_), .Y(mai_mai_n174_));
  NOi31      m158(.An(mai_mai_n174_), .B(mai_mai_n151_), .C(mai_mai_n172_), .Y(mai_mai_n175_));
  NO3        m159(.A(mai_mai_n175_), .B(mai_mai_n169_), .C(mai_mai_n165_), .Y(mai_mai_n176_));
  NO2        m160(.A(mai_mai_n176_), .B(mai_mai_n40_), .Y(mai_mai_n177_));
  NO2        m161(.A(mai_mai_n168_), .B(mai_mai_n71_), .Y(mai_mai_n178_));
  INV        m162(.A(mai_mai_n124_), .Y(mai_mai_n179_));
  NO2        m163(.A(mai_mai_n103_), .B(mai_mai_n17_), .Y(mai_mai_n180_));
  NA3        m164(.A(mai_mai_n174_), .B(mai_mai_n179_), .C(mai_mai_n39_), .Y(mai_mai_n181_));
  OAI210     m165(.A0(mai_mai_n167_), .A1(mai_mai_n131_), .B0(mai_mai_n181_), .Y(mai_mai_n182_));
  NO2        m166(.A(mai_mai_n182_), .B(mai_mai_n178_), .Y(mai_mai_n183_));
  NO2        m167(.A(mai_mai_n183_), .B(x3), .Y(mai_mai_n184_));
  NO3        m168(.A(mai_mai_n184_), .B(mai_mai_n177_), .C(mai_mai_n164_), .Y(mai03));
  NO2        m169(.A(mai_mai_n45_), .B(x3), .Y(mai_mai_n186_));
  NO2        m170(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n187_));
  NA2        m171(.A(mai_mai_n59_), .B(mai_mai_n186_), .Y(mai_mai_n188_));
  NO2        m172(.A(mai_mai_n73_), .B(x6), .Y(mai_mai_n189_));
  NA2        m173(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n190_));
  NO2        m174(.A(mai_mai_n190_), .B(x4), .Y(mai_mai_n191_));
  NO2        m175(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n192_));
  AO220      m176(.A0(mai_mai_n192_), .A1(mai_mai_n191_), .B0(mai_mai_n189_), .B1(mai_mai_n51_), .Y(mai_mai_n193_));
  NA2        m177(.A(mai_mai_n193_), .B(mai_mai_n58_), .Y(mai_mai_n194_));
  NA2        m178(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n195_));
  NA2        m179(.A(x9), .B(mai_mai_n50_), .Y(mai_mai_n196_));
  NA2        m180(.A(mai_mai_n190_), .B(mai_mai_n76_), .Y(mai_mai_n197_));
  AOI210     m181(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n172_), .Y(mai_mai_n198_));
  NA2        m182(.A(mai_mai_n198_), .B(mai_mai_n197_), .Y(mai_mai_n199_));
  NO3        m183(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n200_));
  NO2        m184(.A(x5), .B(x1), .Y(mai_mai_n201_));
  AOI220     m185(.A0(mai_mai_n201_), .A1(mai_mai_n17_), .B0(mai_mai_n100_), .B1(x5), .Y(mai_mai_n202_));
  NO2        m186(.A(mai_mai_n195_), .B(mai_mai_n166_), .Y(mai_mai_n203_));
  INV        m187(.A(mai_mai_n203_), .Y(mai_mai_n204_));
  OAI210     m188(.A0(mai_mai_n202_), .A1(mai_mai_n60_), .B0(mai_mai_n204_), .Y(mai_mai_n205_));
  AOI220     m189(.A0(mai_mai_n205_), .A1(mai_mai_n45_), .B0(mai_mai_n200_), .B1(mai_mai_n124_), .Y(mai_mai_n206_));
  NA4        m190(.A(mai_mai_n206_), .B(mai_mai_n199_), .C(mai_mai_n194_), .D(mai_mai_n188_), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n208_));
  NA2        m192(.A(mai_mai_n208_), .B(mai_mai_n19_), .Y(mai_mai_n209_));
  NO2        m193(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n210_));
  NO2        m194(.A(mai_mai_n210_), .B(x6), .Y(mai_mai_n211_));
  NOi21      m195(.An(mai_mai_n79_), .B(mai_mai_n211_), .Y(mai_mai_n212_));
  NA2        m196(.A(mai_mai_n58_), .B(mai_mai_n89_), .Y(mai_mai_n213_));
  NA3        m197(.A(mai_mai_n213_), .B(mai_mai_n210_), .C(x6), .Y(mai_mai_n214_));
  AOI210     m198(.A0(mai_mai_n214_), .A1(mai_mai_n212_), .B0(mai_mai_n148_), .Y(mai_mai_n215_));
  AO210      m199(.A0(mai_mai_n215_), .A1(mai_mai_n209_), .B0(mai_mai_n171_), .Y(mai_mai_n216_));
  NA2        m200(.A(mai_mai_n40_), .B(mai_mai_n50_), .Y(mai_mai_n217_));
  OAI210     m201(.A0(mai_mai_n217_), .A1(mai_mai_n25_), .B0(mai_mai_n167_), .Y(mai_mai_n218_));
  NO3        m202(.A(mai_mai_n173_), .B(mai_mai_n58_), .C(x6), .Y(mai_mai_n219_));
  AOI220     m203(.A0(mai_mai_n219_), .A1(mai_mai_n218_), .B0(mai_mai_n136_), .B1(mai_mai_n88_), .Y(mai_mai_n220_));
  NA2        m204(.A(x6), .B(mai_mai_n45_), .Y(mai_mai_n221_));
  OAI210     m205(.A0(mai_mai_n115_), .A1(mai_mai_n74_), .B0(x4), .Y(mai_mai_n222_));
  AOI210     m206(.A0(mai_mai_n222_), .A1(mai_mai_n221_), .B0(mai_mai_n73_), .Y(mai_mai_n223_));
  NA2        m207(.A(mai_mai_n187_), .B(mai_mai_n129_), .Y(mai_mai_n224_));
  OAI210     m208(.A0(mai_mai_n89_), .A1(mai_mai_n35_), .B0(mai_mai_n63_), .Y(mai_mai_n225_));
  NA2        m209(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n226_));
  OAI210     m210(.A0(mai_mai_n226_), .A1(mai_mai_n223_), .B0(x2), .Y(mai_mai_n227_));
  NA3        m211(.A(mai_mai_n227_), .B(mai_mai_n220_), .C(mai_mai_n216_), .Y(mai_mai_n228_));
  AOI210     m212(.A0(mai_mai_n207_), .A1(x8), .B0(mai_mai_n228_), .Y(mai_mai_n229_));
  NO2        m213(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n230_));
  AOI210     m214(.A0(mai_mai_n211_), .A1(mai_mai_n151_), .B0(mai_mai_n230_), .Y(mai_mai_n231_));
  NO2        m215(.A(mai_mai_n231_), .B(x2), .Y(mai_mai_n232_));
  NO2        m216(.A(x4), .B(mai_mai_n50_), .Y(mai_mai_n233_));
  AOI220     m217(.A0(mai_mai_n191_), .A1(mai_mai_n180_), .B0(mai_mai_n233_), .B1(mai_mai_n63_), .Y(mai_mai_n234_));
  NA3        m218(.A(mai_mai_n25_), .B(x3), .C(x2), .Y(mai_mai_n235_));
  NO2        m219(.A(mai_mai_n235_), .B(mai_mai_n413_), .Y(mai_mai_n236_));
  NA2        m220(.A(mai_mai_n236_), .B(mai_mai_n119_), .Y(mai_mai_n237_));
  NA2        m221(.A(mai_mai_n195_), .B(x6), .Y(mai_mai_n238_));
  NO2        m222(.A(mai_mai_n195_), .B(x6), .Y(mai_mai_n239_));
  NAi21      m223(.An(mai_mai_n159_), .B(mai_mai_n239_), .Y(mai_mai_n240_));
  NA3        m224(.A(mai_mai_n240_), .B(mai_mai_n238_), .C(mai_mai_n141_), .Y(mai_mai_n241_));
  NA4        m225(.A(mai_mai_n241_), .B(mai_mai_n237_), .C(mai_mai_n234_), .D(mai_mai_n148_), .Y(mai_mai_n242_));
  NA2        m226(.A(mai_mai_n187_), .B(mai_mai_n210_), .Y(mai_mai_n243_));
  NO2        m227(.A(x9), .B(x6), .Y(mai_mai_n244_));
  NO2        m228(.A(mai_mai_n135_), .B(mai_mai_n18_), .Y(mai_mai_n245_));
  NAi21      m229(.An(mai_mai_n245_), .B(mai_mai_n235_), .Y(mai_mai_n246_));
  NAi21      m230(.An(x1), .B(x4), .Y(mai_mai_n247_));
  AOI210     m231(.A0(x3), .A1(x2), .B0(mai_mai_n45_), .Y(mai_mai_n248_));
  OAI210     m232(.A0(mai_mai_n135_), .A1(x3), .B0(mai_mai_n248_), .Y(mai_mai_n249_));
  AOI220     m233(.A0(mai_mai_n249_), .A1(mai_mai_n247_), .B0(mai_mai_n246_), .B1(mai_mai_n244_), .Y(mai_mai_n250_));
  NA2        m234(.A(mai_mai_n250_), .B(mai_mai_n243_), .Y(mai_mai_n251_));
  NA2        m235(.A(mai_mai_n58_), .B(x2), .Y(mai_mai_n252_));
  NO2        m236(.A(mai_mai_n252_), .B(mai_mai_n243_), .Y(mai_mai_n253_));
  NO3        m237(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n254_));
  NA2        m238(.A(x6), .B(x2), .Y(mai_mai_n255_));
  INV        m239(.A(mai_mai_n254_), .Y(mai_mai_n256_));
  OAI210     m240(.A0(mai_mai_n256_), .A1(mai_mai_n40_), .B0(mai_mai_n412_), .Y(mai_mai_n257_));
  OAI210     m241(.A0(mai_mai_n257_), .A1(mai_mai_n253_), .B0(mai_mai_n251_), .Y(mai_mai_n258_));
  NA2        m242(.A(x4), .B(x0), .Y(mai_mai_n259_));
  NA2        m243(.A(mai_mai_n189_), .B(mai_mai_n39_), .Y(mai_mai_n260_));
  AOI210     m244(.A0(mai_mai_n260_), .A1(mai_mai_n258_), .B0(x8), .Y(mai_mai_n261_));
  NA2        m245(.A(mai_mai_n201_), .B(x6), .Y(mai_mai_n262_));
  INV        m246(.A(mai_mai_n170_), .Y(mai_mai_n263_));
  OAI210     m247(.A0(mai_mai_n263_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n264_));
  AOI210     m248(.A0(mai_mai_n264_), .A1(mai_mai_n262_), .B0(mai_mai_n217_), .Y(mai_mai_n265_));
  NO4        m249(.A(mai_mai_n265_), .B(mai_mai_n261_), .C(mai_mai_n242_), .D(mai_mai_n232_), .Y(mai_mai_n266_));
  NO2        m250(.A(mai_mai_n159_), .B(x1), .Y(mai_mai_n267_));
  NO3        m251(.A(mai_mai_n267_), .B(x3), .C(mai_mai_n35_), .Y(mai_mai_n268_));
  OAI210     m252(.A0(mai_mai_n268_), .A1(mai_mai_n239_), .B0(x2), .Y(mai_mai_n269_));
  OAI210     m253(.A0(mai_mai_n263_), .A1(x6), .B0(mai_mai_n41_), .Y(mai_mai_n270_));
  AOI210     m254(.A0(mai_mai_n270_), .A1(mai_mai_n269_), .B0(mai_mai_n179_), .Y(mai_mai_n271_));
  NOi21      m255(.An(mai_mai_n255_), .B(mai_mai_n17_), .Y(mai_mai_n272_));
  NA3        m256(.A(mai_mai_n272_), .B(mai_mai_n201_), .C(mai_mai_n37_), .Y(mai_mai_n273_));
  AOI210     m257(.A0(mai_mai_n35_), .A1(mai_mai_n50_), .B0(x0), .Y(mai_mai_n274_));
  NA3        m258(.A(mai_mai_n274_), .B(mai_mai_n157_), .C(mai_mai_n31_), .Y(mai_mai_n275_));
  NA2        m259(.A(x3), .B(x2), .Y(mai_mai_n276_));
  AOI220     m260(.A0(mai_mai_n276_), .A1(mai_mai_n217_), .B0(mai_mai_n275_), .B1(mai_mai_n273_), .Y(mai_mai_n277_));
  NAi21      m261(.An(x4), .B(x0), .Y(mai_mai_n278_));
  NO3        m262(.A(mai_mai_n278_), .B(mai_mai_n41_), .C(x2), .Y(mai_mai_n279_));
  OAI210     m263(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n279_), .Y(mai_mai_n280_));
  NO2        m264(.A(x9), .B(x8), .Y(mai_mai_n281_));
  NA3        m265(.A(mai_mai_n281_), .B(mai_mai_n35_), .C(mai_mai_n50_), .Y(mai_mai_n282_));
  OAI210     m266(.A0(mai_mai_n274_), .A1(mai_mai_n272_), .B0(mai_mai_n282_), .Y(mai_mai_n283_));
  AOI220     m267(.A0(mai_mai_n283_), .A1(mai_mai_n77_), .B0(mai_mai_n18_), .B1(mai_mai_n30_), .Y(mai_mai_n284_));
  AOI210     m268(.A0(mai_mai_n284_), .A1(mai_mai_n280_), .B0(mai_mai_n25_), .Y(mai_mai_n285_));
  NA3        m269(.A(mai_mai_n35_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n286_));
  OAI210     m270(.A0(mai_mai_n274_), .A1(mai_mai_n272_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  INV        m271(.A(mai_mai_n203_), .Y(mai_mai_n288_));
  NA2        m272(.A(mai_mai_n35_), .B(mai_mai_n40_), .Y(mai_mai_n289_));
  OR2        m273(.A(mai_mai_n289_), .B(mai_mai_n259_), .Y(mai_mai_n290_));
  OAI220     m274(.A0(mai_mai_n290_), .A1(mai_mai_n156_), .B0(mai_mai_n221_), .B1(mai_mai_n288_), .Y(mai_mai_n291_));
  AO210      m275(.A0(mai_mai_n287_), .A1(mai_mai_n144_), .B0(mai_mai_n291_), .Y(mai_mai_n292_));
  NO4        m276(.A(mai_mai_n292_), .B(mai_mai_n285_), .C(mai_mai_n277_), .D(mai_mai_n271_), .Y(mai_mai_n293_));
  OAI210     m277(.A0(mai_mai_n266_), .A1(mai_mai_n229_), .B0(mai_mai_n293_), .Y(mai04));
  NA2        m278(.A(mai_mai_n254_), .B(mai_mai_n80_), .Y(mai_mai_n295_));
  INV        m279(.A(mai_mai_n278_), .Y(mai_mai_n296_));
  NO2        m280(.A(mai_mai_n276_), .B(mai_mai_n192_), .Y(mai_mai_n297_));
  NA2        m281(.A(mai_mai_n297_), .B(x6), .Y(mai_mai_n298_));
  NO2        m282(.A(mai_mai_n196_), .B(mai_mai_n109_), .Y(mai_mai_n299_));
  NO3        m283(.A(mai_mai_n413_), .B(mai_mai_n116_), .C(mai_mai_n18_), .Y(mai_mai_n300_));
  NO2        m284(.A(mai_mai_n300_), .B(mai_mai_n299_), .Y(mai_mai_n301_));
  OAI210     m285(.A0(mai_mai_n114_), .A1(mai_mai_n103_), .B0(mai_mai_n170_), .Y(mai_mai_n302_));
  NA3        m286(.A(mai_mai_n302_), .B(x6), .C(x3), .Y(mai_mai_n303_));
  OAI210     m287(.A0(mai_mai_n252_), .A1(mai_mai_n286_), .B0(mai_mai_n289_), .Y(mai_mai_n304_));
  INV        m288(.A(mai_mai_n304_), .Y(mai_mai_n305_));
  NA4        m289(.A(mai_mai_n414_), .B(mai_mai_n305_), .C(mai_mai_n303_), .D(mai_mai_n301_), .Y(mai_mai_n306_));
  OAI210     m290(.A0(mai_mai_n108_), .A1(x3), .B0(mai_mai_n279_), .Y(mai_mai_n307_));
  NA3        m291(.A(mai_mai_n213_), .B(mai_mai_n200_), .C(mai_mai_n79_), .Y(mai_mai_n308_));
  NA3        m292(.A(mai_mai_n308_), .B(mai_mai_n307_), .C(mai_mai_n148_), .Y(mai_mai_n309_));
  AOI210     m293(.A0(mai_mai_n306_), .A1(x4), .B0(mai_mai_n309_), .Y(mai_mai_n310_));
  NA3        m294(.A(mai_mai_n296_), .B(mai_mai_n196_), .C(mai_mai_n89_), .Y(mai_mai_n311_));
  NOi21      m295(.An(x4), .B(x0), .Y(mai_mai_n312_));
  XO2        m296(.A(x4), .B(x0), .Y(mai_mai_n313_));
  OAI210     m297(.A0(mai_mai_n313_), .A1(mai_mai_n113_), .B0(mai_mai_n247_), .Y(mai_mai_n314_));
  AOI220     m298(.A0(mai_mai_n314_), .A1(x8), .B0(mai_mai_n312_), .B1(mai_mai_n90_), .Y(mai_mai_n315_));
  AOI210     m299(.A0(mai_mai_n315_), .A1(mai_mai_n311_), .B0(x3), .Y(mai_mai_n316_));
  INV        m300(.A(mai_mai_n90_), .Y(mai_mai_n317_));
  NO2        m301(.A(mai_mai_n89_), .B(x4), .Y(mai_mai_n318_));
  AOI220     m302(.A0(mai_mai_n318_), .A1(mai_mai_n41_), .B0(mai_mai_n122_), .B1(mai_mai_n317_), .Y(mai_mai_n319_));
  NO3        m303(.A(mai_mai_n313_), .B(mai_mai_n159_), .C(x2), .Y(mai_mai_n320_));
  NO3        m304(.A(mai_mai_n213_), .B(mai_mai_n28_), .C(mai_mai_n24_), .Y(mai_mai_n321_));
  NO2        m305(.A(mai_mai_n321_), .B(mai_mai_n320_), .Y(mai_mai_n322_));
  NA4        m306(.A(mai_mai_n322_), .B(mai_mai_n319_), .C(mai_mai_n209_), .D(x6), .Y(mai_mai_n323_));
  OAI220     m307(.A0(mai_mai_n278_), .A1(mai_mai_n87_), .B0(mai_mai_n172_), .B1(mai_mai_n89_), .Y(mai_mai_n324_));
  NO2        m308(.A(mai_mai_n40_), .B(x0), .Y(mai_mai_n325_));
  OR2        m309(.A(mai_mai_n318_), .B(mai_mai_n325_), .Y(mai_mai_n326_));
  NO2        m310(.A(mai_mai_n146_), .B(mai_mai_n103_), .Y(mai_mai_n327_));
  AOI220     m311(.A0(mai_mai_n327_), .A1(mai_mai_n326_), .B0(mai_mai_n324_), .B1(mai_mai_n57_), .Y(mai_mai_n328_));
  NO2        m312(.A(mai_mai_n146_), .B(mai_mai_n76_), .Y(mai_mai_n329_));
  NO2        m313(.A(mai_mai_n34_), .B(x2), .Y(mai_mai_n330_));
  NOi21      m314(.An(mai_mai_n119_), .B(mai_mai_n27_), .Y(mai_mai_n331_));
  AOI210     m315(.A0(mai_mai_n330_), .A1(mai_mai_n329_), .B0(mai_mai_n331_), .Y(mai_mai_n332_));
  OAI210     m316(.A0(mai_mai_n328_), .A1(mai_mai_n58_), .B0(mai_mai_n332_), .Y(mai_mai_n333_));
  OAI220     m317(.A0(mai_mai_n333_), .A1(x6), .B0(mai_mai_n323_), .B1(mai_mai_n316_), .Y(mai_mai_n334_));
  INV        m318(.A(mai_mai_n290_), .Y(mai_mai_n335_));
  AOI210     m319(.A0(mai_mai_n335_), .A1(mai_mai_n18_), .B0(mai_mai_n148_), .Y(mai_mai_n336_));
  AO220      m320(.A0(mai_mai_n336_), .A1(mai_mai_n334_), .B0(mai_mai_n310_), .B1(mai_mai_n298_), .Y(mai_mai_n337_));
  NA2        m321(.A(mai_mai_n330_), .B(x6), .Y(mai_mai_n338_));
  AOI210     m322(.A0(x6), .A1(x1), .B0(mai_mai_n147_), .Y(mai_mai_n339_));
  NA2        m323(.A(mai_mai_n318_), .B(x0), .Y(mai_mai_n340_));
  NA2        m324(.A(mai_mai_n79_), .B(x6), .Y(mai_mai_n341_));
  OAI210     m325(.A0(mai_mai_n340_), .A1(mai_mai_n339_), .B0(mai_mai_n341_), .Y(mai_mai_n342_));
  NA2        m326(.A(mai_mai_n342_), .B(mai_mai_n338_), .Y(mai_mai_n343_));
  NA3        m327(.A(mai_mai_n343_), .B(mai_mai_n337_), .C(mai_mai_n295_), .Y(mai_mai_n344_));
  NA3        m328(.A(mai_mai_n108_), .B(mai_mai_n186_), .C(mai_mai_n148_), .Y(mai_mai_n345_));
  OAI210     m329(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n217_), .Y(mai_mai_n346_));
  AO220      m330(.A0(mai_mai_n346_), .A1(mai_mai_n145_), .B0(mai_mai_n107_), .B1(x4), .Y(mai_mai_n347_));
  NA3        m331(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n348_));
  NA2        m332(.A(mai_mai_n208_), .B(x0), .Y(mai_mai_n349_));
  OAI220     m333(.A0(mai_mai_n349_), .A1(mai_mai_n196_), .B0(mai_mai_n348_), .B1(mai_mai_n317_), .Y(mai_mai_n350_));
  AOI210     m334(.A0(mai_mai_n347_), .A1(mai_mai_n115_), .B0(mai_mai_n350_), .Y(mai_mai_n351_));
  AOI210     m335(.A0(mai_mai_n351_), .A1(mai_mai_n345_), .B0(mai_mai_n25_), .Y(mai_mai_n352_));
  NA3        m336(.A(mai_mai_n117_), .B(mai_mai_n208_), .C(x0), .Y(mai_mai_n353_));
  OAI210     m337(.A0(mai_mai_n186_), .A1(mai_mai_n64_), .B0(mai_mai_n192_), .Y(mai_mai_n354_));
  NO2        m338(.A(mai_mai_n354_), .B(mai_mai_n25_), .Y(mai_mai_n355_));
  NA2        m339(.A(mai_mai_n355_), .B(mai_mai_n145_), .Y(mai_mai_n356_));
  NAi31      m340(.An(mai_mai_n47_), .B(mai_mai_n267_), .C(mai_mai_n171_), .Y(mai_mai_n357_));
  NA3        m341(.A(mai_mai_n357_), .B(mai_mai_n356_), .C(mai_mai_n353_), .Y(mai_mai_n358_));
  OAI210     m342(.A0(mai_mai_n358_), .A1(mai_mai_n352_), .B0(x6), .Y(mai_mai_n359_));
  OAI210     m343(.A0(mai_mai_n159_), .A1(mai_mai_n45_), .B0(mai_mai_n130_), .Y(mai_mai_n360_));
  AOI210     m344(.A0(mai_mai_n37_), .A1(mai_mai_n31_), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  NO2        m345(.A(mai_mai_n148_), .B(x0), .Y(mai_mai_n362_));
  AOI220     m346(.A0(mai_mai_n362_), .A1(mai_mai_n208_), .B0(mai_mai_n186_), .B1(mai_mai_n148_), .Y(mai_mai_n363_));
  INV        m347(.A(x1), .Y(mai_mai_n364_));
  OAI210     m348(.A0(mai_mai_n363_), .A1(x8), .B0(mai_mai_n364_), .Y(mai_mai_n365_));
  NO4        m349(.A(x8), .B(mai_mai_n278_), .C(x9), .D(x2), .Y(mai_mai_n366_));
  NOi21      m350(.An(mai_mai_n121_), .B(mai_mai_n172_), .Y(mai_mai_n367_));
  NO3        m351(.A(mai_mai_n367_), .B(mai_mai_n366_), .C(mai_mai_n18_), .Y(mai_mai_n368_));
  NA2        m352(.A(mai_mai_n329_), .B(mai_mai_n148_), .Y(mai_mai_n369_));
  NA3        m353(.A(mai_mai_n369_), .B(mai_mai_n368_), .C(mai_mai_n47_), .Y(mai_mai_n370_));
  OAI210     m354(.A0(mai_mai_n365_), .A1(mai_mai_n361_), .B0(mai_mai_n370_), .Y(mai_mai_n371_));
  NOi31      m355(.An(mai_mai_n362_), .B(mai_mai_n31_), .C(x8), .Y(mai_mai_n372_));
  INV        m356(.A(mai_mai_n128_), .Y(mai_mai_n373_));
  NO3        m357(.A(mai_mai_n373_), .B(mai_mai_n121_), .C(mai_mai_n40_), .Y(mai_mai_n374_));
  NOi31      m358(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n375_));
  AOI220     m359(.A0(mai_mai_n375_), .A1(mai_mai_n312_), .B0(mai_mai_n122_), .B1(x3), .Y(mai_mai_n376_));
  AOI210     m360(.A0(mai_mai_n247_), .A1(mai_mai_n56_), .B0(x0), .Y(mai_mai_n377_));
  OAI210     m361(.A0(mai_mai_n377_), .A1(x3), .B0(mai_mai_n376_), .Y(mai_mai_n378_));
  NO3        m362(.A(mai_mai_n378_), .B(mai_mai_n374_), .C(x2), .Y(mai_mai_n379_));
  OAI220     m363(.A0(mai_mai_n313_), .A1(mai_mai_n281_), .B0(mai_mai_n278_), .B1(mai_mai_n40_), .Y(mai_mai_n380_));
  INV        m364(.A(mai_mai_n348_), .Y(mai_mai_n381_));
  AOI220     m365(.A0(mai_mai_n381_), .A1(mai_mai_n89_), .B0(mai_mai_n380_), .B1(mai_mai_n148_), .Y(mai_mai_n382_));
  NO2        m366(.A(mai_mai_n382_), .B(mai_mai_n50_), .Y(mai_mai_n383_));
  NO3        m367(.A(mai_mai_n383_), .B(mai_mai_n379_), .C(mai_mai_n372_), .Y(mai_mai_n384_));
  AOI210     m368(.A0(mai_mai_n384_), .A1(mai_mai_n371_), .B0(mai_mai_n25_), .Y(mai_mai_n385_));
  NA4        m369(.A(mai_mai_n30_), .B(mai_mai_n89_), .C(x2), .D(mai_mai_n17_), .Y(mai_mai_n386_));
  NO3        m370(.A(mai_mai_n64_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n387_));
  NA2        m371(.A(mai_mai_n387_), .B(mai_mai_n248_), .Y(mai_mai_n388_));
  NO2        m372(.A(mai_mai_n388_), .B(mai_mai_n100_), .Y(mai_mai_n389_));
  NO3        m373(.A(mai_mai_n252_), .B(mai_mai_n170_), .C(mai_mai_n37_), .Y(mai_mai_n390_));
  OAI210     m374(.A0(mai_mai_n390_), .A1(mai_mai_n389_), .B0(x7), .Y(mai_mai_n391_));
  NA2        m375(.A(mai_mai_n213_), .B(x7), .Y(mai_mai_n392_));
  NA3        m376(.A(mai_mai_n392_), .B(mai_mai_n147_), .C(mai_mai_n129_), .Y(mai_mai_n393_));
  NA3        m377(.A(mai_mai_n393_), .B(mai_mai_n391_), .C(mai_mai_n386_), .Y(mai_mai_n394_));
  OAI210     m378(.A0(mai_mai_n394_), .A1(mai_mai_n385_), .B0(mai_mai_n35_), .Y(mai_mai_n395_));
  NA2        m379(.A(mai_mai_n325_), .B(mai_mai_n171_), .Y(mai_mai_n396_));
  NO2        m380(.A(mai_mai_n156_), .B(mai_mai_n40_), .Y(mai_mai_n397_));
  NA2        m381(.A(x3), .B(mai_mai_n50_), .Y(mai_mai_n398_));
  AOI210     m382(.A0(x2), .A1(mai_mai_n27_), .B0(mai_mai_n68_), .Y(mai_mai_n399_));
  NO3        m383(.A(mai_mai_n375_), .B(x3), .C(mai_mai_n50_), .Y(mai_mai_n400_));
  NO2        m384(.A(mai_mai_n400_), .B(mai_mai_n399_), .Y(mai_mai_n401_));
  OAI210     m385(.A0(mai_mai_n149_), .A1(mai_mai_n398_), .B0(mai_mai_n401_), .Y(mai_mai_n402_));
  AOI220     m386(.A0(mai_mai_n402_), .A1(x0), .B0(mai_mai_n397_), .B1(mai_mai_n130_), .Y(mai_mai_n403_));
  AOI210     m387(.A0(mai_mai_n403_), .A1(mai_mai_n396_), .B0(mai_mai_n221_), .Y(mai_mai_n404_));
  INV        m388(.A(x5), .Y(mai_mai_n405_));
  NO4        m389(.A(mai_mai_n103_), .B(mai_mai_n405_), .C(mai_mai_n56_), .D(mai_mai_n31_), .Y(mai_mai_n406_));
  NO2        m390(.A(mai_mai_n406_), .B(mai_mai_n404_), .Y(mai_mai_n407_));
  NA3        m391(.A(mai_mai_n407_), .B(mai_mai_n395_), .C(mai_mai_n359_), .Y(mai_mai_n408_));
  AOI210     m392(.A0(mai_mai_n344_), .A1(mai_mai_n25_), .B0(mai_mai_n408_), .Y(mai05));
  INV        m393(.A(x4), .Y(mai_mai_n412_));
  INV        m394(.A(x6), .Y(mai_mai_n413_));
  INV        m395(.A(mai_mai_n74_), .Y(mai_mai_n414_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  INV        u005(.A(men_men_n19_), .Y(men_men_n22_));
  NA2        u006(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n23_));
  INV        u007(.A(x5), .Y(men_men_n24_));
  NA2        u008(.A(x7), .B(x6), .Y(men_men_n25_));
  NA2        u009(.A(x8), .B(x3), .Y(men_men_n26_));
  NA2        u010(.A(x4), .B(x2), .Y(men_men_n27_));
  NO4        u011(.A(men_men_n27_), .B(men_men_n26_), .C(men_men_n25_), .D(men_men_n24_), .Y(men_men_n28_));
  NO2        u012(.A(men_men_n28_), .B(men_men_n23_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  NOi21      u015(.An(men_men_n22_), .B(men_men_n29_), .Y(men00));
  NO2        u016(.A(x1), .B(x0), .Y(men_men_n33_));
  INV        u017(.A(x6), .Y(men_men_n34_));
  NO2        u018(.A(men_men_n34_), .B(men_men_n24_), .Y(men_men_n35_));
  AN2        u019(.A(x8), .B(x7), .Y(men_men_n36_));
  NA3        u020(.A(men_men_n36_), .B(men_men_n35_), .C(men_men_n33_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  AOI210     u022(.A0(men_men_n37_), .A1(men_men_n22_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n35_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n50_));
  NA2        u034(.A(men_men_n50_), .B(men_men_n33_), .Y(men_men_n51_));
  INV        u035(.A(x2), .Y(men_men_n52_));
  NO2        u036(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  OAI210     u039(.A0(men_men_n51_), .A1(men_men_n31_), .B0(men_men_n55_), .Y(men_men_n56_));
  NO3        u040(.A(men_men_n56_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u041(.A(x8), .B(x7), .Y(men_men_n58_));
  NA2        u042(.A(men_men_n41_), .B(x1), .Y(men_men_n59_));
  INV        u043(.A(x9), .Y(men_men_n60_));
  NO2        u044(.A(men_men_n60_), .B(men_men_n34_), .Y(men_men_n61_));
  INV        u045(.A(men_men_n61_), .Y(men_men_n62_));
  NO3        u046(.A(men_men_n62_), .B(men_men_n59_), .C(men_men_n58_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n59_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  OA210      u051(.A0(men_men_n66_), .A1(men_men_n65_), .B0(men_men_n64_), .Y(men_men_n68_));
  OAI210     u052(.A0(men_men_n42_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n54_), .A1(men_men_n20_), .B0(men_men_n69_), .Y(men_men_n70_));
  NAi31      u054(.An(x1), .B(x9), .C(x5), .Y(men_men_n71_));
  OAI220     u055(.A0(men_men_n71_), .A1(men_men_n41_), .B0(men_men_n70_), .B1(men_men_n68_), .Y(men_men_n72_));
  OAI210     u056(.A0(men_men_n72_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n73_));
  NA2        u057(.A(men_men_n46_), .B(x2), .Y(men_men_n74_));
  OAI210     u058(.A0(men_men_n74_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n75_));
  NA2        u059(.A(x5), .B(x3), .Y(men_men_n76_));
  NO2        u060(.A(x8), .B(x6), .Y(men_men_n77_));
  NO2        u061(.A(men_men_n76_), .B(men_men_n52_), .Y(men_men_n78_));
  NAi21      u062(.An(x4), .B(x3), .Y(men_men_n79_));
  INV        u063(.A(men_men_n79_), .Y(men_men_n80_));
  NO2        u064(.A(x4), .B(x2), .Y(men_men_n81_));
  NO2        u065(.A(men_men_n81_), .B(x3), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n79_), .B(men_men_n18_), .Y(men_men_n83_));
  NO3        u067(.A(men_men_n83_), .B(men_men_n78_), .C(men_men_n75_), .Y(men_men_n84_));
  NO4        u068(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .D(x1), .Y(men_men_n85_));
  INV        u069(.A(x4), .Y(men_men_n86_));
  NA2        u070(.A(men_men_n85_), .B(men_men_n86_), .Y(men_men_n87_));
  NA2        u071(.A(x3), .B(men_men_n18_), .Y(men_men_n88_));
  NO2        u072(.A(men_men_n88_), .B(men_men_n24_), .Y(men_men_n89_));
  INV        u073(.A(x8), .Y(men_men_n90_));
  NA2        u074(.A(x2), .B(x1), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n89_), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n25_), .Y(men_men_n94_));
  AOI210     u078(.A0(men_men_n54_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n95_));
  OAI210     u079(.A0(men_men_n43_), .A1(men_men_n35_), .B0(men_men_n46_), .Y(men_men_n96_));
  NO3        u080(.A(men_men_n96_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n97_));
  NA2        u081(.A(x4), .B(men_men_n41_), .Y(men_men_n98_));
  NO2        u082(.A(men_men_n46_), .B(men_men_n52_), .Y(men_men_n99_));
  OAI210     u083(.A0(men_men_n99_), .A1(men_men_n41_), .B0(men_men_n18_), .Y(men_men_n100_));
  AOI210     u084(.A0(men_men_n98_), .A1(men_men_n50_), .B0(men_men_n100_), .Y(men_men_n101_));
  NO2        u085(.A(x3), .B(x2), .Y(men_men_n102_));
  NA2        u086(.A(men_men_n102_), .B(men_men_n24_), .Y(men_men_n103_));
  AOI210     u087(.A0(x8), .A1(x6), .B0(men_men_n103_), .Y(men_men_n104_));
  NA2        u088(.A(men_men_n52_), .B(x1), .Y(men_men_n105_));
  OAI210     u089(.A0(men_men_n105_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n106_));
  NO4        u090(.A(men_men_n106_), .B(men_men_n104_), .C(men_men_n101_), .D(men_men_n97_), .Y(men_men_n107_));
  AO220      u091(.A0(men_men_n107_), .A1(men_men_n87_), .B0(men_men_n84_), .B1(men_men_n73_), .Y(men02));
  NO2        u092(.A(x3), .B(men_men_n52_), .Y(men_men_n109_));
  NA2        u093(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n110_));
  NA2        u094(.A(men_men_n41_), .B(x0), .Y(men_men_n111_));
  OAI210     u095(.A0(x4), .A1(men_men_n110_), .B0(men_men_n111_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n112_), .B(x1), .Y(men_men_n113_));
  NO3        u097(.A(men_men_n113_), .B(x7), .C(x5), .Y(men_men_n114_));
  NA2        u098(.A(x9), .B(x2), .Y(men_men_n115_));
  OR2        u099(.A(x8), .B(x0), .Y(men_men_n116_));
  NAi21      u100(.An(x2), .B(x8), .Y(men_men_n117_));
  INV        u101(.A(men_men_n117_), .Y(men_men_n118_));
  NO2        u102(.A(x4), .B(x1), .Y(men_men_n119_));
  NOi21      u103(.An(x0), .B(x1), .Y(men_men_n120_));
  NO3        u104(.A(x9), .B(x8), .C(x7), .Y(men_men_n121_));
  NOi21      u105(.An(x0), .B(x4), .Y(men_men_n122_));
  NAi21      u106(.An(x8), .B(x7), .Y(men_men_n123_));
  NO2        u107(.A(men_men_n123_), .B(men_men_n60_), .Y(men_men_n124_));
  AOI220     u108(.A0(men_men_n124_), .A1(men_men_n122_), .B0(men_men_n121_), .B1(men_men_n120_), .Y(men_men_n125_));
  NO2        u109(.A(men_men_n125_), .B(men_men_n76_), .Y(men_men_n126_));
  NO2        u110(.A(x5), .B(men_men_n46_), .Y(men_men_n127_));
  NA2        u111(.A(x2), .B(men_men_n18_), .Y(men_men_n128_));
  AOI210     u112(.A0(men_men_n128_), .A1(men_men_n105_), .B0(men_men_n111_), .Y(men_men_n129_));
  OAI210     u113(.A0(men_men_n129_), .A1(men_men_n33_), .B0(men_men_n127_), .Y(men_men_n130_));
  NAi21      u114(.An(x0), .B(x4), .Y(men_men_n131_));
  NO2        u115(.A(men_men_n131_), .B(x1), .Y(men_men_n132_));
  NO2        u116(.A(x7), .B(x0), .Y(men_men_n133_));
  NO2        u117(.A(men_men_n81_), .B(men_men_n99_), .Y(men_men_n134_));
  NO2        u118(.A(men_men_n134_), .B(x3), .Y(men_men_n135_));
  OAI210     u119(.A0(men_men_n133_), .A1(men_men_n132_), .B0(men_men_n135_), .Y(men_men_n136_));
  NA2        u120(.A(x5), .B(x0), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n46_), .B(x2), .Y(men_men_n138_));
  NA3        u122(.A(men_men_n136_), .B(men_men_n130_), .C(men_men_n34_), .Y(men_men_n139_));
  NO3        u123(.A(men_men_n139_), .B(men_men_n126_), .C(men_men_n114_), .Y(men_men_n140_));
  NO2        u124(.A(men_men_n27_), .B(men_men_n24_), .Y(men_men_n141_));
  AOI220     u125(.A0(men_men_n120_), .A1(men_men_n141_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n142_));
  NO2        u126(.A(men_men_n142_), .B(men_men_n58_), .Y(men_men_n143_));
  NA2        u127(.A(x7), .B(x3), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n98_), .B(x5), .Y(men_men_n145_));
  NO2        u129(.A(x9), .B(x7), .Y(men_men_n146_));
  NOi21      u130(.An(x8), .B(x0), .Y(men_men_n147_));
  OA210      u131(.A0(men_men_n146_), .A1(x1), .B0(men_men_n147_), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n41_), .B(x2), .Y(men_men_n149_));
  INV        u133(.A(x7), .Y(men_men_n150_));
  NA2        u134(.A(men_men_n150_), .B(men_men_n18_), .Y(men_men_n151_));
  AOI220     u135(.A0(men_men_n151_), .A1(men_men_n149_), .B0(men_men_n109_), .B1(men_men_n36_), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n24_), .B(x4), .Y(men_men_n153_));
  NO2        u137(.A(men_men_n153_), .B(men_men_n122_), .Y(men_men_n154_));
  NO2        u138(.A(men_men_n154_), .B(men_men_n152_), .Y(men_men_n155_));
  AOI210     u139(.A0(men_men_n148_), .A1(men_men_n145_), .B0(men_men_n155_), .Y(men_men_n156_));
  OAI210     u140(.A0(men_men_n144_), .A1(men_men_n48_), .B0(men_men_n156_), .Y(men_men_n157_));
  NA2        u141(.A(x5), .B(x1), .Y(men_men_n158_));
  INV        u142(.A(men_men_n158_), .Y(men_men_n159_));
  AOI210     u143(.A0(men_men_n159_), .A1(men_men_n122_), .B0(men_men_n34_), .Y(men_men_n160_));
  NO2        u144(.A(men_men_n60_), .B(men_men_n90_), .Y(men_men_n161_));
  NAi21      u145(.An(x2), .B(x7), .Y(men_men_n162_));
  NAi31      u146(.An(men_men_n76_), .B(men_men_n36_), .C(men_men_n33_), .Y(men_men_n163_));
  NA2        u147(.A(men_men_n163_), .B(men_men_n160_), .Y(men_men_n164_));
  NO3        u148(.A(men_men_n164_), .B(men_men_n157_), .C(men_men_n143_), .Y(men_men_n165_));
  NO2        u149(.A(men_men_n165_), .B(men_men_n140_), .Y(men_men_n166_));
  NO2        u150(.A(men_men_n137_), .B(men_men_n134_), .Y(men_men_n167_));
  NA2        u151(.A(men_men_n24_), .B(men_men_n18_), .Y(men_men_n168_));
  NA2        u152(.A(men_men_n24_), .B(men_men_n17_), .Y(men_men_n169_));
  NA3        u153(.A(men_men_n169_), .B(men_men_n168_), .C(men_men_n23_), .Y(men_men_n170_));
  AN2        u154(.A(men_men_n170_), .B(men_men_n138_), .Y(men_men_n171_));
  NA2        u155(.A(x8), .B(x0), .Y(men_men_n172_));
  NO2        u156(.A(men_men_n150_), .B(men_men_n24_), .Y(men_men_n173_));
  NO2        u157(.A(men_men_n120_), .B(x4), .Y(men_men_n174_));
  NA2        u158(.A(men_men_n174_), .B(men_men_n173_), .Y(men_men_n175_));
  AOI210     u159(.A0(men_men_n172_), .A1(men_men_n128_), .B0(men_men_n175_), .Y(men_men_n176_));
  NA2        u160(.A(x2), .B(x0), .Y(men_men_n177_));
  NA2        u161(.A(x4), .B(x1), .Y(men_men_n178_));
  NAi21      u162(.An(men_men_n119_), .B(men_men_n178_), .Y(men_men_n179_));
  NOi31      u163(.An(men_men_n179_), .B(men_men_n153_), .C(men_men_n177_), .Y(men_men_n180_));
  NO4        u164(.A(men_men_n180_), .B(men_men_n176_), .C(men_men_n171_), .D(men_men_n167_), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n181_), .B(men_men_n41_), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n170_), .B(men_men_n74_), .Y(men_men_n183_));
  INV        u167(.A(men_men_n127_), .Y(men_men_n184_));
  NO2        u168(.A(men_men_n105_), .B(men_men_n17_), .Y(men_men_n185_));
  AOI210     u169(.A0(men_men_n33_), .A1(men_men_n90_), .B0(men_men_n185_), .Y(men_men_n186_));
  NO3        u170(.A(men_men_n186_), .B(men_men_n184_), .C(x7), .Y(men_men_n187_));
  NA3        u171(.A(men_men_n179_), .B(men_men_n184_), .C(men_men_n40_), .Y(men_men_n188_));
  OAI210     u172(.A0(men_men_n169_), .A1(men_men_n134_), .B0(men_men_n188_), .Y(men_men_n189_));
  NO3        u173(.A(men_men_n189_), .B(men_men_n187_), .C(men_men_n183_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n190_), .B(x3), .Y(men_men_n191_));
  NO3        u175(.A(men_men_n191_), .B(men_men_n182_), .C(men_men_n166_), .Y(men03));
  NO2        u176(.A(men_men_n46_), .B(x3), .Y(men_men_n193_));
  NO2        u177(.A(x6), .B(men_men_n24_), .Y(men_men_n194_));
  INV        u178(.A(men_men_n194_), .Y(men_men_n195_));
  NO2        u179(.A(men_men_n52_), .B(x1), .Y(men_men_n196_));
  OAI210     u180(.A0(men_men_n196_), .A1(men_men_n24_), .B0(men_men_n61_), .Y(men_men_n197_));
  OAI220     u181(.A0(men_men_n197_), .A1(men_men_n17_), .B0(men_men_n195_), .B1(men_men_n105_), .Y(men_men_n198_));
  NA2        u182(.A(men_men_n198_), .B(men_men_n193_), .Y(men_men_n199_));
  NA2        u183(.A(x6), .B(men_men_n24_), .Y(men_men_n200_));
  NO2        u184(.A(men_men_n200_), .B(x4), .Y(men_men_n201_));
  NO2        u185(.A(men_men_n18_), .B(x0), .Y(men_men_n202_));
  NA2        u186(.A(x3), .B(men_men_n17_), .Y(men_men_n203_));
  NO2        u187(.A(men_men_n203_), .B(men_men_n200_), .Y(men_men_n204_));
  NA2        u188(.A(x9), .B(men_men_n52_), .Y(men_men_n205_));
  NA2        u189(.A(men_men_n205_), .B(x4), .Y(men_men_n206_));
  NA2        u190(.A(men_men_n200_), .B(men_men_n79_), .Y(men_men_n207_));
  AOI210     u191(.A0(men_men_n24_), .A1(x3), .B0(men_men_n177_), .Y(men_men_n208_));
  AOI220     u192(.A0(men_men_n208_), .A1(men_men_n207_), .B0(men_men_n206_), .B1(men_men_n204_), .Y(men_men_n209_));
  NO2        u193(.A(x5), .B(x1), .Y(men_men_n210_));
  AOI220     u194(.A0(men_men_n210_), .A1(men_men_n17_), .B0(men_men_n102_), .B1(x5), .Y(men_men_n211_));
  NO2        u195(.A(men_men_n203_), .B(men_men_n168_), .Y(men_men_n212_));
  NO3        u196(.A(x3), .B(x2), .C(x1), .Y(men_men_n213_));
  NO2        u197(.A(men_men_n213_), .B(men_men_n212_), .Y(men_men_n214_));
  OAI210     u198(.A0(men_men_n211_), .A1(men_men_n62_), .B0(men_men_n214_), .Y(men_men_n215_));
  NA2        u199(.A(men_men_n215_), .B(men_men_n46_), .Y(men_men_n216_));
  NA3        u200(.A(men_men_n216_), .B(men_men_n209_), .C(men_men_n199_), .Y(men_men_n217_));
  NO2        u201(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n218_));
  NA2        u202(.A(men_men_n218_), .B(men_men_n19_), .Y(men_men_n219_));
  NO2        u203(.A(x3), .B(men_men_n17_), .Y(men_men_n220_));
  NO2        u204(.A(men_men_n220_), .B(x6), .Y(men_men_n221_));
  NOi21      u205(.An(men_men_n81_), .B(men_men_n221_), .Y(men_men_n222_));
  NO2        u206(.A(men_men_n222_), .B(men_men_n150_), .Y(men_men_n223_));
  OR2        u207(.A(men_men_n223_), .B(men_men_n173_), .Y(men_men_n224_));
  NA2        u208(.A(men_men_n41_), .B(men_men_n52_), .Y(men_men_n225_));
  INV        u209(.A(men_men_n169_), .Y(men_men_n226_));
  NO2        u210(.A(men_men_n178_), .B(x6), .Y(men_men_n227_));
  AOI220     u211(.A0(men_men_n227_), .A1(men_men_n226_), .B0(men_men_n138_), .B1(men_men_n89_), .Y(men_men_n228_));
  NA2        u212(.A(x6), .B(men_men_n46_), .Y(men_men_n229_));
  NO2        u213(.A(men_men_n229_), .B(men_men_n76_), .Y(men_men_n230_));
  NO2        u214(.A(men_men_n158_), .B(men_men_n41_), .Y(men_men_n231_));
  OAI210     u215(.A0(men_men_n231_), .A1(men_men_n212_), .B0(men_men_n432_), .Y(men_men_n232_));
  NA2        u216(.A(men_men_n194_), .B(men_men_n132_), .Y(men_men_n233_));
  NA3        u217(.A(men_men_n203_), .B(men_men_n127_), .C(x6), .Y(men_men_n234_));
  OAI210     u218(.A0(men_men_n90_), .A1(men_men_n34_), .B0(men_men_n65_), .Y(men_men_n235_));
  NA4        u219(.A(men_men_n235_), .B(men_men_n234_), .C(men_men_n233_), .D(men_men_n232_), .Y(men_men_n236_));
  OAI210     u220(.A0(men_men_n236_), .A1(men_men_n230_), .B0(x2), .Y(men_men_n237_));
  NA3        u221(.A(men_men_n237_), .B(men_men_n228_), .C(men_men_n224_), .Y(men_men_n238_));
  AOI210     u222(.A0(men_men_n217_), .A1(x8), .B0(men_men_n238_), .Y(men_men_n239_));
  NO2        u223(.A(men_men_n90_), .B(x3), .Y(men_men_n240_));
  NA2        u224(.A(men_men_n240_), .B(men_men_n201_), .Y(men_men_n241_));
  NO3        u225(.A(men_men_n88_), .B(men_men_n77_), .C(men_men_n24_), .Y(men_men_n242_));
  AOI210     u226(.A0(men_men_n221_), .A1(men_men_n153_), .B0(men_men_n242_), .Y(men_men_n243_));
  AOI210     u227(.A0(men_men_n243_), .A1(men_men_n241_), .B0(x2), .Y(men_men_n244_));
  NO2        u228(.A(x4), .B(men_men_n52_), .Y(men_men_n245_));
  AOI220     u229(.A0(men_men_n201_), .A1(men_men_n185_), .B0(men_men_n245_), .B1(men_men_n65_), .Y(men_men_n246_));
  NA2        u230(.A(men_men_n60_), .B(x6), .Y(men_men_n247_));
  NA3        u231(.A(men_men_n24_), .B(x3), .C(x2), .Y(men_men_n248_));
  AOI210     u232(.A0(men_men_n248_), .A1(men_men_n137_), .B0(men_men_n247_), .Y(men_men_n249_));
  NA2        u233(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n250_));
  NO2        u234(.A(men_men_n250_), .B(men_men_n24_), .Y(men_men_n251_));
  OAI210     u235(.A0(men_men_n251_), .A1(men_men_n249_), .B0(men_men_n119_), .Y(men_men_n252_));
  NA2        u236(.A(men_men_n203_), .B(x6), .Y(men_men_n253_));
  NO2        u237(.A(men_men_n203_), .B(x6), .Y(men_men_n254_));
  NA2        u238(.A(men_men_n253_), .B(men_men_n141_), .Y(men_men_n255_));
  NA4        u239(.A(men_men_n255_), .B(men_men_n252_), .C(men_men_n246_), .D(men_men_n150_), .Y(men_men_n256_));
  NA2        u240(.A(men_men_n194_), .B(men_men_n220_), .Y(men_men_n257_));
  NO2        u241(.A(x9), .B(x6), .Y(men_men_n258_));
  NO2        u242(.A(men_men_n137_), .B(men_men_n18_), .Y(men_men_n259_));
  NAi21      u243(.An(men_men_n259_), .B(men_men_n248_), .Y(men_men_n260_));
  NAi21      u244(.An(x1), .B(x4), .Y(men_men_n261_));
  AOI210     u245(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n262_));
  OAI210     u246(.A0(men_men_n137_), .A1(x3), .B0(men_men_n262_), .Y(men_men_n263_));
  AOI220     u247(.A0(men_men_n263_), .A1(men_men_n261_), .B0(men_men_n260_), .B1(men_men_n258_), .Y(men_men_n264_));
  NA2        u248(.A(men_men_n264_), .B(men_men_n257_), .Y(men_men_n265_));
  NA2        u249(.A(men_men_n60_), .B(x2), .Y(men_men_n266_));
  NO2        u250(.A(men_men_n266_), .B(men_men_n257_), .Y(men_men_n267_));
  NO3        u251(.A(x9), .B(x6), .C(x0), .Y(men_men_n268_));
  NA2        u252(.A(men_men_n105_), .B(men_men_n24_), .Y(men_men_n269_));
  NA2        u253(.A(x6), .B(x2), .Y(men_men_n270_));
  NO2        u254(.A(men_men_n270_), .B(men_men_n168_), .Y(men_men_n271_));
  AOI210     u255(.A0(men_men_n269_), .A1(men_men_n268_), .B0(men_men_n271_), .Y(men_men_n272_));
  OAI220     u256(.A0(men_men_n272_), .A1(men_men_n41_), .B0(men_men_n174_), .B1(men_men_n44_), .Y(men_men_n273_));
  OAI210     u257(.A0(men_men_n273_), .A1(men_men_n267_), .B0(men_men_n265_), .Y(men_men_n274_));
  NO2        u258(.A(x3), .B(men_men_n200_), .Y(men_men_n275_));
  NA2        u259(.A(x4), .B(x0), .Y(men_men_n276_));
  NO2        u260(.A(men_men_n71_), .B(x6), .Y(men_men_n277_));
  AOI210     u261(.A0(men_men_n275_), .A1(men_men_n40_), .B0(men_men_n277_), .Y(men_men_n278_));
  AOI210     u262(.A0(men_men_n278_), .A1(men_men_n274_), .B0(x8), .Y(men_men_n279_));
  NA2        u263(.A(men_men_n259_), .B(x6), .Y(men_men_n280_));
  NA2        u264(.A(x4), .B(men_men_n20_), .Y(men_men_n281_));
  AOI210     u265(.A0(men_men_n281_), .A1(men_men_n280_), .B0(men_men_n225_), .Y(men_men_n282_));
  NO4        u266(.A(men_men_n282_), .B(men_men_n279_), .C(men_men_n256_), .D(men_men_n244_), .Y(men_men_n283_));
  NO2        u267(.A(men_men_n161_), .B(x1), .Y(men_men_n284_));
  NO3        u268(.A(men_men_n284_), .B(x3), .C(men_men_n34_), .Y(men_men_n285_));
  OAI210     u269(.A0(men_men_n285_), .A1(men_men_n254_), .B0(x2), .Y(men_men_n286_));
  OAI210     u270(.A0(x0), .A1(x6), .B0(men_men_n42_), .Y(men_men_n287_));
  AOI210     u271(.A0(men_men_n287_), .A1(men_men_n286_), .B0(men_men_n184_), .Y(men_men_n288_));
  NOi21      u272(.An(men_men_n270_), .B(men_men_n17_), .Y(men_men_n289_));
  NA3        u273(.A(men_men_n289_), .B(men_men_n210_), .C(men_men_n38_), .Y(men_men_n290_));
  AOI210     u274(.A0(men_men_n34_), .A1(men_men_n52_), .B0(x0), .Y(men_men_n291_));
  NA3        u275(.A(men_men_n291_), .B(men_men_n159_), .C(men_men_n31_), .Y(men_men_n292_));
  NA2        u276(.A(x3), .B(x2), .Y(men_men_n293_));
  AOI220     u277(.A0(men_men_n293_), .A1(men_men_n225_), .B0(men_men_n292_), .B1(men_men_n290_), .Y(men_men_n294_));
  NAi21      u278(.An(x4), .B(x0), .Y(men_men_n295_));
  NO3        u279(.A(men_men_n295_), .B(men_men_n42_), .C(x2), .Y(men_men_n296_));
  OAI210     u280(.A0(x6), .A1(men_men_n18_), .B0(men_men_n296_), .Y(men_men_n297_));
  OAI220     u281(.A0(men_men_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n298_));
  NO2        u282(.A(x9), .B(x8), .Y(men_men_n299_));
  NA3        u283(.A(men_men_n299_), .B(men_men_n34_), .C(men_men_n52_), .Y(men_men_n300_));
  OAI210     u284(.A0(men_men_n291_), .A1(men_men_n289_), .B0(men_men_n300_), .Y(men_men_n301_));
  AOI220     u285(.A0(men_men_n301_), .A1(men_men_n80_), .B0(men_men_n298_), .B1(men_men_n30_), .Y(men_men_n302_));
  AOI210     u286(.A0(men_men_n302_), .A1(men_men_n297_), .B0(men_men_n24_), .Y(men_men_n303_));
  NA3        u287(.A(men_men_n34_), .B(x1), .C(men_men_n17_), .Y(men_men_n304_));
  OAI210     u288(.A0(men_men_n291_), .A1(men_men_n289_), .B0(men_men_n304_), .Y(men_men_n305_));
  INV        u289(.A(men_men_n212_), .Y(men_men_n306_));
  NA2        u290(.A(men_men_n34_), .B(men_men_n41_), .Y(men_men_n307_));
  OR2        u291(.A(men_men_n307_), .B(men_men_n276_), .Y(men_men_n308_));
  OAI220     u292(.A0(men_men_n308_), .A1(men_men_n158_), .B0(men_men_n229_), .B1(men_men_n306_), .Y(men_men_n309_));
  AO210      u293(.A0(men_men_n305_), .A1(men_men_n145_), .B0(men_men_n309_), .Y(men_men_n310_));
  NO4        u294(.A(men_men_n310_), .B(men_men_n303_), .C(men_men_n294_), .D(men_men_n288_), .Y(men_men_n311_));
  OAI210     u295(.A0(men_men_n283_), .A1(men_men_n239_), .B0(men_men_n311_), .Y(men04));
  OAI210     u296(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n313_));
  NA3        u297(.A(men_men_n313_), .B(men_men_n268_), .C(men_men_n82_), .Y(men_men_n314_));
  NO2        u298(.A(x2), .B(x1), .Y(men_men_n315_));
  OAI210     u299(.A0(men_men_n250_), .A1(men_men_n315_), .B0(men_men_n34_), .Y(men_men_n316_));
  NO2        u300(.A(men_men_n315_), .B(men_men_n295_), .Y(men_men_n317_));
  AOI210     u301(.A0(men_men_n60_), .A1(x4), .B0(men_men_n110_), .Y(men_men_n318_));
  OAI210     u302(.A0(men_men_n318_), .A1(men_men_n317_), .B0(men_men_n240_), .Y(men_men_n319_));
  NO2        u303(.A(men_men_n266_), .B(men_men_n88_), .Y(men_men_n320_));
  NO2        u304(.A(men_men_n320_), .B(men_men_n34_), .Y(men_men_n321_));
  NO2        u305(.A(men_men_n293_), .B(men_men_n202_), .Y(men_men_n322_));
  INV        u306(.A(men_men_n88_), .Y(men_men_n323_));
  OAI210     u307(.A0(men_men_n323_), .A1(men_men_n322_), .B0(men_men_n90_), .Y(men_men_n324_));
  NA3        u308(.A(men_men_n324_), .B(men_men_n321_), .C(men_men_n319_), .Y(men_men_n325_));
  NA2        u309(.A(men_men_n325_), .B(men_men_n316_), .Y(men_men_n326_));
  NO2        u310(.A(men_men_n205_), .B(men_men_n111_), .Y(men_men_n327_));
  NO3        u311(.A(men_men_n247_), .B(men_men_n117_), .C(men_men_n18_), .Y(men_men_n328_));
  NO2        u312(.A(men_men_n328_), .B(men_men_n327_), .Y(men_men_n329_));
  NOi21      u313(.An(men_men_n147_), .B(men_men_n128_), .Y(men_men_n330_));
  AOI210     u314(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n331_));
  OAI220     u315(.A0(men_men_n331_), .A1(men_men_n307_), .B0(men_men_n266_), .B1(men_men_n304_), .Y(men_men_n332_));
  AOI210     u316(.A0(men_men_n330_), .A1(men_men_n61_), .B0(men_men_n332_), .Y(men_men_n333_));
  NA2        u317(.A(men_men_n320_), .B(men_men_n90_), .Y(men_men_n334_));
  NA3        u318(.A(men_men_n334_), .B(men_men_n333_), .C(men_men_n329_), .Y(men_men_n335_));
  OAI210     u319(.A0(x1), .A1(x3), .B0(men_men_n296_), .Y(men_men_n336_));
  NA2        u320(.A(men_men_n336_), .B(men_men_n150_), .Y(men_men_n337_));
  AOI210     u321(.A0(men_men_n335_), .A1(x4), .B0(men_men_n337_), .Y(men_men_n338_));
  NA3        u322(.A(men_men_n317_), .B(men_men_n205_), .C(men_men_n90_), .Y(men_men_n339_));
  XO2        u323(.A(x4), .B(x0), .Y(men_men_n340_));
  OAI210     u324(.A0(men_men_n340_), .A1(men_men_n115_), .B0(men_men_n261_), .Y(men_men_n341_));
  NA2        u325(.A(men_men_n341_), .B(x8), .Y(men_men_n342_));
  AOI210     u326(.A0(men_men_n342_), .A1(men_men_n339_), .B0(x3), .Y(men_men_n343_));
  NO2        u327(.A(men_men_n90_), .B(x4), .Y(men_men_n344_));
  NA2        u328(.A(men_men_n344_), .B(men_men_n42_), .Y(men_men_n345_));
  NO3        u329(.A(men_men_n340_), .B(men_men_n161_), .C(x2), .Y(men_men_n346_));
  NO3        u330(.A(x8), .B(men_men_n27_), .C(men_men_n23_), .Y(men_men_n347_));
  NO2        u331(.A(men_men_n347_), .B(men_men_n346_), .Y(men_men_n348_));
  NA4        u332(.A(men_men_n348_), .B(men_men_n345_), .C(men_men_n219_), .D(x6), .Y(men_men_n349_));
  NO2        u333(.A(men_men_n177_), .B(men_men_n90_), .Y(men_men_n350_));
  OR2        u334(.A(men_men_n344_), .B(x3), .Y(men_men_n351_));
  NO2        u335(.A(men_men_n147_), .B(men_men_n105_), .Y(men_men_n352_));
  AOI220     u336(.A0(men_men_n352_), .A1(men_men_n351_), .B0(men_men_n350_), .B1(men_men_n59_), .Y(men_men_n353_));
  NO2        u337(.A(men_men_n147_), .B(men_men_n79_), .Y(men_men_n354_));
  INV        u338(.A(men_men_n353_), .Y(men_men_n355_));
  OAI220     u339(.A0(men_men_n355_), .A1(x6), .B0(men_men_n349_), .B1(men_men_n343_), .Y(men_men_n356_));
  OAI210     u340(.A0(men_men_n61_), .A1(men_men_n46_), .B0(men_men_n40_), .Y(men_men_n357_));
  OAI210     u341(.A0(men_men_n357_), .A1(men_men_n90_), .B0(men_men_n308_), .Y(men_men_n358_));
  AOI210     u342(.A0(men_men_n358_), .A1(men_men_n18_), .B0(men_men_n150_), .Y(men_men_n359_));
  AO220      u343(.A0(men_men_n359_), .A1(men_men_n356_), .B0(men_men_n338_), .B1(men_men_n326_), .Y(men_men_n360_));
  NA2        u344(.A(men_men_n213_), .B(men_men_n47_), .Y(men_men_n361_));
  NA3        u345(.A(men_men_n361_), .B(men_men_n360_), .C(men_men_n314_), .Y(men_men_n362_));
  NA3        u346(.A(x2), .B(men_men_n193_), .C(men_men_n150_), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n363_), .B(men_men_n24_), .Y(men_men_n364_));
  NA3        u348(.A(men_men_n118_), .B(men_men_n218_), .C(x0), .Y(men_men_n365_));
  OAI210     u349(.A0(men_men_n193_), .A1(men_men_n66_), .B0(men_men_n202_), .Y(men_men_n366_));
  NA3        u350(.A(men_men_n196_), .B(men_men_n220_), .C(x8), .Y(men_men_n367_));
  AOI210     u351(.A0(men_men_n367_), .A1(men_men_n366_), .B0(men_men_n24_), .Y(men_men_n368_));
  AOI210     u352(.A0(men_men_n117_), .A1(men_men_n116_), .B0(men_men_n40_), .Y(men_men_n369_));
  NOi31      u353(.An(men_men_n369_), .B(x3), .C(men_men_n178_), .Y(men_men_n370_));
  OAI210     u354(.A0(men_men_n370_), .A1(men_men_n368_), .B0(men_men_n146_), .Y(men_men_n371_));
  NAi31      u355(.An(men_men_n48_), .B(men_men_n284_), .C(men_men_n173_), .Y(men_men_n372_));
  NA3        u356(.A(men_men_n372_), .B(men_men_n371_), .C(men_men_n365_), .Y(men_men_n373_));
  OAI210     u357(.A0(men_men_n373_), .A1(men_men_n364_), .B0(x6), .Y(men_men_n374_));
  INV        u358(.A(men_men_n133_), .Y(men_men_n375_));
  NA3        u359(.A(men_men_n53_), .B(men_men_n36_), .C(men_men_n30_), .Y(men_men_n376_));
  AOI220     u360(.A0(men_men_n376_), .A1(men_men_n375_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n377_));
  AOI220     u361(.A0(men_men_n433_), .A1(men_men_n218_), .B0(men_men_n193_), .B1(men_men_n150_), .Y(men_men_n378_));
  AOI210     u362(.A0(men_men_n124_), .A1(men_men_n245_), .B0(x1), .Y(men_men_n379_));
  OAI210     u363(.A0(men_men_n378_), .A1(x8), .B0(men_men_n379_), .Y(men_men_n380_));
  NAi31      u364(.An(x2), .B(x8), .C(x0), .Y(men_men_n381_));
  OAI210     u365(.A0(men_men_n381_), .A1(x4), .B0(men_men_n162_), .Y(men_men_n382_));
  NA3        u366(.A(men_men_n382_), .B(men_men_n144_), .C(x9), .Y(men_men_n383_));
  NO4        u367(.A(men_men_n123_), .B(men_men_n295_), .C(x9), .D(x2), .Y(men_men_n384_));
  NOi21      u368(.An(men_men_n121_), .B(men_men_n177_), .Y(men_men_n385_));
  NO3        u369(.A(men_men_n385_), .B(men_men_n384_), .C(men_men_n18_), .Y(men_men_n386_));
  NO3        u370(.A(x9), .B(men_men_n150_), .C(x0), .Y(men_men_n387_));
  AOI220     u371(.A0(men_men_n387_), .A1(men_men_n240_), .B0(men_men_n354_), .B1(men_men_n150_), .Y(men_men_n388_));
  NA4        u372(.A(men_men_n388_), .B(men_men_n386_), .C(men_men_n383_), .D(men_men_n48_), .Y(men_men_n389_));
  OAI210     u373(.A0(men_men_n380_), .A1(men_men_n377_), .B0(men_men_n389_), .Y(men_men_n390_));
  NOi31      u374(.An(men_men_n433_), .B(men_men_n31_), .C(x8), .Y(men_men_n391_));
  AOI210     u375(.A0(men_men_n36_), .A1(x9), .B0(men_men_n131_), .Y(men_men_n392_));
  NO3        u376(.A(men_men_n392_), .B(men_men_n121_), .C(men_men_n41_), .Y(men_men_n393_));
  AOI210     u377(.A0(men_men_n261_), .A1(men_men_n58_), .B0(men_men_n120_), .Y(men_men_n394_));
  NO2        u378(.A(men_men_n394_), .B(x3), .Y(men_men_n395_));
  NO3        u379(.A(men_men_n395_), .B(men_men_n393_), .C(x2), .Y(men_men_n396_));
  NO2        u380(.A(men_men_n396_), .B(men_men_n391_), .Y(men_men_n397_));
  AOI210     u381(.A0(men_men_n397_), .A1(men_men_n390_), .B0(men_men_n24_), .Y(men_men_n398_));
  NO3        u382(.A(men_men_n60_), .B(x4), .C(x1), .Y(men_men_n399_));
  NO3        u383(.A(men_men_n66_), .B(men_men_n18_), .C(x0), .Y(men_men_n400_));
  AOI220     u384(.A0(men_men_n400_), .A1(men_men_n262_), .B0(men_men_n399_), .B1(men_men_n369_), .Y(men_men_n401_));
  NO2        u385(.A(men_men_n401_), .B(men_men_n102_), .Y(men_men_n402_));
  NA2        u386(.A(men_men_n402_), .B(x7), .Y(men_men_n403_));
  NA2        u387(.A(x8), .B(x7), .Y(men_men_n404_));
  NA3        u388(.A(men_men_n404_), .B(men_men_n149_), .C(men_men_n132_), .Y(men_men_n405_));
  NA2        u389(.A(men_men_n405_), .B(men_men_n403_), .Y(men_men_n406_));
  OAI210     u390(.A0(men_men_n406_), .A1(men_men_n398_), .B0(men_men_n34_), .Y(men_men_n407_));
  NO2        u391(.A(men_men_n387_), .B(men_men_n202_), .Y(men_men_n408_));
  NO4        u392(.A(men_men_n408_), .B(men_men_n76_), .C(x4), .D(men_men_n52_), .Y(men_men_n409_));
  NA2        u393(.A(men_men_n250_), .B(men_men_n21_), .Y(men_men_n410_));
  NO2        u394(.A(men_men_n158_), .B(men_men_n133_), .Y(men_men_n411_));
  NA2        u395(.A(men_men_n411_), .B(men_men_n410_), .Y(men_men_n412_));
  AOI210     u396(.A0(men_men_n412_), .A1(men_men_n163_), .B0(men_men_n27_), .Y(men_men_n413_));
  AOI220     u397(.A0(x3), .A1(men_men_n90_), .B0(men_men_n147_), .B1(men_men_n196_), .Y(men_men_n414_));
  NA3        u398(.A(men_men_n414_), .B(men_men_n381_), .C(men_men_n88_), .Y(men_men_n415_));
  NA2        u399(.A(men_men_n415_), .B(men_men_n173_), .Y(men_men_n416_));
  OAI220     u400(.A0(x3), .A1(men_men_n67_), .B0(men_men_n158_), .B1(men_men_n41_), .Y(men_men_n417_));
  AOI210     u401(.A0(men_men_n162_), .A1(men_men_n26_), .B0(men_men_n71_), .Y(men_men_n418_));
  OAI210     u402(.A0(men_men_n146_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n419_));
  NO2        u403(.A(x3), .B(men_men_n52_), .Y(men_men_n420_));
  AOI210     u404(.A0(men_men_n420_), .A1(men_men_n419_), .B0(men_men_n418_), .Y(men_men_n421_));
  INV        u405(.A(men_men_n421_), .Y(men_men_n422_));
  AOI220     u406(.A0(men_men_n422_), .A1(x0), .B0(men_men_n417_), .B1(men_men_n133_), .Y(men_men_n423_));
  AOI210     u407(.A0(men_men_n423_), .A1(men_men_n416_), .B0(men_men_n229_), .Y(men_men_n424_));
  NA2        u408(.A(x9), .B(x5), .Y(men_men_n425_));
  NO4        u409(.A(men_men_n105_), .B(men_men_n425_), .C(men_men_n58_), .D(men_men_n31_), .Y(men_men_n426_));
  NO4        u410(.A(men_men_n426_), .B(men_men_n424_), .C(men_men_n413_), .D(men_men_n409_), .Y(men_men_n427_));
  NA3        u411(.A(men_men_n427_), .B(men_men_n407_), .C(men_men_n374_), .Y(men_men_n428_));
  AOI210     u412(.A0(men_men_n362_), .A1(men_men_n24_), .B0(men_men_n428_), .Y(men05));
  INV        u413(.A(x6), .Y(men_men_n432_));
  INV        u414(.A(x0), .Y(men_men_n433_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule