library verilog;
use verilog.vl_types.all;
entity contmisterioso_vlg_vec_tst is
end contmisterioso_vlg_vec_tst;
