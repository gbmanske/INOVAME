// Benchmark "top" written by ABC on Fri Jun 21 17:49:20 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n138_, new_new_n139_,
    new_new_n140_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1078_, new_new_n1079_,
    new_new_n1080_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(mai1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n51_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g0062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g0063(.A(i_6_), .Y(new_new_n86_));
  OR4        g0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g0065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g0066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  AOI210     g0067(.A0(new_new_n88_), .A1(new_new_n86_), .B0(new_new_n89_), .Y(new_new_n90_));
  OAI210     g0068(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n90_), .Y(new_new_n91_));
  NAi21      g0069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g0070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g0071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n63_), .Y(new_new_n94_));
  NA2        g0072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  INV        g0073(.A(new_new_n94_), .Y(new_new_n96_));
  AOI210     g0074(.A0(new_new_n96_), .A1(new_new_n91_), .B0(new_new_n80_), .Y(new_new_n97_));
  AN3        g0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n98_));
  NAi21      g0076(.An(i_6_), .B(i_11_), .Y(new_new_n99_));
  NO2        g0077(.A(i_5_), .B(i_8_), .Y(new_new_n100_));
  NOi21      g0078(.An(new_new_n100_), .B(new_new_n99_), .Y(new_new_n101_));
  AOI220     g0079(.A0(new_new_n101_), .A1(new_new_n62_), .B0(new_new_n98_), .B1(new_new_n32_), .Y(new_new_n102_));
  INV        g0080(.A(i_7_), .Y(new_new_n103_));
  NA2        g0081(.A(new_new_n47_), .B(new_new_n103_), .Y(new_new_n104_));
  NO2        g0082(.A(i_0_), .B(i_5_), .Y(new_new_n105_));
  NO2        g0083(.A(new_new_n105_), .B(new_new_n86_), .Y(new_new_n106_));
  NA2        g0084(.A(i_12_), .B(i_3_), .Y(new_new_n107_));
  INV        g0085(.A(new_new_n107_), .Y(new_new_n108_));
  NA3        g0086(.A(new_new_n108_), .B(new_new_n106_), .C(new_new_n104_), .Y(new_new_n109_));
  NAi21      g0087(.An(i_7_), .B(i_11_), .Y(new_new_n110_));
  AN2        g0088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g0089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g0090(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n113_));
  NO2        g0091(.A(i_8_), .B(new_new_n103_), .Y(new_new_n114_));
  NO3        g0092(.A(new_new_n114_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n115_));
  NA2        g0093(.A(i_12_), .B(i_7_), .Y(new_new_n116_));
  NA2        g0094(.A(i_11_), .B(i_12_), .Y(new_new_n117_));
  INV        g0095(.A(new_new_n117_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n118_), .B(new_new_n115_), .Y(new_new_n119_));
  NA3        g0097(.A(new_new_n119_), .B(new_new_n109_), .C(new_new_n102_), .Y(new_new_n120_));
  NOi21      g0098(.An(i_1_), .B(i_5_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n121_), .B(i_11_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n123_));
  NA2        g0101(.A(i_7_), .B(new_new_n25_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(new_new_n123_), .Y(new_new_n125_));
  NO2        g0103(.A(new_new_n125_), .B(new_new_n47_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n127_));
  NAi21      g0105(.An(i_3_), .B(i_8_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n62_), .Y(new_new_n129_));
  NOi31      g0107(.An(new_new_n129_), .B(new_new_n127_), .C(new_new_n126_), .Y(new_new_n130_));
  NO2        g0108(.A(i_1_), .B(new_new_n86_), .Y(new_new_n131_));
  NO2        g0109(.A(i_6_), .B(i_5_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(i_3_), .Y(new_new_n133_));
  AO210      g0111(.A0(new_new_n133_), .A1(new_new_n48_), .B0(new_new_n131_), .Y(new_new_n134_));
  OAI220     g0112(.A0(new_new_n134_), .A1(new_new_n110_), .B0(new_new_n130_), .B1(new_new_n122_), .Y(new_new_n135_));
  NO3        g0113(.A(new_new_n135_), .B(new_new_n120_), .C(new_new_n97_), .Y(new_new_n136_));
  NA3        g0114(.A(new_new_n136_), .B(new_new_n79_), .C(new_new_n56_), .Y(mai2));
  NO2        g0115(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n138_));
  NA2        g0116(.A(i_6_), .B(new_new_n25_), .Y(new_new_n139_));
  NA2        g0117(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n140_));
  NA4        g0118(.A(new_new_n140_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(mai0));
  AN2        g0119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(i_6_), .Y(new_new_n143_));
  NO2        g0121(.A(i_12_), .B(i_13_), .Y(new_new_n144_));
  NAi21      g0122(.An(i_5_), .B(i_11_), .Y(new_new_n145_));
  NOi21      g0123(.An(new_new_n144_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g0124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NA2        g0125(.A(i_2_), .B(i_3_), .Y(new_new_n148_));
  NO2        g0126(.A(new_new_n148_), .B(i_4_), .Y(new_new_n149_));
  NA3        g0127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  AN2        g0128(.A(new_new_n144_), .B(new_new_n83_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(new_new_n27_), .Y(new_new_n152_));
  NA2        g0130(.A(i_1_), .B(i_5_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n73_), .B(new_new_n47_), .Y(new_new_n154_));
  NA2        g0132(.A(new_new_n154_), .B(new_new_n36_), .Y(new_new_n155_));
  NO3        g0133(.A(new_new_n155_), .B(new_new_n153_), .C(new_new_n152_), .Y(new_new_n156_));
  OR2        g0134(.A(i_0_), .B(i_1_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n158_));
  NAi32      g0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NAi21      g0137(.An(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  NOi21      g0138(.An(i_4_), .B(i_10_), .Y(new_new_n161_));
  NA2        g0139(.A(new_new_n161_), .B(new_new_n40_), .Y(new_new_n162_));
  NO2        g0140(.A(i_3_), .B(i_5_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  OAI210     g0143(.A0(new_new_n165_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n166_));
  NO2        g0144(.A(new_new_n166_), .B(new_new_n156_), .Y(new_new_n167_));
  AOI210     g0145(.A0(new_new_n167_), .A1(new_new_n150_), .B0(new_new_n143_), .Y(new_new_n168_));
  NA3        g0146(.A(new_new_n73_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n169_));
  NA2        g0147(.A(i_3_), .B(new_new_n49_), .Y(new_new_n170_));
  NOi21      g0148(.An(i_4_), .B(i_9_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_11_), .B(i_13_), .Y(new_new_n172_));
  NA2        g0150(.A(new_new_n172_), .B(new_new_n171_), .Y(new_new_n173_));
  OR2        g0151(.A(new_new_n173_), .B(new_new_n170_), .Y(new_new_n174_));
  NO2        g0152(.A(i_4_), .B(i_5_), .Y(new_new_n175_));
  NAi21      g0153(.An(i_12_), .B(i_11_), .Y(new_new_n176_));
  NO2        g0154(.A(new_new_n176_), .B(i_13_), .Y(new_new_n177_));
  NA3        g0155(.A(new_new_n177_), .B(new_new_n175_), .C(new_new_n83_), .Y(new_new_n178_));
  AOI210     g0156(.A0(new_new_n178_), .A1(new_new_n174_), .B0(new_new_n169_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n180_));
  NA2        g0158(.A(new_new_n180_), .B(new_new_n47_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n36_), .B(i_5_), .Y(new_new_n182_));
  NAi31      g0160(.An(new_new_n182_), .B(new_new_n151_), .C(i_11_), .Y(new_new_n183_));
  NA2        g0161(.A(i_3_), .B(i_5_), .Y(new_new_n184_));
  OR2        g0162(.A(new_new_n184_), .B(new_new_n173_), .Y(new_new_n185_));
  AOI210     g0163(.A0(new_new_n185_), .A1(new_new_n183_), .B0(new_new_n181_), .Y(new_new_n186_));
  NO2        g0164(.A(new_new_n73_), .B(i_5_), .Y(new_new_n187_));
  NO2        g0165(.A(i_13_), .B(i_10_), .Y(new_new_n188_));
  NA3        g0166(.A(new_new_n188_), .B(new_new_n187_), .C(new_new_n45_), .Y(new_new_n189_));
  NO2        g0167(.A(i_2_), .B(i_1_), .Y(new_new_n190_));
  NA2        g0168(.A(new_new_n190_), .B(i_3_), .Y(new_new_n191_));
  NAi21      g0169(.An(i_4_), .B(i_12_), .Y(new_new_n192_));
  NO4        g0170(.A(new_new_n192_), .B(new_new_n191_), .C(new_new_n189_), .D(new_new_n25_), .Y(new_new_n193_));
  NO3        g0171(.A(new_new_n193_), .B(new_new_n186_), .C(new_new_n179_), .Y(new_new_n194_));
  INV        g0172(.A(i_8_), .Y(new_new_n195_));
  NO2        g0173(.A(new_new_n195_), .B(i_7_), .Y(new_new_n196_));
  NA2        g0174(.A(new_new_n196_), .B(i_6_), .Y(new_new_n197_));
  NO3        g0175(.A(i_3_), .B(new_new_n86_), .C(new_new_n49_), .Y(new_new_n198_));
  NA2        g0176(.A(new_new_n198_), .B(new_new_n114_), .Y(new_new_n199_));
  NO3        g0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n200_));
  NA3        g0178(.A(new_new_n200_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n201_));
  NO3        g0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n202_));
  OAI210     g0180(.A0(new_new_n98_), .A1(i_12_), .B0(new_new_n202_), .Y(new_new_n203_));
  AOI210     g0181(.A0(new_new_n203_), .A1(new_new_n201_), .B0(new_new_n199_), .Y(new_new_n204_));
  NO2        g0182(.A(i_3_), .B(i_8_), .Y(new_new_n205_));
  NO3        g0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n206_));
  NA3        g0184(.A(new_new_n206_), .B(new_new_n205_), .C(new_new_n40_), .Y(new_new_n207_));
  NO2        g0185(.A(new_new_n105_), .B(new_new_n58_), .Y(new_new_n208_));
  NO2        g0186(.A(i_13_), .B(i_9_), .Y(new_new_n209_));
  NA3        g0187(.A(new_new_n209_), .B(i_6_), .C(new_new_n195_), .Y(new_new_n210_));
  NAi21      g0188(.An(i_12_), .B(i_3_), .Y(new_new_n211_));
  NO2        g0189(.A(new_new_n45_), .B(i_5_), .Y(new_new_n212_));
  NO3        g0190(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n213_));
  NA3        g0191(.A(new_new_n213_), .B(new_new_n212_), .C(i_10_), .Y(new_new_n214_));
  NO2        g0192(.A(new_new_n214_), .B(new_new_n210_), .Y(new_new_n215_));
  AOI210     g0193(.A0(new_new_n215_), .A1(i_7_), .B0(new_new_n204_), .Y(new_new_n216_));
  OAI220     g0194(.A0(new_new_n216_), .A1(i_4_), .B0(new_new_n197_), .B1(new_new_n194_), .Y(new_new_n217_));
  NAi21      g0195(.An(i_12_), .B(i_7_), .Y(new_new_n218_));
  NA3        g0196(.A(i_13_), .B(new_new_n195_), .C(i_10_), .Y(new_new_n219_));
  NO2        g0197(.A(new_new_n219_), .B(new_new_n218_), .Y(new_new_n220_));
  NA2        g0198(.A(i_0_), .B(i_5_), .Y(new_new_n221_));
  NA2        g0199(.A(new_new_n221_), .B(new_new_n106_), .Y(new_new_n222_));
  OAI220     g0200(.A0(new_new_n222_), .A1(new_new_n191_), .B0(new_new_n181_), .B1(new_new_n133_), .Y(new_new_n223_));
  NAi31      g0201(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n36_), .B(i_13_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n226_));
  NO2        g0204(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n227_));
  NA3        g0205(.A(new_new_n227_), .B(new_new_n226_), .C(new_new_n225_), .Y(new_new_n228_));
  INV        g0206(.A(i_13_), .Y(new_new_n229_));
  NO2        g0207(.A(i_12_), .B(new_new_n229_), .Y(new_new_n230_));
  NA3        g0208(.A(new_new_n230_), .B(new_new_n200_), .C(new_new_n198_), .Y(new_new_n231_));
  OAI210     g0209(.A0(new_new_n228_), .A1(new_new_n224_), .B0(new_new_n231_), .Y(new_new_n232_));
  AOI220     g0210(.A0(new_new_n232_), .A1(new_new_n142_), .B0(new_new_n223_), .B1(new_new_n220_), .Y(new_new_n233_));
  NO2        g0211(.A(i_12_), .B(new_new_n37_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n184_), .B(i_4_), .Y(new_new_n235_));
  NA2        g0213(.A(new_new_n235_), .B(new_new_n234_), .Y(new_new_n236_));
  OR2        g0214(.A(i_8_), .B(i_7_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n237_), .B(new_new_n86_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n54_), .B(i_1_), .Y(new_new_n239_));
  NA2        g0217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  INV        g0218(.A(i_12_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n45_), .B(new_new_n241_), .Y(new_new_n242_));
  NO3        g0220(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n243_));
  NA2        g0221(.A(i_2_), .B(i_1_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n240_), .B(new_new_n236_), .Y(new_new_n245_));
  NO3        g0223(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n246_));
  NAi21      g0224(.An(i_4_), .B(i_3_), .Y(new_new_n247_));
  NO2        g0225(.A(new_new_n247_), .B(new_new_n75_), .Y(new_new_n248_));
  NO2        g0226(.A(i_0_), .B(i_6_), .Y(new_new_n249_));
  NOi41      g0227(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n250_));
  NA2        g0228(.A(new_new_n250_), .B(new_new_n249_), .Y(new_new_n251_));
  NO2        g0229(.A(new_new_n244_), .B(new_new_n184_), .Y(new_new_n252_));
  NAi21      g0230(.An(new_new_n251_), .B(new_new_n252_), .Y(new_new_n253_));
  INV        g0231(.A(new_new_n253_), .Y(new_new_n254_));
  AOI220     g0232(.A0(new_new_n254_), .A1(new_new_n40_), .B0(new_new_n245_), .B1(new_new_n209_), .Y(new_new_n255_));
  NO2        g0233(.A(i_11_), .B(new_new_n229_), .Y(new_new_n256_));
  NOi21      g0234(.An(i_1_), .B(i_6_), .Y(new_new_n257_));
  NAi21      g0235(.An(i_3_), .B(i_7_), .Y(new_new_n258_));
  NA2        g0236(.A(new_new_n241_), .B(i_9_), .Y(new_new_n259_));
  OR4        g0237(.A(new_new_n259_), .B(new_new_n258_), .C(new_new_n257_), .D(new_new_n187_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n261_));
  NO2        g0239(.A(i_12_), .B(i_3_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n73_), .B(i_5_), .Y(new_new_n263_));
  NA2        g0241(.A(i_3_), .B(i_9_), .Y(new_new_n264_));
  NAi21      g0242(.An(i_7_), .B(i_10_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n266_));
  NA3        g0244(.A(new_new_n266_), .B(new_new_n263_), .C(new_new_n64_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n267_), .B(new_new_n260_), .Y(new_new_n268_));
  NA3        g0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n269_));
  INV        g0247(.A(new_new_n143_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n241_), .B(i_13_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n271_), .B(new_new_n75_), .Y(new_new_n272_));
  AOI220     g0250(.A0(new_new_n272_), .A1(new_new_n270_), .B0(new_new_n268_), .B1(new_new_n256_), .Y(new_new_n273_));
  NO2        g0251(.A(new_new_n237_), .B(new_new_n37_), .Y(new_new_n274_));
  NA2        g0252(.A(i_12_), .B(i_6_), .Y(new_new_n275_));
  OR2        g0253(.A(i_13_), .B(i_9_), .Y(new_new_n276_));
  NO2        g0254(.A(new_new_n247_), .B(i_2_), .Y(new_new_n277_));
  NA2        g0255(.A(new_new_n256_), .B(i_9_), .Y(new_new_n278_));
  NA2        g0256(.A(new_new_n154_), .B(new_new_n63_), .Y(new_new_n279_));
  NO3        g0257(.A(i_11_), .B(new_new_n229_), .C(new_new_n25_), .Y(new_new_n280_));
  NO2        g0258(.A(new_new_n258_), .B(i_8_), .Y(new_new_n281_));
  NO2        g0259(.A(i_6_), .B(new_new_n49_), .Y(new_new_n282_));
  NA3        g0260(.A(new_new_n282_), .B(new_new_n281_), .C(new_new_n280_), .Y(new_new_n283_));
  NO3        g0261(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n284_));
  NA3        g0262(.A(new_new_n284_), .B(new_new_n274_), .C(new_new_n230_), .Y(new_new_n285_));
  AOI210     g0263(.A0(new_new_n285_), .A1(new_new_n283_), .B0(new_new_n279_), .Y(new_new_n286_));
  INV        g0264(.A(new_new_n286_), .Y(new_new_n287_));
  NA4        g0265(.A(new_new_n287_), .B(new_new_n273_), .C(new_new_n255_), .D(new_new_n233_), .Y(new_new_n288_));
  NO3        g0266(.A(i_12_), .B(new_new_n229_), .C(new_new_n37_), .Y(new_new_n289_));
  INV        g0267(.A(new_new_n289_), .Y(new_new_n290_));
  NA2        g0268(.A(i_8_), .B(new_new_n103_), .Y(new_new_n291_));
  NOi21      g0269(.An(new_new_n163_), .B(new_new_n86_), .Y(new_new_n292_));
  NO3        g0270(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n293_));
  AOI220     g0271(.A0(new_new_n293_), .A1(new_new_n198_), .B0(new_new_n292_), .B1(new_new_n239_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n294_), .B(new_new_n291_), .Y(new_new_n295_));
  NO3        g0273(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n296_));
  NO2        g0274(.A(new_new_n244_), .B(i_0_), .Y(new_new_n297_));
  AOI220     g0275(.A0(new_new_n297_), .A1(new_new_n196_), .B0(new_new_n296_), .B1(new_new_n142_), .Y(new_new_n298_));
  NA2        g0276(.A(new_new_n282_), .B(new_new_n26_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n299_), .B(new_new_n298_), .Y(new_new_n300_));
  NA2        g0278(.A(i_0_), .B(i_1_), .Y(new_new_n301_));
  NO2        g0279(.A(new_new_n301_), .B(i_2_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n59_), .B(i_6_), .Y(new_new_n303_));
  NA3        g0281(.A(new_new_n303_), .B(new_new_n302_), .C(new_new_n163_), .Y(new_new_n304_));
  OAI210     g0282(.A0(new_new_n165_), .A1(new_new_n143_), .B0(new_new_n304_), .Y(new_new_n305_));
  NO3        g0283(.A(new_new_n305_), .B(new_new_n300_), .C(new_new_n295_), .Y(new_new_n306_));
  NO2        g0284(.A(i_3_), .B(i_10_), .Y(new_new_n307_));
  NA3        g0285(.A(new_new_n307_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n308_));
  NO2        g0286(.A(i_2_), .B(new_new_n103_), .Y(new_new_n309_));
  NA2        g0287(.A(i_1_), .B(new_new_n36_), .Y(new_new_n310_));
  NO2        g0288(.A(new_new_n310_), .B(i_8_), .Y(new_new_n311_));
  NA2        g0289(.A(new_new_n311_), .B(new_new_n309_), .Y(new_new_n312_));
  AN2        g0290(.A(i_3_), .B(i_10_), .Y(new_new_n313_));
  NA4        g0291(.A(new_new_n313_), .B(new_new_n200_), .C(new_new_n177_), .D(new_new_n175_), .Y(new_new_n314_));
  NO2        g0292(.A(i_5_), .B(new_new_n37_), .Y(new_new_n315_));
  NO2        g0293(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n316_));
  OR2        g0294(.A(new_new_n312_), .B(new_new_n308_), .Y(new_new_n317_));
  OAI220     g0295(.A0(new_new_n317_), .A1(i_6_), .B0(new_new_n306_), .B1(new_new_n290_), .Y(new_new_n318_));
  NO4        g0296(.A(new_new_n318_), .B(new_new_n288_), .C(new_new_n217_), .D(new_new_n168_), .Y(new_new_n319_));
  NO3        g0297(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n320_));
  NO2        g0298(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n321_));
  NA2        g0299(.A(new_new_n297_), .B(new_new_n321_), .Y(new_new_n322_));
  NO3        g0300(.A(i_6_), .B(new_new_n195_), .C(i_7_), .Y(new_new_n323_));
  NA2        g0301(.A(new_new_n323_), .B(new_new_n200_), .Y(new_new_n324_));
  AOI210     g0302(.A0(new_new_n324_), .A1(new_new_n322_), .B0(new_new_n170_), .Y(new_new_n325_));
  NO2        g0303(.A(i_2_), .B(i_3_), .Y(new_new_n326_));
  OR2        g0304(.A(i_0_), .B(i_5_), .Y(new_new_n327_));
  NA2        g0305(.A(new_new_n221_), .B(new_new_n327_), .Y(new_new_n328_));
  NA4        g0306(.A(new_new_n328_), .B(new_new_n238_), .C(new_new_n326_), .D(i_1_), .Y(new_new_n329_));
  NA3        g0307(.A(new_new_n297_), .B(new_new_n292_), .C(new_new_n114_), .Y(new_new_n330_));
  NAi21      g0308(.An(i_8_), .B(i_7_), .Y(new_new_n331_));
  NO2        g0309(.A(new_new_n331_), .B(i_6_), .Y(new_new_n332_));
  NO2        g0310(.A(new_new_n157_), .B(new_new_n47_), .Y(new_new_n333_));
  NA3        g0311(.A(new_new_n333_), .B(new_new_n332_), .C(new_new_n163_), .Y(new_new_n334_));
  NA3        g0312(.A(new_new_n334_), .B(new_new_n330_), .C(new_new_n329_), .Y(new_new_n335_));
  OAI210     g0313(.A0(new_new_n335_), .A1(new_new_n325_), .B0(i_4_), .Y(new_new_n336_));
  NO2        g0314(.A(i_12_), .B(i_10_), .Y(new_new_n337_));
  NOi21      g0315(.An(i_5_), .B(i_0_), .Y(new_new_n338_));
  NO3        g0316(.A(new_new_n310_), .B(new_new_n338_), .C(new_new_n128_), .Y(new_new_n339_));
  NA4        g0317(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n340_));
  NA2        g0318(.A(new_new_n339_), .B(new_new_n337_), .Y(new_new_n341_));
  NO2        g0319(.A(i_6_), .B(i_8_), .Y(new_new_n342_));
  NOi21      g0320(.An(i_0_), .B(i_2_), .Y(new_new_n343_));
  AN2        g0321(.A(new_new_n343_), .B(new_new_n342_), .Y(new_new_n344_));
  NO2        g0322(.A(i_1_), .B(i_7_), .Y(new_new_n345_));
  AO220      g0323(.A0(new_new_n345_), .A1(new_new_n344_), .B0(new_new_n332_), .B1(new_new_n239_), .Y(new_new_n346_));
  NA3        g0324(.A(new_new_n346_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n347_));
  NA3        g0325(.A(new_new_n347_), .B(new_new_n341_), .C(new_new_n336_), .Y(new_new_n348_));
  NO3        g0326(.A(new_new_n237_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n349_));
  NO3        g0327(.A(new_new_n331_), .B(i_2_), .C(i_1_), .Y(new_new_n350_));
  OAI210     g0328(.A0(new_new_n350_), .A1(new_new_n349_), .B0(i_6_), .Y(new_new_n351_));
  NA3        g0329(.A(new_new_n257_), .B(new_new_n309_), .C(new_new_n195_), .Y(new_new_n352_));
  AOI210     g0330(.A0(new_new_n352_), .A1(new_new_n351_), .B0(new_new_n328_), .Y(new_new_n353_));
  NOi21      g0331(.An(new_new_n153_), .B(new_new_n106_), .Y(new_new_n354_));
  NA2        g0332(.A(new_new_n353_), .B(i_3_), .Y(new_new_n355_));
  INV        g0333(.A(new_new_n84_), .Y(new_new_n356_));
  NO2        g0334(.A(new_new_n301_), .B(new_new_n81_), .Y(new_new_n357_));
  NA2        g0335(.A(new_new_n357_), .B(new_new_n132_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n95_), .B(new_new_n195_), .Y(new_new_n359_));
  NA2        g0337(.A(new_new_n359_), .B(new_new_n63_), .Y(new_new_n360_));
  AOI210     g0338(.A0(new_new_n360_), .A1(new_new_n358_), .B0(new_new_n356_), .Y(new_new_n361_));
  NO2        g0339(.A(new_new_n195_), .B(i_9_), .Y(new_new_n362_));
  NA3        g0340(.A(new_new_n362_), .B(new_new_n208_), .C(new_new_n157_), .Y(new_new_n363_));
  NO2        g0341(.A(new_new_n361_), .B(new_new_n300_), .Y(new_new_n364_));
  AOI210     g0342(.A0(new_new_n364_), .A1(new_new_n355_), .B0(new_new_n162_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n348_), .A1(new_new_n320_), .B0(new_new_n365_), .Y(new_new_n366_));
  NOi32      g0344(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n367_));
  INV        g0345(.A(new_new_n367_), .Y(new_new_n368_));
  NAi21      g0346(.An(i_0_), .B(i_6_), .Y(new_new_n369_));
  NAi21      g0347(.An(i_1_), .B(i_5_), .Y(new_new_n370_));
  NA2        g0348(.A(new_new_n370_), .B(new_new_n369_), .Y(new_new_n371_));
  NA2        g0349(.A(new_new_n371_), .B(new_new_n25_), .Y(new_new_n372_));
  OAI210     g0350(.A0(new_new_n372_), .A1(new_new_n159_), .B0(new_new_n251_), .Y(new_new_n373_));
  NAi41      g0351(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n374_));
  OAI220     g0352(.A0(new_new_n374_), .A1(new_new_n370_), .B0(new_new_n224_), .B1(new_new_n159_), .Y(new_new_n375_));
  AOI210     g0353(.A0(new_new_n374_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n376_));
  NOi32      g0354(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n377_));
  OR2        g0355(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n378_));
  NO2        g0356(.A(i_1_), .B(new_new_n103_), .Y(new_new_n379_));
  NAi21      g0357(.An(i_3_), .B(i_4_), .Y(new_new_n380_));
  NO2        g0358(.A(new_new_n380_), .B(i_9_), .Y(new_new_n381_));
  AN2        g0359(.A(i_6_), .B(i_7_), .Y(new_new_n382_));
  OAI210     g0360(.A0(new_new_n382_), .A1(new_new_n379_), .B0(new_new_n381_), .Y(new_new_n383_));
  NA2        g0361(.A(i_2_), .B(i_7_), .Y(new_new_n384_));
  NO2        g0362(.A(new_new_n380_), .B(i_10_), .Y(new_new_n385_));
  NA3        g0363(.A(new_new_n385_), .B(new_new_n384_), .C(new_new_n249_), .Y(new_new_n386_));
  AOI210     g0364(.A0(new_new_n386_), .A1(new_new_n383_), .B0(new_new_n187_), .Y(new_new_n387_));
  AOI210     g0365(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n388_));
  OAI210     g0366(.A0(new_new_n388_), .A1(new_new_n190_), .B0(new_new_n385_), .Y(new_new_n389_));
  AOI220     g0367(.A0(new_new_n385_), .A1(new_new_n345_), .B0(new_new_n243_), .B1(new_new_n190_), .Y(new_new_n390_));
  AOI210     g0368(.A0(new_new_n390_), .A1(new_new_n389_), .B0(i_5_), .Y(new_new_n391_));
  NO4        g0369(.A(new_new_n391_), .B(new_new_n387_), .C(new_new_n378_), .D(new_new_n373_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n392_), .B(new_new_n368_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n394_));
  AN2        g0372(.A(i_12_), .B(i_5_), .Y(new_new_n395_));
  NO2        g0373(.A(i_4_), .B(new_new_n26_), .Y(new_new_n396_));
  NA2        g0374(.A(new_new_n396_), .B(new_new_n395_), .Y(new_new_n397_));
  NO2        g0375(.A(i_11_), .B(i_6_), .Y(new_new_n398_));
  NA3        g0376(.A(new_new_n398_), .B(new_new_n333_), .C(new_new_n229_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n399_), .B(new_new_n397_), .Y(new_new_n400_));
  NO2        g0378(.A(new_new_n247_), .B(i_5_), .Y(new_new_n401_));
  NO2        g0379(.A(i_5_), .B(i_10_), .Y(new_new_n402_));
  AOI220     g0380(.A0(new_new_n402_), .A1(new_new_n277_), .B0(new_new_n401_), .B1(new_new_n200_), .Y(new_new_n403_));
  NA2        g0381(.A(new_new_n144_), .B(new_new_n46_), .Y(new_new_n404_));
  NO2        g0382(.A(new_new_n404_), .B(new_new_n403_), .Y(new_new_n405_));
  OAI210     g0383(.A0(new_new_n405_), .A1(new_new_n400_), .B0(new_new_n394_), .Y(new_new_n406_));
  NO2        g0384(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n150_), .B(new_new_n86_), .Y(new_new_n408_));
  OAI210     g0386(.A0(new_new_n408_), .A1(new_new_n400_), .B0(new_new_n407_), .Y(new_new_n409_));
  NO3        g0387(.A(new_new_n86_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n410_));
  NO2        g0388(.A(i_3_), .B(new_new_n103_), .Y(new_new_n411_));
  NA4        g0389(.A(new_new_n307_), .B(new_new_n93_), .C(new_new_n75_), .D(new_new_n55_), .Y(new_new_n412_));
  NO2        g0390(.A(i_11_), .B(i_12_), .Y(new_new_n413_));
  NA2        g0391(.A(new_new_n413_), .B(new_new_n36_), .Y(new_new_n414_));
  NO2        g0392(.A(new_new_n412_), .B(new_new_n414_), .Y(new_new_n415_));
  NA2        g0393(.A(new_new_n402_), .B(new_new_n241_), .Y(new_new_n416_));
  NA3        g0394(.A(new_new_n114_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n417_));
  NO2        g0395(.A(new_new_n417_), .B(new_new_n224_), .Y(new_new_n418_));
  NAi21      g0396(.An(i_13_), .B(i_0_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n419_), .B(new_new_n244_), .Y(new_new_n420_));
  OAI210     g0398(.A0(new_new_n418_), .A1(new_new_n415_), .B0(new_new_n420_), .Y(new_new_n421_));
  NA3        g0399(.A(new_new_n421_), .B(new_new_n409_), .C(new_new_n406_), .Y(new_new_n422_));
  NA2        g0400(.A(new_new_n45_), .B(new_new_n229_), .Y(new_new_n423_));
  NO3        g0401(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n424_));
  NO2        g0402(.A(i_0_), .B(i_11_), .Y(new_new_n425_));
  INV        g0403(.A(i_5_), .Y(new_new_n426_));
  AN2        g0404(.A(i_1_), .B(i_6_), .Y(new_new_n427_));
  NOi21      g0405(.An(i_2_), .B(i_12_), .Y(new_new_n428_));
  NA2        g0406(.A(new_new_n428_), .B(new_new_n427_), .Y(new_new_n429_));
  NO2        g0407(.A(new_new_n429_), .B(new_new_n426_), .Y(new_new_n430_));
  NA2        g0408(.A(new_new_n142_), .B(i_9_), .Y(new_new_n431_));
  NO2        g0409(.A(new_new_n431_), .B(i_4_), .Y(new_new_n432_));
  NA2        g0410(.A(new_new_n430_), .B(new_new_n432_), .Y(new_new_n433_));
  NAi21      g0411(.An(i_9_), .B(i_4_), .Y(new_new_n434_));
  OR2        g0412(.A(i_13_), .B(i_10_), .Y(new_new_n435_));
  NO3        g0413(.A(new_new_n435_), .B(new_new_n117_), .C(new_new_n434_), .Y(new_new_n436_));
  OR2        g0414(.A(new_new_n219_), .B(new_new_n218_), .Y(new_new_n437_));
  NO2        g0415(.A(new_new_n103_), .B(new_new_n25_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n289_), .B(new_new_n438_), .Y(new_new_n439_));
  NA2        g0417(.A(new_new_n282_), .B(new_new_n213_), .Y(new_new_n440_));
  OAI220     g0418(.A0(new_new_n440_), .A1(new_new_n437_), .B0(new_new_n439_), .B1(new_new_n354_), .Y(new_new_n441_));
  INV        g0419(.A(new_new_n441_), .Y(new_new_n442_));
  AOI210     g0420(.A0(new_new_n442_), .A1(new_new_n433_), .B0(new_new_n26_), .Y(new_new_n443_));
  NA2        g0421(.A(new_new_n330_), .B(new_new_n329_), .Y(new_new_n444_));
  AOI220     g0422(.A0(new_new_n303_), .A1(new_new_n293_), .B0(new_new_n297_), .B1(new_new_n321_), .Y(new_new_n445_));
  NO2        g0423(.A(new_new_n445_), .B(new_new_n170_), .Y(new_new_n446_));
  NO2        g0424(.A(new_new_n184_), .B(new_new_n86_), .Y(new_new_n447_));
  AOI220     g0425(.A0(new_new_n447_), .A1(new_new_n302_), .B0(new_new_n284_), .B1(new_new_n213_), .Y(new_new_n448_));
  NO2        g0426(.A(new_new_n448_), .B(new_new_n291_), .Y(new_new_n449_));
  NO3        g0427(.A(new_new_n449_), .B(new_new_n446_), .C(new_new_n444_), .Y(new_new_n450_));
  NA2        g0428(.A(new_new_n198_), .B(new_new_n98_), .Y(new_new_n451_));
  NA3        g0429(.A(new_new_n333_), .B(new_new_n163_), .C(new_new_n86_), .Y(new_new_n452_));
  AOI210     g0430(.A0(new_new_n452_), .A1(new_new_n451_), .B0(new_new_n331_), .Y(new_new_n453_));
  NA2        g0431(.A(new_new_n195_), .B(i_10_), .Y(new_new_n454_));
  NA3        g0432(.A(new_new_n263_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n303_), .B(new_new_n239_), .Y(new_new_n456_));
  OAI220     g0434(.A0(new_new_n456_), .A1(new_new_n184_), .B0(new_new_n455_), .B1(new_new_n454_), .Y(new_new_n457_));
  NO2        g0435(.A(i_3_), .B(new_new_n49_), .Y(new_new_n458_));
  NA3        g0436(.A(new_new_n345_), .B(new_new_n344_), .C(new_new_n458_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n323_), .B(new_new_n328_), .Y(new_new_n460_));
  OAI210     g0438(.A0(new_new_n460_), .A1(new_new_n191_), .B0(new_new_n459_), .Y(new_new_n461_));
  NO3        g0439(.A(new_new_n461_), .B(new_new_n457_), .C(new_new_n453_), .Y(new_new_n462_));
  AOI210     g0440(.A0(new_new_n462_), .A1(new_new_n450_), .B0(new_new_n278_), .Y(new_new_n463_));
  NO4        g0441(.A(new_new_n463_), .B(new_new_n443_), .C(new_new_n422_), .D(new_new_n393_), .Y(new_new_n464_));
  NO2        g0442(.A(new_new_n63_), .B(i_4_), .Y(new_new_n465_));
  NO2        g0443(.A(new_new_n73_), .B(i_13_), .Y(new_new_n466_));
  NO2        g0444(.A(i_10_), .B(i_9_), .Y(new_new_n467_));
  NAi21      g0445(.An(i_12_), .B(i_8_), .Y(new_new_n468_));
  NO2        g0446(.A(new_new_n468_), .B(i_3_), .Y(new_new_n469_));
  NO2        g0447(.A(new_new_n47_), .B(i_4_), .Y(new_new_n470_));
  NA2        g0448(.A(new_new_n470_), .B(new_new_n106_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n471_), .B(new_new_n207_), .Y(new_new_n472_));
  NA2        g0450(.A(new_new_n316_), .B(i_0_), .Y(new_new_n473_));
  NO3        g0451(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n275_), .B(new_new_n99_), .Y(new_new_n475_));
  NA2        g0453(.A(new_new_n475_), .B(new_new_n474_), .Y(new_new_n476_));
  NA2        g0454(.A(i_8_), .B(i_9_), .Y(new_new_n477_));
  AOI210     g0455(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n478_));
  OR2        g0456(.A(new_new_n478_), .B(new_new_n477_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n289_), .B(new_new_n208_), .Y(new_new_n480_));
  NO2        g0458(.A(new_new_n480_), .B(new_new_n479_), .Y(new_new_n481_));
  NA2        g0459(.A(new_new_n256_), .B(new_new_n315_), .Y(new_new_n482_));
  NO3        g0460(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n483_));
  AOI210     g0461(.A0(new_new_n262_), .A1(new_new_n190_), .B0(new_new_n483_), .Y(new_new_n484_));
  NO2        g0462(.A(new_new_n484_), .B(new_new_n482_), .Y(new_new_n485_));
  NO3        g0463(.A(new_new_n485_), .B(new_new_n481_), .C(new_new_n472_), .Y(new_new_n486_));
  OR2        g0464(.A(new_new_n301_), .B(new_new_n210_), .Y(new_new_n487_));
  OA210      g0465(.A0(new_new_n363_), .A1(new_new_n103_), .B0(new_new_n304_), .Y(new_new_n488_));
  OA220      g0466(.A0(new_new_n488_), .A1(new_new_n162_), .B0(new_new_n487_), .B1(new_new_n236_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n98_), .B(i_13_), .Y(new_new_n490_));
  NA2        g0468(.A(new_new_n447_), .B(new_new_n394_), .Y(new_new_n491_));
  NO2        g0469(.A(i_2_), .B(i_13_), .Y(new_new_n492_));
  NA3        g0470(.A(new_new_n492_), .B(new_new_n161_), .C(new_new_n101_), .Y(new_new_n493_));
  OAI220     g0471(.A0(new_new_n493_), .A1(new_new_n241_), .B0(new_new_n491_), .B1(new_new_n490_), .Y(new_new_n494_));
  NO3        g0472(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n495_));
  NO2        g0473(.A(i_6_), .B(i_7_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n496_), .B(new_new_n495_), .Y(new_new_n497_));
  NO2        g0475(.A(i_11_), .B(i_1_), .Y(new_new_n498_));
  NO2        g0476(.A(new_new_n73_), .B(i_3_), .Y(new_new_n499_));
  OR2        g0477(.A(i_11_), .B(i_8_), .Y(new_new_n500_));
  NOi21      g0478(.An(i_2_), .B(i_7_), .Y(new_new_n501_));
  NAi31      g0479(.An(new_new_n500_), .B(new_new_n501_), .C(new_new_n499_), .Y(new_new_n502_));
  NO2        g0480(.A(new_new_n435_), .B(i_6_), .Y(new_new_n503_));
  NA3        g0481(.A(new_new_n503_), .B(new_new_n465_), .C(new_new_n75_), .Y(new_new_n504_));
  NO2        g0482(.A(new_new_n504_), .B(new_new_n502_), .Y(new_new_n505_));
  NO2        g0483(.A(i_3_), .B(new_new_n195_), .Y(new_new_n506_));
  NO2        g0484(.A(i_6_), .B(i_10_), .Y(new_new_n507_));
  NA4        g0485(.A(new_new_n507_), .B(new_new_n320_), .C(new_new_n506_), .D(new_new_n241_), .Y(new_new_n508_));
  NO2        g0486(.A(new_new_n508_), .B(new_new_n155_), .Y(new_new_n509_));
  NA3        g0487(.A(new_new_n250_), .B(new_new_n172_), .C(new_new_n132_), .Y(new_new_n510_));
  NA2        g0488(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n511_));
  NO2        g0489(.A(new_new_n157_), .B(i_3_), .Y(new_new_n512_));
  NAi31      g0490(.An(new_new_n511_), .B(new_new_n512_), .C(new_new_n230_), .Y(new_new_n513_));
  NA3        g0491(.A(new_new_n407_), .B(new_new_n180_), .C(new_new_n149_), .Y(new_new_n514_));
  NA3        g0492(.A(new_new_n514_), .B(new_new_n513_), .C(new_new_n510_), .Y(new_new_n515_));
  NO4        g0493(.A(new_new_n515_), .B(new_new_n509_), .C(new_new_n505_), .D(new_new_n494_), .Y(new_new_n516_));
  NA2        g0494(.A(new_new_n474_), .B(new_new_n395_), .Y(new_new_n517_));
  NA2        g0495(.A(new_new_n483_), .B(new_new_n402_), .Y(new_new_n518_));
  NO2        g0496(.A(new_new_n518_), .B(new_new_n228_), .Y(new_new_n519_));
  NAi21      g0497(.An(new_new_n219_), .B(new_new_n413_), .Y(new_new_n520_));
  NO2        g0498(.A(new_new_n26_), .B(i_5_), .Y(new_new_n521_));
  NO2        g0499(.A(i_0_), .B(new_new_n86_), .Y(new_new_n522_));
  NA3        g0500(.A(new_new_n522_), .B(new_new_n521_), .C(new_new_n142_), .Y(new_new_n523_));
  OR3        g0501(.A(new_new_n310_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n524_));
  NO2        g0502(.A(new_new_n524_), .B(new_new_n523_), .Y(new_new_n525_));
  NA2        g0503(.A(new_new_n27_), .B(i_10_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n320_), .B(new_new_n243_), .Y(new_new_n527_));
  OAI220     g0505(.A0(new_new_n527_), .A1(new_new_n455_), .B0(new_new_n526_), .B1(new_new_n490_), .Y(new_new_n528_));
  NA4        g0506(.A(new_new_n313_), .B(new_new_n227_), .C(new_new_n73_), .D(new_new_n241_), .Y(new_new_n529_));
  NO2        g0507(.A(new_new_n529_), .B(new_new_n497_), .Y(new_new_n530_));
  NO4        g0508(.A(new_new_n530_), .B(new_new_n528_), .C(new_new_n525_), .D(new_new_n519_), .Y(new_new_n531_));
  NA4        g0509(.A(new_new_n531_), .B(new_new_n516_), .C(new_new_n489_), .D(new_new_n486_), .Y(new_new_n532_));
  NA3        g0510(.A(new_new_n313_), .B(new_new_n177_), .C(new_new_n175_), .Y(new_new_n533_));
  OAI210     g0511(.A0(new_new_n308_), .A1(new_new_n182_), .B0(new_new_n533_), .Y(new_new_n534_));
  AN2        g0512(.A(new_new_n293_), .B(new_new_n238_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n535_), .B(new_new_n534_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n122_), .B(new_new_n113_), .Y(new_new_n537_));
  AN2        g0515(.A(new_new_n537_), .B(new_new_n474_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n320_), .B(new_new_n164_), .Y(new_new_n539_));
  OAI210     g0517(.A0(new_new_n539_), .A1(new_new_n236_), .B0(new_new_n314_), .Y(new_new_n540_));
  AOI220     g0518(.A0(new_new_n540_), .A1(new_new_n332_), .B0(new_new_n538_), .B1(new_new_n316_), .Y(new_new_n541_));
  NA2        g0519(.A(new_new_n395_), .B(new_new_n229_), .Y(new_new_n542_));
  NA2        g0520(.A(new_new_n367_), .B(new_new_n73_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n382_), .B(new_new_n377_), .Y(new_new_n544_));
  AO210      g0522(.A0(new_new_n543_), .A1(new_new_n542_), .B0(new_new_n544_), .Y(new_new_n545_));
  NO2        g0523(.A(new_new_n36_), .B(i_8_), .Y(new_new_n546_));
  AOI210     g0524(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n436_), .Y(new_new_n547_));
  NA2        g0525(.A(new_new_n547_), .B(new_new_n545_), .Y(new_new_n548_));
  INV        g0526(.A(new_new_n548_), .Y(new_new_n549_));
  NO2        g0527(.A(i_7_), .B(new_new_n201_), .Y(new_new_n550_));
  OR2        g0528(.A(new_new_n184_), .B(i_4_), .Y(new_new_n551_));
  NO2        g0529(.A(new_new_n551_), .B(new_new_n86_), .Y(new_new_n552_));
  NA2        g0530(.A(new_new_n552_), .B(new_new_n550_), .Y(new_new_n553_));
  NA4        g0531(.A(new_new_n553_), .B(new_new_n549_), .C(new_new_n541_), .D(new_new_n536_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n401_), .B(new_new_n302_), .Y(new_new_n555_));
  OAI210     g0533(.A0(new_new_n397_), .A1(new_new_n169_), .B0(new_new_n555_), .Y(new_new_n556_));
  NO2        g0534(.A(i_12_), .B(new_new_n195_), .Y(new_new_n557_));
  NA2        g0535(.A(new_new_n557_), .B(new_new_n229_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n1080_), .B(new_new_n558_), .Y(new_new_n559_));
  NOi31      g0537(.An(new_new_n323_), .B(new_new_n435_), .C(new_new_n38_), .Y(new_new_n560_));
  OAI210     g0538(.A0(new_new_n560_), .A1(new_new_n559_), .B0(new_new_n556_), .Y(new_new_n561_));
  NO2        g0539(.A(i_8_), .B(i_7_), .Y(new_new_n562_));
  OAI210     g0540(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n563_), .B(new_new_n227_), .Y(new_new_n564_));
  AOI220     g0542(.A0(new_new_n333_), .A1(new_new_n40_), .B0(new_new_n239_), .B1(new_new_n209_), .Y(new_new_n565_));
  OAI220     g0543(.A0(new_new_n565_), .A1(new_new_n551_), .B0(new_new_n564_), .B1(new_new_n247_), .Y(new_new_n566_));
  NA2        g0544(.A(new_new_n45_), .B(i_10_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n567_), .B(i_6_), .Y(new_new_n568_));
  NA3        g0546(.A(new_new_n568_), .B(new_new_n566_), .C(new_new_n562_), .Y(new_new_n569_));
  AOI220     g0547(.A0(new_new_n447_), .A1(new_new_n333_), .B0(new_new_n252_), .B1(new_new_n249_), .Y(new_new_n570_));
  OAI220     g0548(.A0(new_new_n570_), .A1(new_new_n271_), .B0(new_new_n490_), .B1(new_new_n133_), .Y(new_new_n571_));
  NA2        g0549(.A(new_new_n571_), .B(new_new_n274_), .Y(new_new_n572_));
  NOi31      g0550(.An(new_new_n297_), .B(new_new_n308_), .C(new_new_n182_), .Y(new_new_n573_));
  NA3        g0551(.A(new_new_n313_), .B(new_new_n175_), .C(new_new_n98_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n225_), .B(new_new_n45_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n157_), .B(i_5_), .Y(new_new_n576_));
  NA3        g0554(.A(new_new_n576_), .B(new_new_n423_), .C(new_new_n326_), .Y(new_new_n577_));
  OAI210     g0555(.A0(new_new_n577_), .A1(new_new_n575_), .B0(new_new_n574_), .Y(new_new_n578_));
  OAI210     g0556(.A0(new_new_n578_), .A1(new_new_n573_), .B0(new_new_n483_), .Y(new_new_n579_));
  NA4        g0557(.A(new_new_n579_), .B(new_new_n572_), .C(new_new_n569_), .D(new_new_n561_), .Y(new_new_n580_));
  NA3        g0558(.A(new_new_n221_), .B(new_new_n71_), .C(new_new_n45_), .Y(new_new_n581_));
  NA2        g0559(.A(new_new_n289_), .B(new_new_n84_), .Y(new_new_n582_));
  AOI210     g0560(.A0(new_new_n581_), .A1(new_new_n358_), .B0(new_new_n582_), .Y(new_new_n583_));
  NA2        g0561(.A(new_new_n303_), .B(new_new_n293_), .Y(new_new_n584_));
  NO2        g0562(.A(new_new_n584_), .B(new_new_n174_), .Y(new_new_n585_));
  NA2        g0563(.A(new_new_n227_), .B(new_new_n226_), .Y(new_new_n586_));
  NA2        g0564(.A(new_new_n467_), .B(new_new_n225_), .Y(new_new_n587_));
  NO2        g0565(.A(new_new_n586_), .B(new_new_n587_), .Y(new_new_n588_));
  AOI210     g0566(.A0(i_6_), .A1(new_new_n47_), .B0(new_new_n379_), .Y(new_new_n589_));
  NA2        g0567(.A(i_0_), .B(new_new_n49_), .Y(new_new_n590_));
  NA3        g0568(.A(new_new_n557_), .B(new_new_n280_), .C(new_new_n590_), .Y(new_new_n591_));
  NO2        g0569(.A(new_new_n589_), .B(new_new_n591_), .Y(new_new_n592_));
  NO4        g0570(.A(new_new_n592_), .B(new_new_n588_), .C(new_new_n585_), .D(new_new_n583_), .Y(new_new_n593_));
  NO4        g0571(.A(new_new_n257_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n594_));
  NO3        g0572(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n237_), .B(new_new_n36_), .Y(new_new_n596_));
  AN2        g0574(.A(new_new_n596_), .B(new_new_n595_), .Y(new_new_n597_));
  OA210      g0575(.A0(new_new_n597_), .A1(new_new_n594_), .B0(new_new_n367_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n435_), .B(i_1_), .Y(new_new_n599_));
  NOi31      g0577(.An(new_new_n599_), .B(new_new_n475_), .C(new_new_n73_), .Y(new_new_n600_));
  AN4        g0578(.A(new_new_n600_), .B(new_new_n432_), .C(new_new_n521_), .D(i_2_), .Y(new_new_n601_));
  NO2        g0579(.A(new_new_n445_), .B(new_new_n178_), .Y(new_new_n602_));
  NO3        g0580(.A(new_new_n602_), .B(new_new_n601_), .C(new_new_n598_), .Y(new_new_n603_));
  NOi21      g0581(.An(i_10_), .B(i_6_), .Y(new_new_n604_));
  NO2        g0582(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n605_));
  NO2        g0583(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n606_));
  NA2        g0584(.A(new_new_n323_), .B(new_new_n164_), .Y(new_new_n607_));
  AOI220     g0585(.A0(new_new_n607_), .A1(new_new_n456_), .B0(new_new_n185_), .B1(new_new_n183_), .Y(new_new_n608_));
  NOi31      g0586(.An(new_new_n146_), .B(i_1_), .C(new_new_n340_), .Y(new_new_n609_));
  NO2        g0587(.A(new_new_n609_), .B(new_new_n608_), .Y(new_new_n610_));
  NO2        g0588(.A(new_new_n543_), .B(new_new_n390_), .Y(new_new_n611_));
  INV        g0589(.A(new_new_n326_), .Y(new_new_n612_));
  NO2        g0590(.A(i_12_), .B(new_new_n86_), .Y(new_new_n613_));
  NA2        g0591(.A(new_new_n175_), .B(i_0_), .Y(new_new_n614_));
  NO3        g0592(.A(new_new_n614_), .B(new_new_n351_), .C(new_new_n308_), .Y(new_new_n615_));
  OR2        g0593(.A(i_2_), .B(i_5_), .Y(new_new_n616_));
  OR2        g0594(.A(new_new_n616_), .B(new_new_n427_), .Y(new_new_n617_));
  AOI210     g0595(.A0(new_new_n384_), .A1(new_new_n249_), .B0(new_new_n200_), .Y(new_new_n618_));
  AOI210     g0596(.A0(new_new_n618_), .A1(new_new_n617_), .B0(new_new_n520_), .Y(new_new_n619_));
  NO3        g0597(.A(new_new_n619_), .B(new_new_n615_), .C(new_new_n611_), .Y(new_new_n620_));
  NA4        g0598(.A(new_new_n620_), .B(new_new_n610_), .C(new_new_n603_), .D(new_new_n593_), .Y(new_new_n621_));
  NO4        g0599(.A(new_new_n621_), .B(new_new_n580_), .C(new_new_n554_), .D(new_new_n532_), .Y(new_new_n622_));
  NA4        g0600(.A(new_new_n622_), .B(new_new_n464_), .C(new_new_n366_), .D(new_new_n319_), .Y(mai7));
  NO2        g0601(.A(new_new_n95_), .B(new_new_n55_), .Y(new_new_n624_));
  NO2        g0602(.A(new_new_n110_), .B(new_new_n92_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n396_), .B(new_new_n625_), .Y(new_new_n626_));
  NA2        g0604(.A(new_new_n507_), .B(new_new_n84_), .Y(new_new_n627_));
  NA2        g0605(.A(i_11_), .B(new_new_n195_), .Y(new_new_n628_));
  INV        g0606(.A(new_new_n626_), .Y(new_new_n629_));
  NA3        g0607(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n241_), .B(i_4_), .Y(new_new_n631_));
  NA2        g0609(.A(new_new_n631_), .B(i_8_), .Y(new_new_n632_));
  NO2        g0610(.A(new_new_n107_), .B(new_new_n630_), .Y(new_new_n633_));
  NA2        g0611(.A(i_2_), .B(new_new_n86_), .Y(new_new_n634_));
  OAI210     g0612(.A0(new_new_n89_), .A1(new_new_n205_), .B0(new_new_n206_), .Y(new_new_n635_));
  NO2        g0613(.A(i_7_), .B(new_new_n37_), .Y(new_new_n636_));
  NA2        g0614(.A(i_4_), .B(i_8_), .Y(new_new_n637_));
  AOI210     g0615(.A0(new_new_n637_), .A1(new_new_n313_), .B0(new_new_n636_), .Y(new_new_n638_));
  OAI220     g0616(.A0(new_new_n638_), .A1(new_new_n634_), .B0(new_new_n635_), .B1(i_13_), .Y(new_new_n639_));
  NO4        g0617(.A(new_new_n639_), .B(new_new_n633_), .C(new_new_n629_), .D(new_new_n624_), .Y(new_new_n640_));
  AOI210     g0618(.A0(new_new_n128_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n641_));
  AOI210     g0619(.A0(new_new_n641_), .A1(new_new_n241_), .B0(new_new_n161_), .Y(new_new_n642_));
  OR2        g0620(.A(i_6_), .B(i_10_), .Y(new_new_n643_));
  NO2        g0621(.A(new_new_n643_), .B(new_new_n23_), .Y(new_new_n644_));
  OR3        g0622(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n645_));
  NO3        g0623(.A(new_new_n645_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n646_));
  INV        g0624(.A(new_new_n202_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n646_), .B(new_new_n644_), .Y(new_new_n648_));
  OA220      g0626(.A0(new_new_n648_), .A1(new_new_n612_), .B0(new_new_n642_), .B1(new_new_n276_), .Y(new_new_n649_));
  AOI210     g0627(.A0(new_new_n649_), .A1(new_new_n640_), .B0(new_new_n63_), .Y(new_new_n650_));
  NOi21      g0628(.An(i_11_), .B(i_7_), .Y(new_new_n651_));
  AO210      g0629(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n652_), .B(new_new_n651_), .Y(new_new_n653_));
  NA2        g0631(.A(new_new_n653_), .B(new_new_n209_), .Y(new_new_n654_));
  NA3        g0632(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n655_));
  NAi31      g0633(.An(new_new_n655_), .B(new_new_n218_), .C(i_11_), .Y(new_new_n656_));
  AOI210     g0634(.A0(new_new_n656_), .A1(new_new_n654_), .B0(new_new_n63_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n88_), .B(new_new_n63_), .Y(new_new_n658_));
  AO210      g0636(.A0(new_new_n658_), .A1(new_new_n390_), .B0(new_new_n41_), .Y(new_new_n659_));
  NA2        g0637(.A(new_new_n230_), .B(new_new_n63_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n63_), .B(i_9_), .Y(new_new_n661_));
  NO2        g0639(.A(i_1_), .B(i_12_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n660_), .B(new_new_n659_), .Y(new_new_n663_));
  OAI210     g0641(.A0(new_new_n663_), .A1(new_new_n657_), .B0(i_6_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n655_), .B(new_new_n110_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n665_), .B(new_new_n613_), .Y(new_new_n666_));
  NO2        g0644(.A(new_new_n241_), .B(new_new_n86_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n667_), .B(i_11_), .Y(new_new_n668_));
  NA2        g0646(.A(new_new_n666_), .B(new_new_n476_), .Y(new_new_n669_));
  NO4        g0647(.A(new_new_n218_), .B(new_new_n128_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n670_));
  NA2        g0648(.A(new_new_n670_), .B(new_new_n661_), .Y(new_new_n671_));
  NA2        g0649(.A(new_new_n241_), .B(i_6_), .Y(new_new_n672_));
  NA2        g0650(.A(i_1_), .B(new_new_n266_), .Y(new_new_n673_));
  OAI210     g0651(.A0(new_new_n673_), .A1(new_new_n45_), .B0(new_new_n671_), .Y(new_new_n674_));
  NA3        g0652(.A(new_new_n562_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n138_), .B(i_9_), .Y(new_new_n676_));
  NA3        g0654(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n677_));
  NO2        g0655(.A(new_new_n47_), .B(i_1_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n676_), .B(new_new_n1078_), .Y(new_new_n679_));
  NA3        g0657(.A(new_new_n661_), .B(new_new_n326_), .C(i_6_), .Y(new_new_n680_));
  NO2        g0658(.A(new_new_n680_), .B(new_new_n23_), .Y(new_new_n681_));
  AOI210     g0659(.A0(new_new_n498_), .A1(new_new_n438_), .B0(new_new_n246_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n682_), .B(new_new_n634_), .Y(new_new_n683_));
  NAi21      g0661(.An(new_new_n675_), .B(new_new_n94_), .Y(new_new_n684_));
  NA2        g0662(.A(new_new_n678_), .B(new_new_n275_), .Y(new_new_n685_));
  NO2        g0663(.A(i_11_), .B(new_new_n37_), .Y(new_new_n686_));
  NA2        g0664(.A(new_new_n686_), .B(new_new_n24_), .Y(new_new_n687_));
  OAI210     g0665(.A0(new_new_n687_), .A1(new_new_n685_), .B0(new_new_n684_), .Y(new_new_n688_));
  OR4        g0666(.A(new_new_n688_), .B(new_new_n683_), .C(new_new_n681_), .D(new_new_n679_), .Y(new_new_n689_));
  NO3        g0667(.A(new_new_n689_), .B(new_new_n674_), .C(new_new_n669_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n241_), .B(new_new_n103_), .Y(new_new_n691_));
  NO2        g0669(.A(new_new_n691_), .B(new_new_n651_), .Y(new_new_n692_));
  NA2        g0670(.A(new_new_n692_), .B(i_1_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n693_), .B(new_new_n645_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n434_), .B(new_new_n86_), .Y(new_new_n695_));
  NA2        g0673(.A(new_new_n694_), .B(new_new_n47_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n237_), .B(new_new_n45_), .Y(new_new_n697_));
  NO3        g0675(.A(new_new_n697_), .B(new_new_n316_), .C(new_new_n242_), .Y(new_new_n698_));
  NO2        g0676(.A(new_new_n117_), .B(new_new_n37_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n699_), .B(i_6_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n86_), .B(i_9_), .Y(new_new_n701_));
  NO2        g0679(.A(new_new_n701_), .B(new_new_n63_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n702_), .B(new_new_n662_), .Y(new_new_n703_));
  NO4        g0681(.A(new_new_n703_), .B(new_new_n700_), .C(new_new_n698_), .D(i_4_), .Y(new_new_n704_));
  NA2        g0682(.A(i_1_), .B(i_3_), .Y(new_new_n705_));
  INV        g0683(.A(new_new_n704_), .Y(new_new_n706_));
  NA4        g0684(.A(new_new_n706_), .B(new_new_n696_), .C(new_new_n690_), .D(new_new_n664_), .Y(new_new_n707_));
  NO3        g0685(.A(new_new_n500_), .B(i_3_), .C(i_7_), .Y(new_new_n708_));
  NOi21      g0686(.An(new_new_n708_), .B(i_10_), .Y(new_new_n709_));
  OA210      g0687(.A0(new_new_n709_), .A1(new_new_n250_), .B0(new_new_n86_), .Y(new_new_n710_));
  NA3        g0688(.A(new_new_n507_), .B(new_new_n546_), .C(new_new_n47_), .Y(new_new_n711_));
  NA3        g0689(.A(new_new_n161_), .B(new_new_n84_), .C(new_new_n86_), .Y(new_new_n712_));
  NA2        g0690(.A(new_new_n712_), .B(new_new_n711_), .Y(new_new_n713_));
  OAI210     g0691(.A0(new_new_n713_), .A1(new_new_n710_), .B0(i_1_), .Y(new_new_n714_));
  AOI210     g0692(.A0(new_new_n275_), .A1(new_new_n99_), .B0(i_1_), .Y(new_new_n715_));
  NO2        g0693(.A(new_new_n380_), .B(i_2_), .Y(new_new_n716_));
  NA2        g0694(.A(new_new_n716_), .B(new_new_n715_), .Y(new_new_n717_));
  OAI210     g0695(.A0(new_new_n680_), .A1(new_new_n468_), .B0(new_new_n717_), .Y(new_new_n718_));
  INV        g0696(.A(new_new_n718_), .Y(new_new_n719_));
  AOI210     g0697(.A0(new_new_n719_), .A1(new_new_n714_), .B0(i_13_), .Y(new_new_n720_));
  OR2        g0698(.A(i_11_), .B(i_7_), .Y(new_new_n721_));
  NA3        g0699(.A(new_new_n721_), .B(new_new_n108_), .C(new_new_n138_), .Y(new_new_n722_));
  AOI220     g0700(.A0(new_new_n492_), .A1(new_new_n161_), .B0(new_new_n470_), .B1(new_new_n138_), .Y(new_new_n723_));
  OAI210     g0701(.A0(new_new_n723_), .A1(new_new_n45_), .B0(new_new_n722_), .Y(new_new_n724_));
  NO2        g0702(.A(new_new_n55_), .B(i_12_), .Y(new_new_n725_));
  INV        g0703(.A(new_new_n725_), .Y(new_new_n726_));
  NO2        g0704(.A(new_new_n501_), .B(new_new_n24_), .Y(new_new_n727_));
  AOI220     g0705(.A0(new_new_n727_), .A1(new_new_n695_), .B0(new_new_n250_), .B1(new_new_n131_), .Y(new_new_n728_));
  OAI220     g0706(.A0(new_new_n728_), .A1(new_new_n41_), .B0(new_new_n726_), .B1(new_new_n95_), .Y(new_new_n729_));
  AOI210     g0707(.A0(new_new_n724_), .A1(new_new_n342_), .B0(new_new_n729_), .Y(new_new_n730_));
  NA2        g0708(.A(new_new_n398_), .B(new_new_n678_), .Y(new_new_n731_));
  NO2        g0709(.A(new_new_n731_), .B(new_new_n247_), .Y(new_new_n732_));
  AOI210     g0710(.A0(new_new_n468_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n733_));
  NOi31      g0711(.An(new_new_n733_), .B(new_new_n627_), .C(new_new_n45_), .Y(new_new_n734_));
  NA2        g0712(.A(new_new_n127_), .B(i_13_), .Y(new_new_n735_));
  NO2        g0713(.A(new_new_n677_), .B(new_new_n116_), .Y(new_new_n736_));
  INV        g0714(.A(new_new_n736_), .Y(new_new_n737_));
  OAI220     g0715(.A0(new_new_n737_), .A1(new_new_n71_), .B0(new_new_n735_), .B1(new_new_n715_), .Y(new_new_n738_));
  NA2        g0716(.A(new_new_n26_), .B(new_new_n195_), .Y(new_new_n739_));
  INV        g0717(.A(i_7_), .Y(new_new_n740_));
  AOI220     g0718(.A0(new_new_n398_), .A1(new_new_n678_), .B0(new_new_n94_), .B1(new_new_n104_), .Y(new_new_n741_));
  NO2        g0719(.A(new_new_n741_), .B(new_new_n632_), .Y(new_new_n742_));
  NO4        g0720(.A(new_new_n742_), .B(new_new_n738_), .C(new_new_n734_), .D(new_new_n732_), .Y(new_new_n743_));
  OR2        g0721(.A(i_11_), .B(i_6_), .Y(new_new_n744_));
  NA3        g0722(.A(new_new_n631_), .B(new_new_n739_), .C(i_7_), .Y(new_new_n745_));
  AOI210     g0723(.A0(new_new_n745_), .A1(new_new_n737_), .B0(new_new_n744_), .Y(new_new_n746_));
  NA3        g0724(.A(new_new_n428_), .B(new_new_n636_), .C(new_new_n99_), .Y(new_new_n747_));
  NA2        g0725(.A(new_new_n668_), .B(i_13_), .Y(new_new_n748_));
  NA2        g0726(.A(new_new_n104_), .B(new_new_n739_), .Y(new_new_n749_));
  NAi21      g0727(.An(i_11_), .B(i_12_), .Y(new_new_n750_));
  NOi41      g0728(.An(new_new_n112_), .B(new_new_n750_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n751_));
  NA2        g0729(.A(new_new_n751_), .B(new_new_n749_), .Y(new_new_n752_));
  NA3        g0730(.A(new_new_n752_), .B(new_new_n748_), .C(new_new_n747_), .Y(new_new_n753_));
  OAI210     g0731(.A0(new_new_n753_), .A1(new_new_n746_), .B0(new_new_n63_), .Y(new_new_n754_));
  NO2        g0732(.A(i_2_), .B(i_12_), .Y(new_new_n755_));
  NA2        g0733(.A(new_new_n379_), .B(new_new_n755_), .Y(new_new_n756_));
  NA2        g0734(.A(i_8_), .B(new_new_n25_), .Y(new_new_n757_));
  NO3        g0735(.A(new_new_n757_), .B(new_new_n396_), .C(new_new_n631_), .Y(new_new_n758_));
  OAI210     g0736(.A0(new_new_n758_), .A1(new_new_n381_), .B0(new_new_n379_), .Y(new_new_n759_));
  NO2        g0737(.A(new_new_n128_), .B(i_2_), .Y(new_new_n760_));
  NA2        g0738(.A(new_new_n759_), .B(new_new_n756_), .Y(new_new_n761_));
  NA3        g0739(.A(new_new_n761_), .B(new_new_n46_), .C(new_new_n229_), .Y(new_new_n762_));
  NA4        g0740(.A(new_new_n762_), .B(new_new_n754_), .C(new_new_n743_), .D(new_new_n730_), .Y(new_new_n763_));
  OR4        g0741(.A(new_new_n763_), .B(new_new_n720_), .C(new_new_n707_), .D(new_new_n650_), .Y(mai5));
  NA2        g0742(.A(new_new_n692_), .B(new_new_n277_), .Y(new_new_n765_));
  AN2        g0743(.A(new_new_n24_), .B(i_10_), .Y(new_new_n766_));
  NA3        g0744(.A(new_new_n766_), .B(new_new_n755_), .C(new_new_n110_), .Y(new_new_n767_));
  NO2        g0745(.A(new_new_n632_), .B(i_11_), .Y(new_new_n768_));
  NA2        g0746(.A(new_new_n89_), .B(new_new_n768_), .Y(new_new_n769_));
  NA3        g0747(.A(new_new_n769_), .B(new_new_n767_), .C(new_new_n765_), .Y(new_new_n770_));
  NO3        g0748(.A(i_11_), .B(new_new_n241_), .C(i_13_), .Y(new_new_n771_));
  NO2        g0749(.A(new_new_n124_), .B(new_new_n23_), .Y(new_new_n772_));
  NA2        g0750(.A(i_12_), .B(i_8_), .Y(new_new_n773_));
  OAI210     g0751(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n773_), .Y(new_new_n774_));
  INV        g0752(.A(new_new_n467_), .Y(new_new_n775_));
  AOI220     g0753(.A0(new_new_n326_), .A1(new_new_n606_), .B0(new_new_n774_), .B1(new_new_n772_), .Y(new_new_n776_));
  INV        g0754(.A(new_new_n776_), .Y(new_new_n777_));
  NO2        g0755(.A(new_new_n777_), .B(new_new_n770_), .Y(new_new_n778_));
  INV        g0756(.A(new_new_n172_), .Y(new_new_n779_));
  INV        g0757(.A(new_new_n250_), .Y(new_new_n780_));
  OAI210     g0758(.A0(new_new_n716_), .A1(new_new_n469_), .B0(new_new_n112_), .Y(new_new_n781_));
  AOI210     g0759(.A0(new_new_n781_), .A1(new_new_n780_), .B0(new_new_n779_), .Y(new_new_n782_));
  NO2        g0760(.A(new_new_n477_), .B(new_new_n26_), .Y(new_new_n783_));
  NO2        g0761(.A(new_new_n783_), .B(new_new_n438_), .Y(new_new_n784_));
  NA2        g0762(.A(new_new_n784_), .B(i_2_), .Y(new_new_n785_));
  INV        g0763(.A(new_new_n785_), .Y(new_new_n786_));
  AOI210     g0764(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n435_), .Y(new_new_n787_));
  AOI210     g0765(.A0(new_new_n787_), .A1(new_new_n786_), .B0(new_new_n782_), .Y(new_new_n788_));
  NO2        g0766(.A(new_new_n192_), .B(new_new_n125_), .Y(new_new_n789_));
  OAI210     g0767(.A0(new_new_n789_), .A1(new_new_n772_), .B0(i_2_), .Y(new_new_n790_));
  INV        g0768(.A(new_new_n173_), .Y(new_new_n791_));
  NO3        g0769(.A(new_new_n652_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n792_));
  AOI210     g0770(.A0(new_new_n791_), .A1(new_new_n89_), .B0(new_new_n792_), .Y(new_new_n793_));
  AOI210     g0771(.A0(new_new_n793_), .A1(new_new_n790_), .B0(new_new_n195_), .Y(new_new_n794_));
  OA210      g0772(.A0(new_new_n653_), .A1(new_new_n126_), .B0(i_13_), .Y(new_new_n795_));
  NA2        g0773(.A(new_new_n151_), .B(new_new_n628_), .Y(new_new_n796_));
  NO2        g0774(.A(new_new_n796_), .B(new_new_n384_), .Y(new_new_n797_));
  AOI210     g0775(.A0(new_new_n211_), .A1(new_new_n148_), .B0(new_new_n546_), .Y(new_new_n798_));
  OAI210     g0776(.A0(new_new_n798_), .A1(new_new_n230_), .B0(new_new_n438_), .Y(new_new_n799_));
  NO2        g0777(.A(new_new_n104_), .B(new_new_n45_), .Y(new_new_n800_));
  INV        g0778(.A(new_new_n309_), .Y(new_new_n801_));
  NA4        g0779(.A(new_new_n801_), .B(new_new_n313_), .C(new_new_n124_), .D(new_new_n43_), .Y(new_new_n802_));
  OAI210     g0780(.A0(new_new_n802_), .A1(new_new_n800_), .B0(new_new_n799_), .Y(new_new_n803_));
  NO4        g0781(.A(new_new_n803_), .B(new_new_n797_), .C(new_new_n795_), .D(new_new_n794_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n606_), .B(new_new_n28_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n771_), .B(new_new_n281_), .Y(new_new_n806_));
  NA2        g0784(.A(new_new_n806_), .B(new_new_n805_), .Y(new_new_n807_));
  NO2        g0785(.A(new_new_n62_), .B(i_12_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n808_), .B(new_new_n126_), .Y(new_new_n809_));
  NO2        g0787(.A(new_new_n809_), .B(new_new_n628_), .Y(new_new_n810_));
  AOI220     g0788(.A0(new_new_n810_), .A1(new_new_n36_), .B0(new_new_n807_), .B1(new_new_n47_), .Y(new_new_n811_));
  NA4        g0789(.A(new_new_n811_), .B(new_new_n804_), .C(new_new_n788_), .D(new_new_n778_), .Y(mai6));
  NO3        g0790(.A(new_new_n261_), .B(new_new_n315_), .C(i_1_), .Y(new_new_n813_));
  NO2        g0791(.A(new_new_n187_), .B(new_new_n139_), .Y(new_new_n814_));
  OAI210     g0792(.A0(new_new_n814_), .A1(new_new_n813_), .B0(new_new_n760_), .Y(new_new_n815_));
  NO2        g0793(.A(new_new_n224_), .B(new_new_n511_), .Y(new_new_n816_));
  NO2        g0794(.A(i_11_), .B(i_9_), .Y(new_new_n817_));
  AO210      g0795(.A0(new_new_n1079_), .A1(new_new_n815_), .B0(i_12_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n385_), .B(new_new_n345_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n613_), .B(new_new_n63_), .Y(new_new_n820_));
  NA2        g0798(.A(new_new_n709_), .B(new_new_n71_), .Y(new_new_n821_));
  BUFFER     g0799(.A(new_new_n658_), .Y(new_new_n822_));
  NA4        g0800(.A(new_new_n822_), .B(new_new_n821_), .C(new_new_n820_), .D(new_new_n819_), .Y(new_new_n823_));
  INV        g0801(.A(new_new_n199_), .Y(new_new_n824_));
  AOI220     g0802(.A0(new_new_n824_), .A1(new_new_n817_), .B0(new_new_n823_), .B1(new_new_n73_), .Y(new_new_n825_));
  INV        g0803(.A(new_new_n337_), .Y(new_new_n826_));
  NA2        g0804(.A(new_new_n75_), .B(new_new_n131_), .Y(new_new_n827_));
  INV        g0805(.A(new_new_n124_), .Y(new_new_n828_));
  NA2        g0806(.A(new_new_n828_), .B(new_new_n47_), .Y(new_new_n829_));
  AOI210     g0807(.A0(new_new_n829_), .A1(new_new_n827_), .B0(new_new_n826_), .Y(new_new_n830_));
  NO2        g0808(.A(new_new_n257_), .B(i_9_), .Y(new_new_n831_));
  NA2        g0809(.A(new_new_n831_), .B(new_new_n808_), .Y(new_new_n832_));
  AOI210     g0810(.A0(new_new_n832_), .A1(new_new_n544_), .B0(new_new_n187_), .Y(new_new_n833_));
  NO2        g0811(.A(new_new_n32_), .B(i_11_), .Y(new_new_n834_));
  NA3        g0812(.A(new_new_n834_), .B(new_new_n496_), .C(new_new_n402_), .Y(new_new_n835_));
  NAi32      g0813(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n836_));
  AOI210     g0814(.A0(new_new_n744_), .A1(new_new_n87_), .B0(new_new_n836_), .Y(new_new_n837_));
  OAI210     g0815(.A0(new_new_n708_), .A1(new_new_n596_), .B0(new_new_n595_), .Y(new_new_n838_));
  NAi31      g0816(.An(new_new_n837_), .B(new_new_n838_), .C(new_new_n835_), .Y(new_new_n839_));
  OR3        g0817(.A(new_new_n839_), .B(new_new_n833_), .C(new_new_n830_), .Y(new_new_n840_));
  NO2        g0818(.A(new_new_n721_), .B(i_2_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n842_));
  OAI210     g0820(.A0(new_new_n842_), .A1(new_new_n427_), .B0(new_new_n372_), .Y(new_new_n843_));
  NA2        g0821(.A(new_new_n843_), .B(new_new_n841_), .Y(new_new_n844_));
  AO220      g0822(.A0(new_new_n371_), .A1(new_new_n362_), .B0(new_new_n410_), .B1(new_new_n628_), .Y(new_new_n845_));
  NA3        g0823(.A(new_new_n845_), .B(new_new_n262_), .C(i_7_), .Y(new_new_n846_));
  BUFFER     g0824(.A(new_new_n653_), .Y(new_new_n847_));
  NA3        g0825(.A(new_new_n847_), .B(new_new_n147_), .C(new_new_n69_), .Y(new_new_n848_));
  AO210      g0826(.A0(new_new_n518_), .A1(new_new_n775_), .B0(new_new_n36_), .Y(new_new_n849_));
  NA4        g0827(.A(new_new_n849_), .B(new_new_n848_), .C(new_new_n846_), .D(new_new_n844_), .Y(new_new_n850_));
  OAI210     g0828(.A0(new_new_n667_), .A1(i_11_), .B0(new_new_n87_), .Y(new_new_n851_));
  AOI220     g0829(.A0(new_new_n851_), .A1(new_new_n595_), .B0(new_new_n816_), .B1(new_new_n740_), .Y(new_new_n852_));
  NA2        g0830(.A(new_new_n410_), .B(new_new_n70_), .Y(new_new_n853_));
  NA3        g0831(.A(new_new_n853_), .B(new_new_n852_), .C(new_new_n635_), .Y(new_new_n854_));
  AO210      g0832(.A0(new_new_n546_), .A1(new_new_n47_), .B0(new_new_n88_), .Y(new_new_n855_));
  NA3        g0833(.A(new_new_n855_), .B(new_new_n507_), .C(new_new_n221_), .Y(new_new_n856_));
  AOI210     g0834(.A0(new_new_n469_), .A1(new_new_n467_), .B0(new_new_n594_), .Y(new_new_n857_));
  NA2        g0835(.A(new_new_n113_), .B(new_new_n425_), .Y(new_new_n858_));
  NA2        g0836(.A(new_new_n249_), .B(new_new_n47_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n859_), .B(new_new_n617_), .Y(new_new_n860_));
  NA3        g0838(.A(new_new_n860_), .B(new_new_n337_), .C(i_7_), .Y(new_new_n861_));
  NA4        g0839(.A(new_new_n861_), .B(new_new_n858_), .C(new_new_n857_), .D(new_new_n856_), .Y(new_new_n862_));
  NO4        g0840(.A(new_new_n862_), .B(new_new_n854_), .C(new_new_n850_), .D(new_new_n840_), .Y(new_new_n863_));
  NA4        g0841(.A(new_new_n863_), .B(new_new_n825_), .C(new_new_n818_), .D(new_new_n392_), .Y(mai3));
  NA2        g0842(.A(i_12_), .B(i_10_), .Y(new_new_n865_));
  NA2        g0843(.A(i_6_), .B(i_7_), .Y(new_new_n866_));
  NO2        g0844(.A(new_new_n866_), .B(i_0_), .Y(new_new_n867_));
  NO2        g0845(.A(i_11_), .B(new_new_n241_), .Y(new_new_n868_));
  OAI210     g0846(.A0(new_new_n867_), .A1(new_new_n297_), .B0(new_new_n868_), .Y(new_new_n869_));
  NO2        g0847(.A(new_new_n869_), .B(new_new_n195_), .Y(new_new_n870_));
  NO3        g0848(.A(new_new_n473_), .B(new_new_n92_), .C(new_new_n45_), .Y(new_new_n871_));
  OA210      g0849(.A0(new_new_n871_), .A1(new_new_n870_), .B0(new_new_n175_), .Y(new_new_n872_));
  NA2        g0850(.A(new_new_n428_), .B(new_new_n46_), .Y(new_new_n873_));
  NO4        g0851(.A(new_new_n388_), .B(new_new_n395_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n187_), .B(new_new_n604_), .Y(new_new_n875_));
  NOi31      g0853(.An(new_new_n875_), .B(new_new_n874_), .C(new_new_n39_), .Y(new_new_n876_));
  NA2        g0854(.A(new_new_n733_), .B(new_new_n701_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n343_), .B(new_new_n458_), .Y(new_new_n878_));
  OAI220     g0856(.A0(new_new_n878_), .A1(new_new_n877_), .B0(new_new_n876_), .B1(new_new_n63_), .Y(new_new_n879_));
  NOi21      g0857(.An(i_5_), .B(i_9_), .Y(new_new_n880_));
  NA2        g0858(.A(new_new_n880_), .B(new_new_n466_), .Y(new_new_n881_));
  BUFFER     g0859(.A(new_new_n275_), .Y(new_new_n882_));
  NA2        g0860(.A(new_new_n882_), .B(new_new_n498_), .Y(new_new_n883_));
  NO3        g0861(.A(new_new_n431_), .B(new_new_n275_), .C(new_new_n73_), .Y(new_new_n884_));
  NO2        g0862(.A(new_new_n176_), .B(new_new_n148_), .Y(new_new_n885_));
  AOI210     g0863(.A0(new_new_n885_), .A1(new_new_n249_), .B0(new_new_n884_), .Y(new_new_n886_));
  OAI220     g0864(.A0(new_new_n886_), .A1(new_new_n182_), .B0(new_new_n883_), .B1(new_new_n881_), .Y(new_new_n887_));
  NO3        g0865(.A(new_new_n887_), .B(new_new_n879_), .C(new_new_n872_), .Y(new_new_n888_));
  NA2        g0866(.A(new_new_n187_), .B(new_new_n24_), .Y(new_new_n889_));
  NO2        g0867(.A(new_new_n699_), .B(new_new_n625_), .Y(new_new_n890_));
  NO2        g0868(.A(new_new_n890_), .B(new_new_n889_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n320_), .B(new_new_n129_), .Y(new_new_n892_));
  NAi21      g0870(.An(new_new_n162_), .B(new_new_n458_), .Y(new_new_n893_));
  OAI220     g0871(.A0(new_new_n893_), .A1(new_new_n859_), .B0(new_new_n892_), .B1(new_new_n416_), .Y(new_new_n894_));
  NO2        g0872(.A(new_new_n894_), .B(new_new_n891_), .Y(new_new_n895_));
  NO2        g0873(.A(new_new_n402_), .B(new_new_n301_), .Y(new_new_n896_));
  NA2        g0874(.A(new_new_n896_), .B(new_new_n736_), .Y(new_new_n897_));
  NA2        g0875(.A(new_new_n605_), .B(i_0_), .Y(new_new_n898_));
  NO3        g0876(.A(new_new_n898_), .B(new_new_n397_), .C(new_new_n89_), .Y(new_new_n899_));
  INV        g0877(.A(new_new_n899_), .Y(new_new_n900_));
  INV        g0878(.A(new_new_n496_), .Y(new_new_n901_));
  AN2        g0879(.A(new_new_n98_), .B(new_new_n248_), .Y(new_new_n902_));
  NA2        g0880(.A(new_new_n771_), .B(new_new_n338_), .Y(new_new_n903_));
  INV        g0881(.A(new_new_n58_), .Y(new_new_n904_));
  OAI220     g0882(.A0(new_new_n904_), .A1(new_new_n903_), .B0(new_new_n687_), .B1(new_new_n564_), .Y(new_new_n905_));
  NO2        g0883(.A(new_new_n259_), .B(new_new_n153_), .Y(new_new_n906_));
  NA2        g0884(.A(i_0_), .B(i_10_), .Y(new_new_n907_));
  AN2        g0885(.A(new_new_n906_), .B(i_6_), .Y(new_new_n908_));
  AOI220     g0886(.A0(new_new_n343_), .A1(new_new_n100_), .B0(new_new_n187_), .B1(new_new_n84_), .Y(new_new_n909_));
  NA2        g0887(.A(new_new_n599_), .B(i_4_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n190_), .B(new_new_n205_), .Y(new_new_n911_));
  OAI220     g0889(.A0(new_new_n911_), .A1(new_new_n903_), .B0(new_new_n910_), .B1(new_new_n909_), .Y(new_new_n912_));
  NO4        g0890(.A(new_new_n912_), .B(new_new_n908_), .C(new_new_n905_), .D(new_new_n902_), .Y(new_new_n913_));
  NA4        g0891(.A(new_new_n913_), .B(new_new_n900_), .C(new_new_n897_), .D(new_new_n895_), .Y(new_new_n914_));
  NA2        g0892(.A(i_11_), .B(i_9_), .Y(new_new_n915_));
  NO2        g0893(.A(new_new_n49_), .B(i_7_), .Y(new_new_n916_));
  NA2        g0894(.A(new_new_n407_), .B(new_new_n180_), .Y(new_new_n917_));
  NA2        g0895(.A(new_new_n917_), .B(new_new_n160_), .Y(new_new_n918_));
  NO2        g0896(.A(new_new_n915_), .B(new_new_n73_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n176_), .B(i_0_), .Y(new_new_n920_));
  INV        g0898(.A(new_new_n920_), .Y(new_new_n921_));
  NA2        g0899(.A(new_new_n496_), .B(new_new_n235_), .Y(new_new_n922_));
  AOI210     g0900(.A0(new_new_n382_), .A1(new_new_n42_), .B0(new_new_n424_), .Y(new_new_n923_));
  OAI220     g0901(.A0(new_new_n923_), .A1(new_new_n881_), .B0(new_new_n922_), .B1(new_new_n921_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n924_), .B(new_new_n918_), .Y(new_new_n925_));
  NA2        g0903(.A(new_new_n686_), .B(new_new_n121_), .Y(new_new_n926_));
  NO2        g0904(.A(i_6_), .B(new_new_n926_), .Y(new_new_n927_));
  AOI210     g0905(.A0(new_new_n468_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n928_));
  NA2        g0906(.A(new_new_n172_), .B(new_new_n105_), .Y(new_new_n929_));
  INV        g0907(.A(new_new_n927_), .Y(new_new_n930_));
  NOi21      g0908(.An(i_7_), .B(i_5_), .Y(new_new_n931_));
  NOi31      g0909(.An(new_new_n931_), .B(i_0_), .C(new_new_n750_), .Y(new_new_n932_));
  NA3        g0910(.A(new_new_n932_), .B(new_new_n396_), .C(i_6_), .Y(new_new_n933_));
  OA210      g0911(.A0(new_new_n929_), .A1(new_new_n544_), .B0(new_new_n933_), .Y(new_new_n934_));
  NO3        g0912(.A(new_new_n419_), .B(new_new_n374_), .C(new_new_n370_), .Y(new_new_n935_));
  NO2        g0913(.A(new_new_n269_), .B(new_new_n327_), .Y(new_new_n936_));
  NO2        g0914(.A(new_new_n750_), .B(new_new_n264_), .Y(new_new_n937_));
  AOI210     g0915(.A0(new_new_n937_), .A1(new_new_n936_), .B0(new_new_n935_), .Y(new_new_n938_));
  NA4        g0916(.A(new_new_n938_), .B(new_new_n934_), .C(new_new_n930_), .D(new_new_n925_), .Y(new_new_n939_));
  NO2        g0917(.A(new_new_n889_), .B(new_new_n244_), .Y(new_new_n940_));
  AN2        g0918(.A(new_new_n342_), .B(new_new_n338_), .Y(new_new_n941_));
  AO220      g0919(.A0(new_new_n941_), .A1(new_new_n885_), .B0(new_new_n357_), .B1(new_new_n27_), .Y(new_new_n942_));
  OAI210     g0920(.A0(new_new_n942_), .A1(new_new_n940_), .B0(i_10_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n865_), .B(new_new_n326_), .Y(new_new_n944_));
  NA2        g0922(.A(new_new_n944_), .B(new_new_n919_), .Y(new_new_n945_));
  NA3        g0923(.A(new_new_n495_), .B(new_new_n428_), .C(new_new_n46_), .Y(new_new_n946_));
  OAI210     g0924(.A0(new_new_n893_), .A1(new_new_n901_), .B0(new_new_n946_), .Y(new_new_n947_));
  NO2        g0925(.A(new_new_n262_), .B(new_new_n47_), .Y(new_new_n948_));
  NO2        g0926(.A(new_new_n948_), .B(new_new_n189_), .Y(new_new_n949_));
  AOI220     g0927(.A0(new_new_n949_), .A1(new_new_n496_), .B0(new_new_n947_), .B1(new_new_n73_), .Y(new_new_n950_));
  NA3        g0928(.A(new_new_n842_), .B(new_new_n394_), .C(new_new_n667_), .Y(new_new_n951_));
  NA2        g0929(.A(new_new_n95_), .B(new_new_n45_), .Y(new_new_n952_));
  NO2        g0930(.A(new_new_n75_), .B(new_new_n773_), .Y(new_new_n953_));
  AOI220     g0931(.A0(new_new_n953_), .A1(new_new_n952_), .B0(new_new_n175_), .B1(new_new_n625_), .Y(new_new_n954_));
  AOI210     g0932(.A0(new_new_n954_), .A1(new_new_n951_), .B0(new_new_n48_), .Y(new_new_n955_));
  NO3        g0933(.A(new_new_n616_), .B(new_new_n369_), .C(new_new_n24_), .Y(new_new_n956_));
  AOI210     g0934(.A0(new_new_n727_), .A1(new_new_n576_), .B0(new_new_n956_), .Y(new_new_n957_));
  NAi21      g0935(.An(i_9_), .B(i_5_), .Y(new_new_n958_));
  NO2        g0936(.A(new_new_n958_), .B(new_new_n419_), .Y(new_new_n959_));
  NA2        g0937(.A(new_new_n959_), .B(new_new_n653_), .Y(new_new_n960_));
  OAI220     g0938(.A0(new_new_n960_), .A1(new_new_n86_), .B0(new_new_n957_), .B1(new_new_n173_), .Y(new_new_n961_));
  NO3        g0939(.A(new_new_n961_), .B(new_new_n955_), .C(new_new_n548_), .Y(new_new_n962_));
  NA4        g0940(.A(new_new_n962_), .B(new_new_n950_), .C(new_new_n945_), .D(new_new_n943_), .Y(new_new_n963_));
  NO3        g0941(.A(new_new_n963_), .B(new_new_n939_), .C(new_new_n914_), .Y(new_new_n964_));
  NO2        g0942(.A(i_0_), .B(new_new_n750_), .Y(new_new_n965_));
  NA2        g0943(.A(new_new_n73_), .B(new_new_n45_), .Y(new_new_n966_));
  NA2        g0944(.A(new_new_n907_), .B(new_new_n966_), .Y(new_new_n967_));
  NO3        g0945(.A(new_new_n107_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n968_));
  AO220      g0946(.A0(new_new_n968_), .A1(new_new_n967_), .B0(new_new_n965_), .B1(new_new_n175_), .Y(new_new_n969_));
  NO2        g0947(.A(new_new_n820_), .B(new_new_n929_), .Y(new_new_n970_));
  AOI210     g0948(.A0(new_new_n969_), .A1(new_new_n359_), .B0(new_new_n970_), .Y(new_new_n971_));
  NA2        g0949(.A(new_new_n760_), .B(new_new_n146_), .Y(new_new_n972_));
  INV        g0950(.A(new_new_n972_), .Y(new_new_n973_));
  NA3        g0951(.A(new_new_n973_), .B(new_new_n701_), .C(new_new_n73_), .Y(new_new_n974_));
  NO2        g0952(.A(new_new_n838_), .B(new_new_n419_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n867_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n868_), .B(i_9_), .Y(new_new_n977_));
  AOI210     g0955(.A0(new_new_n976_), .A1(new_new_n523_), .B0(new_new_n977_), .Y(new_new_n978_));
  OAI210     g0956(.A0(new_new_n249_), .A1(i_9_), .B0(new_new_n234_), .Y(new_new_n979_));
  AOI210     g0957(.A0(new_new_n979_), .A1(new_new_n898_), .B0(new_new_n153_), .Y(new_new_n980_));
  NO3        g0958(.A(new_new_n980_), .B(new_new_n978_), .C(new_new_n975_), .Y(new_new_n981_));
  NA3        g0959(.A(new_new_n981_), .B(new_new_n974_), .C(new_new_n971_), .Y(new_new_n982_));
  NA2        g0960(.A(new_new_n941_), .B(new_new_n384_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n308_), .A1(new_new_n162_), .B0(new_new_n983_), .Y(new_new_n984_));
  NA3        g0962(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n916_), .B(new_new_n512_), .Y(new_new_n986_));
  AOI210     g0964(.A0(new_new_n985_), .A1(new_new_n162_), .B0(new_new_n986_), .Y(new_new_n987_));
  NO2        g0965(.A(new_new_n987_), .B(new_new_n984_), .Y(new_new_n988_));
  NO3        g0966(.A(new_new_n907_), .B(new_new_n880_), .C(new_new_n192_), .Y(new_new_n989_));
  AOI220     g0967(.A0(new_new_n989_), .A1(i_11_), .B0(new_new_n600_), .B1(new_new_n75_), .Y(new_new_n990_));
  NO3        g0968(.A(new_new_n212_), .B(new_new_n395_), .C(i_0_), .Y(new_new_n991_));
  OAI210     g0969(.A0(new_new_n991_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n992_));
  INV        g0970(.A(new_new_n221_), .Y(new_new_n993_));
  OAI220     g0971(.A0(new_new_n558_), .A1(new_new_n139_), .B0(new_new_n672_), .B1(new_new_n647_), .Y(new_new_n994_));
  NA3        g0972(.A(new_new_n994_), .B(new_new_n411_), .C(new_new_n993_), .Y(new_new_n995_));
  NA4        g0973(.A(new_new_n995_), .B(new_new_n992_), .C(new_new_n990_), .D(new_new_n988_), .Y(new_new_n996_));
  AOI220     g0974(.A0(new_new_n931_), .A1(new_new_n512_), .B0(new_new_n867_), .B1(new_new_n163_), .Y(new_new_n997_));
  NA2        g0975(.A(new_new_n362_), .B(new_new_n177_), .Y(new_new_n998_));
  OR2        g0976(.A(new_new_n998_), .B(new_new_n997_), .Y(new_new_n999_));
  AOI210     g0977(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n176_), .Y(new_new_n1000_));
  NA3        g0978(.A(new_new_n644_), .B(new_new_n187_), .C(new_new_n84_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n1001_), .B(new_new_n574_), .Y(new_new_n1002_));
  NO3        g0980(.A(new_new_n873_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n1003_));
  NA3        g0981(.A(new_new_n517_), .B(new_new_n510_), .C(new_new_n493_), .Y(new_new_n1004_));
  NO3        g0982(.A(new_new_n1004_), .B(new_new_n1003_), .C(new_new_n1002_), .Y(new_new_n1005_));
  NA3        g0983(.A(new_new_n916_), .B(new_new_n297_), .C(new_new_n234_), .Y(new_new_n1006_));
  INV        g0984(.A(new_new_n1006_), .Y(new_new_n1007_));
  NA3        g0985(.A(new_new_n402_), .B(new_new_n344_), .C(new_new_n225_), .Y(new_new_n1008_));
  OAI210     g0986(.A0(new_new_n875_), .A1(new_new_n675_), .B0(new_new_n1008_), .Y(new_new_n1009_));
  NOi31      g0987(.An(new_new_n401_), .B(new_new_n966_), .C(new_new_n244_), .Y(new_new_n1010_));
  NO3        g0988(.A(new_new_n915_), .B(new_new_n221_), .C(new_new_n192_), .Y(new_new_n1011_));
  NO4        g0989(.A(new_new_n1011_), .B(new_new_n1010_), .C(new_new_n1009_), .D(new_new_n1007_), .Y(new_new_n1012_));
  NA3        g0990(.A(new_new_n1012_), .B(new_new_n1005_), .C(new_new_n999_), .Y(new_new_n1013_));
  INV        g0991(.A(new_new_n646_), .Y(new_new_n1014_));
  NO3        g0992(.A(new_new_n1014_), .B(new_new_n590_), .C(new_new_n356_), .Y(new_new_n1015_));
  NO2        g0993(.A(new_new_n86_), .B(i_5_), .Y(new_new_n1016_));
  NA3        g0994(.A(new_new_n868_), .B(new_new_n111_), .C(new_new_n124_), .Y(new_new_n1017_));
  INV        g0995(.A(new_new_n1017_), .Y(new_new_n1018_));
  AOI210     g0996(.A0(new_new_n1018_), .A1(new_new_n1016_), .B0(new_new_n1015_), .Y(new_new_n1019_));
  NA3        g0997(.A(new_new_n313_), .B(i_5_), .C(new_new_n195_), .Y(new_new_n1020_));
  NA2        g0998(.A(new_new_n1020_), .B(new_new_n247_), .Y(new_new_n1021_));
  NO4        g0999(.A(new_new_n244_), .B(new_new_n212_), .C(i_0_), .D(i_12_), .Y(new_new_n1022_));
  NA2        g1000(.A(new_new_n1022_), .B(new_new_n1021_), .Y(new_new_n1023_));
  AN2        g1001(.A(new_new_n907_), .B(new_new_n153_), .Y(new_new_n1024_));
  NO4        g1002(.A(new_new_n1024_), .B(i_12_), .C(new_new_n675_), .D(new_new_n131_), .Y(new_new_n1025_));
  NA2        g1003(.A(new_new_n1025_), .B(new_new_n221_), .Y(new_new_n1026_));
  NA3        g1004(.A(new_new_n100_), .B(new_new_n604_), .C(i_11_), .Y(new_new_n1027_));
  NO2        g1005(.A(new_new_n1027_), .B(new_new_n155_), .Y(new_new_n1028_));
  NA2        g1006(.A(new_new_n931_), .B(new_new_n492_), .Y(new_new_n1029_));
  NA2        g1007(.A(new_new_n64_), .B(new_new_n103_), .Y(new_new_n1030_));
  OAI220     g1008(.A0(new_new_n1030_), .A1(new_new_n1020_), .B0(new_new_n1029_), .B1(new_new_n702_), .Y(new_new_n1031_));
  AOI210     g1009(.A0(new_new_n1031_), .A1(new_new_n920_), .B0(new_new_n1028_), .Y(new_new_n1032_));
  NA4        g1010(.A(new_new_n1032_), .B(new_new_n1026_), .C(new_new_n1023_), .D(new_new_n1019_), .Y(new_new_n1033_));
  NO4        g1011(.A(new_new_n1033_), .B(new_new_n1013_), .C(new_new_n996_), .D(new_new_n982_), .Y(new_new_n1034_));
  OAI210     g1012(.A0(new_new_n841_), .A1(new_new_n834_), .B0(new_new_n37_), .Y(new_new_n1035_));
  NA3        g1013(.A(new_new_n928_), .B(new_new_n379_), .C(i_5_), .Y(new_new_n1036_));
  NA3        g1014(.A(new_new_n1036_), .B(new_new_n1035_), .C(new_new_n642_), .Y(new_new_n1037_));
  NA2        g1015(.A(new_new_n1037_), .B(new_new_n209_), .Y(new_new_n1038_));
  BUFFER     g1016(.A(new_new_n380_), .Y(new_new_n1039_));
  NA2        g1017(.A(new_new_n188_), .B(new_new_n190_), .Y(new_new_n1040_));
  AO210      g1018(.A0(new_new_n1039_), .A1(new_new_n33_), .B0(new_new_n1040_), .Y(new_new_n1041_));
  OAI210     g1019(.A0(new_new_n646_), .A1(new_new_n644_), .B0(new_new_n326_), .Y(new_new_n1042_));
  NA2        g1020(.A(new_new_n1042_), .B(new_new_n1041_), .Y(new_new_n1043_));
  NO4        g1021(.A(new_new_n237_), .B(new_new_n145_), .C(new_new_n705_), .D(new_new_n37_), .Y(new_new_n1044_));
  INV        g1022(.A(new_new_n1044_), .Y(new_new_n1045_));
  OAI210     g1023(.A0(new_new_n1027_), .A1(new_new_n148_), .B0(new_new_n1045_), .Y(new_new_n1046_));
  AOI210     g1024(.A0(new_new_n1043_), .A1(new_new_n49_), .B0(new_new_n1046_), .Y(new_new_n1047_));
  AOI210     g1025(.A0(new_new_n1047_), .A1(new_new_n1038_), .B0(new_new_n73_), .Y(new_new_n1048_));
  NO2        g1026(.A(new_new_n597_), .B(new_new_n391_), .Y(new_new_n1049_));
  NO2        g1027(.A(new_new_n1049_), .B(new_new_n779_), .Y(new_new_n1050_));
  OAI210     g1028(.A0(new_new_n80_), .A1(new_new_n55_), .B0(new_new_n110_), .Y(new_new_n1051_));
  NA2        g1029(.A(new_new_n1051_), .B(new_new_n76_), .Y(new_new_n1052_));
  AOI210     g1030(.A0(new_new_n1000_), .A1(new_new_n916_), .B0(new_new_n932_), .Y(new_new_n1053_));
  AOI210     g1031(.A0(new_new_n1053_), .A1(new_new_n1052_), .B0(new_new_n705_), .Y(new_new_n1054_));
  NA2        g1032(.A(new_new_n269_), .B(new_new_n57_), .Y(new_new_n1055_));
  AOI220     g1033(.A0(new_new_n1055_), .A1(new_new_n76_), .B0(new_new_n357_), .B1(new_new_n261_), .Y(new_new_n1056_));
  NO2        g1034(.A(new_new_n1056_), .B(new_new_n241_), .Y(new_new_n1057_));
  NA3        g1035(.A(new_new_n98_), .B(new_new_n315_), .C(new_new_n31_), .Y(new_new_n1058_));
  INV        g1036(.A(new_new_n1058_), .Y(new_new_n1059_));
  NO3        g1037(.A(new_new_n1059_), .B(new_new_n1057_), .C(new_new_n1054_), .Y(new_new_n1060_));
  NA2        g1038(.A(new_new_n158_), .B(new_new_n89_), .Y(new_new_n1061_));
  NA3        g1039(.A(new_new_n783_), .B(new_new_n297_), .C(new_new_n80_), .Y(new_new_n1062_));
  AOI210     g1040(.A0(new_new_n1062_), .A1(new_new_n1061_), .B0(i_11_), .Y(new_new_n1063_));
  NA2        g1041(.A(new_new_n637_), .B(new_new_n218_), .Y(new_new_n1064_));
  OAI210     g1042(.A0(new_new_n1064_), .A1(new_new_n928_), .B0(new_new_n209_), .Y(new_new_n1065_));
  NA2        g1043(.A(new_new_n164_), .B(i_5_), .Y(new_new_n1066_));
  NO2        g1044(.A(new_new_n1065_), .B(new_new_n1066_), .Y(new_new_n1067_));
  NO4        g1045(.A(new_new_n958_), .B(new_new_n500_), .C(new_new_n258_), .D(new_new_n257_), .Y(new_new_n1068_));
  NO2        g1046(.A(new_new_n1068_), .B(new_new_n594_), .Y(new_new_n1069_));
  NO2        g1047(.A(new_new_n837_), .B(new_new_n375_), .Y(new_new_n1070_));
  AOI210     g1048(.A0(new_new_n1070_), .A1(new_new_n1069_), .B0(new_new_n41_), .Y(new_new_n1071_));
  NO3        g1049(.A(new_new_n1071_), .B(new_new_n1067_), .C(new_new_n1063_), .Y(new_new_n1072_));
  OAI210     g1050(.A0(new_new_n1060_), .A1(i_4_), .B0(new_new_n1072_), .Y(new_new_n1073_));
  NO3        g1051(.A(new_new_n1073_), .B(new_new_n1050_), .C(new_new_n1048_), .Y(new_new_n1074_));
  NA4        g1052(.A(new_new_n1074_), .B(new_new_n1034_), .C(new_new_n964_), .D(new_new_n888_), .Y(mai4));
  INV        g1053(.A(i_2_), .Y(new_new_n1078_));
  INV        g1054(.A(new_new_n338_), .Y(new_new_n1079_));
  INV        g1055(.A(new_new_n507_), .Y(new_new_n1080_));
endmodule


