//Benchmark atmr_misex3_1774_0.125

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n396_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o000(.A(j), .B(g), .Y(ori_ori_n29_));
  INV        o001(.A(i), .Y(ori_ori_n30_));
  AN2        o002(.A(h), .B(g), .Y(ori_ori_n31_));
  NAi21      o003(.An(n), .B(m), .Y(ori_ori_n32_));
  NOi32      o004(.An(k), .Bn(h), .C(l), .Y(ori_ori_n33_));
  INV        o005(.A(c), .Y(ori_ori_n34_));
  INV        o006(.A(d), .Y(ori_ori_n35_));
  NAi21      o007(.An(i), .B(h), .Y(ori_ori_n36_));
  INV        o008(.A(f), .Y(ori_ori_n37_));
  INV        o009(.A(m), .Y(ori_ori_n38_));
  INV        o010(.A(n), .Y(ori_ori_n39_));
  INV        o011(.A(j), .Y(ori_ori_n40_));
  NAi41      o012(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n41_));
  NOi21      o013(.An(i), .B(h), .Y(ori_ori_n42_));
  NOi21      o014(.An(m), .B(n), .Y(ori_ori_n43_));
  AN2        o015(.A(k), .B(h), .Y(ori_ori_n44_));
  INV        o016(.A(b), .Y(ori_ori_n45_));
  AN2        o017(.A(k), .B(i), .Y(ori_ori_n46_));
  NOi32      o018(.An(f), .Bn(b), .C(e), .Y(ori_ori_n47_));
  NAi21      o019(.An(m), .B(n), .Y(ori_ori_n48_));
  NAi31      o020(.An(j), .B(k), .C(h), .Y(ori_ori_n49_));
  NAi21      o021(.An(e), .B(f), .Y(ori_ori_n50_));
  NAi21      o022(.An(c), .B(d), .Y(ori_ori_n51_));
  NOi21      o023(.An(h), .B(i), .Y(ori_ori_n52_));
  NOi21      o024(.An(k), .B(m), .Y(ori_ori_n53_));
  NA3        o025(.A(ori_ori_n53_), .B(ori_ori_n52_), .C(n), .Y(ori_ori_n54_));
  NAi31      o026(.An(d), .B(f), .C(c), .Y(ori_ori_n55_));
  NAi31      o027(.An(e), .B(f), .C(c), .Y(ori_ori_n56_));
  NA2        o028(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  NA2        o029(.A(j), .B(h), .Y(ori_ori_n58_));
  OR3        o030(.A(n), .B(m), .C(k), .Y(ori_ori_n59_));
  NO2        o031(.A(ori_ori_n59_), .B(ori_ori_n58_), .Y(ori_ori_n60_));
  NAi32      o032(.An(m), .Bn(k), .C(n), .Y(ori_ori_n61_));
  NA2        o033(.A(ori_ori_n60_), .B(ori_ori_n57_), .Y(ori_ori_n62_));
  NO2        o034(.A(n), .B(m), .Y(ori_ori_n63_));
  NA2        o035(.A(ori_ori_n63_), .B(ori_ori_n33_), .Y(ori_ori_n64_));
  NAi21      o036(.An(f), .B(e), .Y(ori_ori_n65_));
  NA2        o037(.A(d), .B(c), .Y(ori_ori_n66_));
  NAi21      o038(.An(h), .B(f), .Y(ori_ori_n67_));
  NOi32      o039(.An(f), .Bn(c), .C(d), .Y(ori_ori_n68_));
  NOi32      o040(.An(f), .Bn(c), .C(e), .Y(ori_ori_n69_));
  NO2        o041(.A(ori_ori_n69_), .B(ori_ori_n68_), .Y(ori_ori_n70_));
  NO3        o042(.A(n), .B(m), .C(j), .Y(ori_ori_n71_));
  NA2        o043(.A(ori_ori_n71_), .B(ori_ori_n44_), .Y(ori_ori_n72_));
  AO210      o044(.A0(ori_ori_n72_), .A1(ori_ori_n64_), .B0(ori_ori_n70_), .Y(ori_ori_n73_));
  NA2        o045(.A(ori_ori_n73_), .B(ori_ori_n62_), .Y(ori_ori_n74_));
  INV        o046(.A(ori_ori_n74_), .Y(ori_ori_n75_));
  NAi31      o047(.An(n), .B(h), .C(g), .Y(ori_ori_n76_));
  INV        o048(.A(f), .Y(ori_ori_n77_));
  INV        o049(.A(g), .Y(ori_ori_n78_));
  NOi31      o050(.An(i), .B(j), .C(h), .Y(ori_ori_n79_));
  NOi21      o051(.An(l), .B(m), .Y(ori_ori_n80_));
  NOi21      o052(.An(n), .B(m), .Y(ori_ori_n81_));
  NAi21      o053(.An(j), .B(h), .Y(ori_ori_n82_));
  XN2        o054(.A(i), .B(h), .Y(ori_ori_n83_));
  NA2        o055(.A(ori_ori_n83_), .B(ori_ori_n82_), .Y(ori_ori_n84_));
  NOi31      o056(.An(k), .B(n), .C(m), .Y(ori_ori_n85_));
  NOi31      o057(.An(ori_ori_n85_), .B(ori_ori_n66_), .C(ori_ori_n65_), .Y(ori_ori_n86_));
  NA2        o058(.A(ori_ori_n86_), .B(ori_ori_n84_), .Y(ori_ori_n87_));
  NAi31      o059(.An(f), .B(e), .C(c), .Y(ori_ori_n88_));
  NO4        o060(.A(ori_ori_n88_), .B(ori_ori_n59_), .C(ori_ori_n58_), .D(ori_ori_n35_), .Y(ori_ori_n89_));
  NAi32      o061(.An(m), .Bn(i), .C(k), .Y(ori_ori_n90_));
  INV        o062(.A(k), .Y(ori_ori_n91_));
  INV        o063(.A(ori_ori_n89_), .Y(ori_ori_n92_));
  AN2        o064(.A(ori_ori_n92_), .B(ori_ori_n87_), .Y(ori_ori_n93_));
  BUFFER     o065(.A(g), .Y(ori_ori_n94_));
  NO2        o066(.A(ori_ori_n94_), .B(ori_ori_n41_), .Y(ori_ori_n95_));
  NA2        o067(.A(ori_ori_n95_), .B(ori_ori_n47_), .Y(ori_ori_n96_));
  NA2        o068(.A(ori_ori_n53_), .B(ori_ori_n42_), .Y(ori_ori_n97_));
  NAi21      o069(.An(h), .B(i), .Y(ori_ori_n98_));
  NA2        o070(.A(ori_ori_n63_), .B(k), .Y(ori_ori_n99_));
  NO2        o071(.A(ori_ori_n99_), .B(ori_ori_n98_), .Y(ori_ori_n100_));
  NA2        o072(.A(ori_ori_n100_), .B(ori_ori_n68_), .Y(ori_ori_n101_));
  NA2        o073(.A(ori_ori_n101_), .B(ori_ori_n96_), .Y(ori_ori_n102_));
  NOi21      o074(.An(ori_ori_n93_), .B(ori_ori_n102_), .Y(ori_ori_n103_));
  INV        o075(.A(c), .Y(ori_ori_n104_));
  NA3        o076(.A(ori_ori_n53_), .B(ori_ori_n52_), .C(ori_ori_n39_), .Y(ori_ori_n105_));
  NO2        o077(.A(ori_ori_n105_), .B(ori_ori_n70_), .Y(ori_ori_n106_));
  NA3        o078(.A(e), .B(c), .C(b), .Y(ori_ori_n107_));
  NAi32      o079(.An(j), .Bn(h), .C(i), .Y(ori_ori_n108_));
  NAi21      o080(.An(m), .B(l), .Y(ori_ori_n109_));
  NAi32      o081(.An(n), .Bn(m), .C(l), .Y(ori_ori_n110_));
  NO2        o082(.A(ori_ori_n110_), .B(ori_ori_n108_), .Y(ori_ori_n111_));
  INV        o083(.A(ori_ori_n106_), .Y(ori_ori_n112_));
  NA2        o084(.A(ori_ori_n100_), .B(ori_ori_n69_), .Y(ori_ori_n113_));
  NAi21      o085(.An(m), .B(k), .Y(ori_ori_n114_));
  NA2        o086(.A(e), .B(c), .Y(ori_ori_n115_));
  NO3        o087(.A(ori_ori_n115_), .B(n), .C(d), .Y(ori_ori_n116_));
  INV        o088(.A(ori_ori_n113_), .Y(ori_ori_n117_));
  NOi31      o089(.An(l), .B(n), .C(m), .Y(ori_ori_n118_));
  NA2        o090(.A(ori_ori_n118_), .B(ori_ori_n79_), .Y(ori_ori_n119_));
  NO2        o091(.A(ori_ori_n119_), .B(ori_ori_n70_), .Y(ori_ori_n120_));
  NAi32      o092(.An(m), .Bn(j), .C(k), .Y(ori_ori_n121_));
  NO2        o093(.A(ori_ori_n120_), .B(ori_ori_n117_), .Y(ori_ori_n122_));
  NA4        o094(.A(ori_ori_n122_), .B(ori_ori_n112_), .C(ori_ori_n103_), .D(ori_ori_n75_), .Y(ori10));
  NAi31      o095(.An(b), .B(f), .C(c), .Y(ori_ori_n124_));
  INV        o096(.A(ori_ori_n124_), .Y(ori_ori_n125_));
  NOi32      o097(.An(k), .Bn(h), .C(j), .Y(ori_ori_n126_));
  NA2        o098(.A(ori_ori_n126_), .B(ori_ori_n81_), .Y(ori_ori_n127_));
  NA2        o099(.A(ori_ori_n54_), .B(ori_ori_n127_), .Y(ori_ori_n128_));
  NA2        o100(.A(ori_ori_n128_), .B(ori_ori_n125_), .Y(ori_ori_n129_));
  AN2        o101(.A(j), .B(h), .Y(ori_ori_n130_));
  NO3        o102(.A(n), .B(m), .C(k), .Y(ori_ori_n131_));
  NA2        o103(.A(ori_ori_n131_), .B(ori_ori_n130_), .Y(ori_ori_n132_));
  NO3        o104(.A(ori_ori_n132_), .B(ori_ori_n51_), .C(ori_ori_n77_), .Y(ori_ori_n133_));
  OR2        o105(.A(m), .B(k), .Y(ori_ori_n134_));
  NO2        o106(.A(ori_ori_n58_), .B(ori_ori_n134_), .Y(ori_ori_n135_));
  NA4        o107(.A(n), .B(f), .C(c), .D(ori_ori_n45_), .Y(ori_ori_n136_));
  NOi21      o108(.An(ori_ori_n135_), .B(ori_ori_n136_), .Y(ori_ori_n137_));
  NO2        o109(.A(ori_ori_n137_), .B(ori_ori_n133_), .Y(ori_ori_n138_));
  NO2        o110(.A(ori_ori_n136_), .B(ori_ori_n109_), .Y(ori_ori_n139_));
  NOi32      o111(.An(f), .Bn(d), .C(c), .Y(ori_ori_n140_));
  NA2        o112(.A(ori_ori_n140_), .B(ori_ori_n111_), .Y(ori_ori_n141_));
  NA3        o113(.A(ori_ori_n141_), .B(ori_ori_n138_), .C(ori_ori_n129_), .Y(ori_ori_n142_));
  INV        o114(.A(e), .Y(ori_ori_n143_));
  INV        o115(.A(ori_ori_n142_), .Y(ori_ori_n144_));
  OR2        o116(.A(n), .B(m), .Y(ori_ori_n145_));
  NO2        o117(.A(ori_ori_n66_), .B(ori_ori_n50_), .Y(ori_ori_n146_));
  NA2        o118(.A(ori_ori_n60_), .B(ori_ori_n146_), .Y(ori_ori_n147_));
  NAi21      o119(.An(k), .B(j), .Y(ori_ori_n148_));
  NAi21      o120(.An(e), .B(d), .Y(ori_ori_n149_));
  INV        o121(.A(ori_ori_n149_), .Y(ori_ori_n150_));
  NO2        o122(.A(ori_ori_n99_), .B(ori_ori_n77_), .Y(ori_ori_n151_));
  NA3        o123(.A(ori_ori_n151_), .B(ori_ori_n150_), .C(ori_ori_n84_), .Y(ori_ori_n152_));
  NA2        o124(.A(ori_ori_n152_), .B(ori_ori_n147_), .Y(ori_ori_n153_));
  NO2        o125(.A(ori_ori_n119_), .B(ori_ori_n77_), .Y(ori_ori_n154_));
  NOi31      o126(.An(n), .B(m), .C(k), .Y(ori_ori_n155_));
  AOI220     o127(.A0(ori_ori_n155_), .A1(ori_ori_n130_), .B0(ori_ori_n81_), .B1(ori_ori_n33_), .Y(ori_ori_n156_));
  NAi31      o128(.An(g), .B(f), .C(c), .Y(ori_ori_n157_));
  INV        o129(.A(ori_ori_n153_), .Y(ori_ori_n158_));
  AN2        o130(.A(e), .B(d), .Y(ori_ori_n159_));
  NO2        o131(.A(ori_ori_n37_), .B(e), .Y(ori_ori_n160_));
  NO4        o132(.A(ori_ori_n67_), .B(ori_ori_n41_), .C(ori_ori_n34_), .D(b), .Y(ori_ori_n161_));
  AOI210     o133(.A0(ori_ori_n90_), .A1(ori_ori_n121_), .B0(ori_ori_n39_), .Y(ori_ori_n162_));
  INV        o134(.A(ori_ori_n161_), .Y(ori_ori_n163_));
  INV        o135(.A(ori_ori_n93_), .Y(ori_ori_n164_));
  XO2        o136(.A(i), .B(h), .Y(ori_ori_n165_));
  NA3        o137(.A(ori_ori_n165_), .B(ori_ori_n53_), .C(n), .Y(ori_ori_n166_));
  NA3        o138(.A(ori_ori_n166_), .B(ori_ori_n156_), .C(ori_ori_n127_), .Y(ori_ori_n167_));
  NOi32      o139(.An(ori_ori_n167_), .Bn(ori_ori_n160_), .C(ori_ori_n104_), .Y(ori_ori_n168_));
  NAi31      o140(.An(c), .B(f), .C(d), .Y(ori_ori_n169_));
  AOI210     o141(.A0(ori_ori_n105_), .A1(ori_ori_n72_), .B0(ori_ori_n169_), .Y(ori_ori_n170_));
  INV        o142(.A(ori_ori_n170_), .Y(ori_ori_n171_));
  NA2        o143(.A(ori_ori_n85_), .B(ori_ori_n42_), .Y(ori_ori_n172_));
  AOI210     o144(.A0(ori_ori_n172_), .A1(ori_ori_n64_), .B0(ori_ori_n169_), .Y(ori_ori_n173_));
  INV        o145(.A(ori_ori_n173_), .Y(ori_ori_n174_));
  NA2        o146(.A(ori_ori_n174_), .B(ori_ori_n171_), .Y(ori_ori_n175_));
  NO3        o147(.A(ori_ori_n175_), .B(ori_ori_n168_), .C(ori_ori_n164_), .Y(ori_ori_n176_));
  NA4        o148(.A(ori_ori_n176_), .B(ori_ori_n163_), .C(ori_ori_n158_), .D(ori_ori_n144_), .Y(ori11));
  INV        o149(.A(j), .Y(ori_ori_n178_));
  NAi32      o150(.An(e), .Bn(b), .C(c), .Y(ori_ori_n179_));
  INV        o151(.A(k), .Y(ori_ori_n180_));
  NO3        o152(.A(ori_ori_n114_), .B(ori_ori_n36_), .C(n), .Y(ori_ori_n181_));
  NA3        o153(.A(ori_ori_n169_), .B(ori_ori_n56_), .C(ori_ori_n55_), .Y(ori_ori_n182_));
  NA2        o154(.A(ori_ori_n157_), .B(ori_ori_n88_), .Y(ori_ori_n183_));
  OR2        o155(.A(ori_ori_n183_), .B(ori_ori_n182_), .Y(ori_ori_n184_));
  NA2        o156(.A(ori_ori_n184_), .B(ori_ori_n181_), .Y(ori_ori_n185_));
  NO2        o157(.A(ori_ori_n185_), .B(ori_ori_n40_), .Y(ori_ori_n186_));
  NOi32      o158(.An(e), .Bn(c), .C(f), .Y(ori_ori_n187_));
  NA2        o159(.A(ori_ori_n187_), .B(ori_ori_n60_), .Y(ori_ori_n188_));
  NA2        o160(.A(ori_ori_n188_), .B(ori_ori_n62_), .Y(ori_ori_n189_));
  NOi31      o161(.An(m), .B(n), .C(k), .Y(ori_ori_n190_));
  NA2        o162(.A(ori_ori_n165_), .B(ori_ori_n53_), .Y(ori_ori_n191_));
  NO3        o163(.A(ori_ori_n136_), .B(ori_ori_n191_), .C(ori_ori_n40_), .Y(ori_ori_n192_));
  INV        o164(.A(ori_ori_n192_), .Y(ori_ori_n193_));
  AN3        o165(.A(f), .B(d), .C(b), .Y(ori_ori_n194_));
  OAI210     o166(.A0(ori_ori_n194_), .A1(ori_ori_n47_), .B0(n), .Y(ori_ori_n195_));
  NA3        o167(.A(ori_ori_n165_), .B(ori_ori_n53_), .C(ori_ori_n78_), .Y(ori_ori_n196_));
  NO2        o168(.A(ori_ori_n195_), .B(ori_ori_n196_), .Y(ori_ori_n197_));
  NA2        o169(.A(ori_ori_n197_), .B(j), .Y(ori_ori_n198_));
  NA2        o170(.A(ori_ori_n198_), .B(ori_ori_n193_), .Y(ori_ori_n199_));
  NO3        o171(.A(ori_ori_n199_), .B(ori_ori_n189_), .C(ori_ori_n186_), .Y(ori_ori_n200_));
  NO3        o172(.A(g), .B(ori_ori_n77_), .C(ori_ori_n34_), .Y(ori_ori_n201_));
  NO2        o173(.A(ori_ori_n172_), .B(ori_ori_n40_), .Y(ori_ori_n202_));
  OAI210     o174(.A0(ori_ori_n202_), .A1(ori_ori_n135_), .B0(ori_ori_n201_), .Y(ori_ori_n203_));
  BUFFER     o175(.A(h), .Y(ori_ori_n204_));
  NA2        o176(.A(ori_ori_n204_), .B(ori_ori_n29_), .Y(ori_ori_n205_));
  INV        o177(.A(ori_ori_n203_), .Y(ori_ori_n206_));
  INV        o178(.A(ori_ori_n48_), .Y(ori_ori_n207_));
  NO3        o179(.A(ori_ori_n140_), .B(ori_ori_n69_), .C(ori_ori_n68_), .Y(ori_ori_n208_));
  NA2        o180(.A(ori_ori_n208_), .B(ori_ori_n88_), .Y(ori_ori_n209_));
  NA3        o181(.A(ori_ori_n209_), .B(ori_ori_n100_), .C(j), .Y(ori_ori_n210_));
  NA2        o182(.A(ori_ori_n210_), .B(ori_ori_n138_), .Y(ori_ori_n211_));
  NO2        o183(.A(ori_ori_n211_), .B(ori_ori_n206_), .Y(ori_ori_n212_));
  NA2        o184(.A(ori_ori_n212_), .B(ori_ori_n200_), .Y(ori08));
  NO2        o185(.A(k), .B(h), .Y(ori_ori_n214_));
  AO210      o186(.A0(ori_ori_n98_), .A1(ori_ori_n148_), .B0(ori_ori_n214_), .Y(ori_ori_n215_));
  NO2        o187(.A(ori_ori_n215_), .B(ori_ori_n109_), .Y(ori_ori_n216_));
  NA2        o188(.A(ori_ori_n187_), .B(ori_ori_n39_), .Y(ori_ori_n217_));
  NA2        o189(.A(ori_ori_n217_), .B(ori_ori_n157_), .Y(ori_ori_n218_));
  NA2        o190(.A(ori_ori_n218_), .B(ori_ori_n216_), .Y(ori_ori_n219_));
  NA4        o191(.A(ori_ori_n80_), .B(k), .C(ori_ori_n30_), .D(h), .Y(ori_ori_n220_));
  INV        o192(.A(ori_ori_n219_), .Y(ori_ori_n221_));
  NA2        o193(.A(ori_ori_n215_), .B(ori_ori_n49_), .Y(ori_ori_n222_));
  NA2        o194(.A(ori_ori_n222_), .B(ori_ori_n139_), .Y(ori_ori_n223_));
  INV        o195(.A(ori_ori_n223_), .Y(ori_ori_n224_));
  NA3        o196(.A(ori_ori_n209_), .B(ori_ori_n118_), .C(ori_ori_n126_), .Y(ori_ori_n225_));
  INV        o197(.A(ori_ori_n225_), .Y(ori_ori_n226_));
  NO3        o198(.A(ori_ori_n226_), .B(ori_ori_n224_), .C(ori_ori_n221_), .Y(ori_ori_n227_));
  NA2        o199(.A(l), .B(ori_ori_n38_), .Y(ori_ori_n228_));
  NO4        o200(.A(ori_ori_n208_), .B(ori_ori_n58_), .C(n), .D(i), .Y(ori_ori_n229_));
  BUFFER     o201(.A(h), .Y(ori_ori_n230_));
  INV        o202(.A(ori_ori_n229_), .Y(ori_ori_n231_));
  NO2        o203(.A(ori_ori_n231_), .B(ori_ori_n228_), .Y(ori_ori_n232_));
  INV        o204(.A(ori_ori_n232_), .Y(ori_ori_n233_));
  NO2        o205(.A(ori_ori_n109_), .B(ori_ori_n49_), .Y(ori_ori_n234_));
  NO2        o206(.A(ori_ori_n220_), .B(ori_ori_n217_), .Y(ori_ori_n235_));
  NO2        o207(.A(ori_ori_n120_), .B(ori_ori_n235_), .Y(ori_ori_n236_));
  INV        o208(.A(ori_ori_n141_), .Y(ori_ori_n237_));
  NO2        o209(.A(ori_ori_n220_), .B(ori_ori_n136_), .Y(ori_ori_n238_));
  NO2        o210(.A(ori_ori_n208_), .B(n), .Y(ori_ori_n239_));
  BUFFER     o211(.A(ori_ori_n234_), .Y(ori_ori_n240_));
  AOI220     o212(.A0(ori_ori_n240_), .A1(ori_ori_n201_), .B0(ori_ori_n239_), .B1(ori_ori_n216_), .Y(ori_ori_n241_));
  INV        o213(.A(ori_ori_n241_), .Y(ori_ori_n242_));
  NO3        o214(.A(ori_ori_n242_), .B(ori_ori_n238_), .C(ori_ori_n237_), .Y(ori_ori_n243_));
  NA4        o215(.A(ori_ori_n243_), .B(ori_ori_n236_), .C(ori_ori_n233_), .D(ori_ori_n227_), .Y(ori09));
  INV        o216(.A(ori_ori_n188_), .Y(ori_ori_n245_));
  NA2        o217(.A(c), .B(ori_ori_n45_), .Y(ori_ori_n246_));
  NO2        o218(.A(ori_ori_n246_), .B(ori_ori_n143_), .Y(ori_ori_n247_));
  NA3        o219(.A(ori_ori_n247_), .B(ori_ori_n167_), .C(f), .Y(ori_ori_n248_));
  INV        o220(.A(ori_ori_n248_), .Y(ori_ori_n249_));
  NO2        o221(.A(ori_ori_n249_), .B(ori_ori_n245_), .Y(ori_ori_n250_));
  NO2        o222(.A(ori_ori_n88_), .B(ori_ori_n82_), .Y(ori_ori_n251_));
  NA2        o223(.A(ori_ori_n251_), .B(ori_ori_n85_), .Y(ori_ori_n252_));
  INV        o224(.A(ori_ori_n252_), .Y(ori_ori_n253_));
  NA2        o225(.A(e), .B(d), .Y(ori_ori_n254_));
  OAI220     o226(.A0(ori_ori_n254_), .A1(c), .B0(ori_ori_n115_), .B1(d), .Y(ori_ori_n255_));
  NA3        o227(.A(ori_ori_n255_), .B(ori_ori_n151_), .C(ori_ori_n165_), .Y(ori_ori_n256_));
  AOI210     o228(.A0(ori_ori_n172_), .A1(ori_ori_n64_), .B0(ori_ori_n88_), .Y(ori_ori_n257_));
  INV        o229(.A(ori_ori_n257_), .Y(ori_ori_n258_));
  NA2        o230(.A(ori_ori_n258_), .B(ori_ori_n256_), .Y(ori_ori_n259_));
  NO2        o231(.A(ori_ori_n259_), .B(ori_ori_n253_), .Y(ori_ori_n260_));
  NA2        o232(.A(ori_ori_n181_), .B(ori_ori_n187_), .Y(ori_ori_n261_));
  AO220      o233(.A0(ori_ori_n151_), .A1(ori_ori_n230_), .B0(ori_ori_n60_), .B1(f), .Y(ori_ori_n262_));
  OAI210     o234(.A0(ori_ori_n262_), .A1(ori_ori_n154_), .B0(ori_ori_n255_), .Y(ori_ori_n263_));
  AN2        o235(.A(ori_ori_n263_), .B(ori_ori_n261_), .Y(ori_ori_n264_));
  NA3        o236(.A(ori_ori_n264_), .B(ori_ori_n260_), .C(ori_ori_n250_), .Y(ori12));
  NO4        o237(.A(ori_ori_n145_), .B(ori_ori_n98_), .C(ori_ori_n180_), .D(ori_ori_n78_), .Y(ori_ori_n266_));
  AOI210     o238(.A0(ori_ori_n90_), .A1(ori_ori_n121_), .B0(ori_ori_n76_), .Y(ori_ori_n267_));
  OR2        o239(.A(ori_ori_n267_), .B(ori_ori_n266_), .Y(ori_ori_n268_));
  AOI210     o240(.A0(ori_ori_n119_), .A1(ori_ori_n132_), .B0(ori_ori_n78_), .Y(ori_ori_n269_));
  OAI210     o241(.A0(ori_ori_n269_), .A1(ori_ori_n268_), .B0(ori_ori_n140_), .Y(ori_ori_n270_));
  INV        o242(.A(ori_ori_n124_), .Y(ori_ori_n271_));
  NA2        o243(.A(ori_ori_n46_), .B(g), .Y(ori_ori_n272_));
  AOI210     o244(.A0(ori_ori_n205_), .A1(ori_ori_n272_), .B0(m), .Y(ori_ori_n273_));
  NA2        o245(.A(ori_ori_n273_), .B(ori_ori_n116_), .Y(ori_ori_n274_));
  NO2        o246(.A(ori_ori_n156_), .B(ori_ori_n78_), .Y(ori_ori_n275_));
  NA2        o247(.A(ori_ori_n88_), .B(ori_ori_n56_), .Y(ori_ori_n276_));
  NO2        o248(.A(ori_ori_n111_), .B(ori_ori_n60_), .Y(ori_ori_n277_));
  NOi31      o249(.An(ori_ori_n276_), .B(ori_ori_n277_), .C(ori_ori_n78_), .Y(ori_ori_n278_));
  NAi21      o250(.An(ori_ori_n179_), .B(ori_ori_n275_), .Y(ori_ori_n279_));
  NA2        o251(.A(ori_ori_n161_), .B(g), .Y(ori_ori_n280_));
  NA2        o252(.A(ori_ori_n280_), .B(ori_ori_n279_), .Y(ori_ori_n281_));
  OAI210     o253(.A0(ori_ori_n267_), .A1(ori_ori_n266_), .B0(ori_ori_n276_), .Y(ori_ori_n282_));
  NA3        o254(.A(ori_ori_n271_), .B(ori_ori_n162_), .C(ori_ori_n31_), .Y(ori_ori_n283_));
  NA2        o255(.A(ori_ori_n283_), .B(ori_ori_n282_), .Y(ori_ori_n284_));
  NO3        o256(.A(ori_ori_n284_), .B(ori_ori_n281_), .C(ori_ori_n278_), .Y(ori_ori_n285_));
  NA3        o257(.A(ori_ori_n285_), .B(ori_ori_n274_), .C(ori_ori_n270_), .Y(ori13));
  NAi21      o258(.An(c), .B(e), .Y(ori_ori_n287_));
  AN2        o259(.A(d), .B(c), .Y(ori_ori_n288_));
  NA2        o260(.A(ori_ori_n288_), .B(ori_ori_n45_), .Y(ori_ori_n289_));
  NAi32      o261(.An(f), .Bn(e), .C(c), .Y(ori_ori_n290_));
  NO3        o262(.A(m), .B(i), .C(h), .Y(ori_ori_n291_));
  NA3        o263(.A(k), .B(j), .C(i), .Y(ori_ori_n292_));
  NO2        o264(.A(f), .B(c), .Y(ori_ori_n293_));
  NOi21      o265(.An(ori_ori_n293_), .B(ori_ori_n145_), .Y(ori_ori_n294_));
  AN3        o266(.A(g), .B(f), .C(c), .Y(ori_ori_n295_));
  NA3        o267(.A(l), .B(k), .C(j), .Y(ori_ori_n296_));
  NA2        o268(.A(i), .B(h), .Y(ori_ori_n297_));
  NO3        o269(.A(ori_ori_n297_), .B(ori_ori_n296_), .C(ori_ori_n48_), .Y(ori_ori_n298_));
  NO2        o270(.A(ori_ori_n107_), .B(ori_ori_n78_), .Y(ori_ori_n299_));
  NOi21      o271(.An(m), .B(n), .Y(ori_ori_n300_));
  NA2        o272(.A(ori_ori_n167_), .B(f), .Y(ori_ori_n301_));
  NO2        o273(.A(ori_ori_n301_), .B(ori_ori_n289_), .Y(ori_ori_n302_));
  INV        o274(.A(ori_ori_n302_), .Y(ori_ori_n303_));
  INV        o275(.A(h), .Y(ori_ori_n304_));
  NA2        o276(.A(ori_ori_n194_), .B(ori_ori_n95_), .Y(ori_ori_n305_));
  NA2        o277(.A(ori_ori_n305_), .B(ori_ori_n303_), .Y(ori01));
  INV        o278(.A(ori_ori_n106_), .Y(ori_ori_n307_));
  NA2        o279(.A(ori_ori_n137_), .B(i), .Y(ori_ori_n308_));
  NA2        o280(.A(ori_ori_n308_), .B(ori_ori_n307_), .Y(ori_ori_n309_));
  INV        o281(.A(ori_ori_n261_), .Y(ori_ori_n310_));
  INV        o282(.A(ori_ori_n252_), .Y(ori_ori_n311_));
  INV        o283(.A(ori_ori_n170_), .Y(ori_ori_n312_));
  OR2        o284(.A(ori_ori_n72_), .B(ori_ori_n70_), .Y(ori_ori_n313_));
  NA2        o285(.A(ori_ori_n313_), .B(ori_ori_n312_), .Y(ori_ori_n314_));
  NO4        o286(.A(ori_ori_n314_), .B(ori_ori_n311_), .C(ori_ori_n310_), .D(ori_ori_n309_), .Y(ori_ori_n315_));
  NA2        o287(.A(ori_ori_n105_), .B(ori_ori_n72_), .Y(ori_ori_n316_));
  NA2        o288(.A(ori_ori_n316_), .B(ori_ori_n201_), .Y(ori_ori_n317_));
  NO3        o289(.A(ori_ori_n297_), .B(ori_ori_n61_), .C(ori_ori_n40_), .Y(ori_ori_n318_));
  NO2        o290(.A(ori_ori_n183_), .B(ori_ori_n182_), .Y(ori_ori_n319_));
  NO4        o291(.A(ori_ori_n297_), .B(ori_ori_n319_), .C(ori_ori_n59_), .D(ori_ori_n40_), .Y(ori_ori_n320_));
  INV        o292(.A(ori_ori_n320_), .Y(ori_ori_n321_));
  NA4        o293(.A(ori_ori_n321_), .B(ori_ori_n129_), .C(ori_ori_n317_), .D(ori_ori_n315_), .Y(ori06));
  NO2        o294(.A(ori_ori_n82_), .B(ori_ori_n41_), .Y(ori_ori_n323_));
  OAI210     o295(.A0(ori_ori_n323_), .A1(ori_ori_n318_), .B0(ori_ori_n125_), .Y(ori_ori_n324_));
  INV        o296(.A(ori_ori_n324_), .Y(ori_ori_n325_));
  NO2        o297(.A(ori_ori_n325_), .B(ori_ori_n102_), .Y(ori_ori_n326_));
  NO2        o298(.A(ori_ori_n172_), .B(ori_ori_n56_), .Y(ori_ori_n327_));
  NO2        o299(.A(ori_ori_n157_), .B(ori_ori_n97_), .Y(ori_ori_n328_));
  NO2        o300(.A(ori_ori_n328_), .B(ori_ori_n327_), .Y(ori_ori_n329_));
  OAI220     o301(.A0(ori_ori_n217_), .A1(ori_ori_n97_), .B0(ori_ori_n169_), .B1(ori_ori_n172_), .Y(ori_ori_n330_));
  NAi21      o302(.An(j), .B(i), .Y(ori_ori_n331_));
  NO4        o303(.A(ori_ori_n319_), .B(ori_ori_n331_), .C(ori_ori_n145_), .D(ori_ori_n91_), .Y(ori_ori_n332_));
  NO3        o304(.A(ori_ori_n332_), .B(ori_ori_n161_), .C(ori_ori_n330_), .Y(ori_ori_n333_));
  NA4        o305(.A(ori_ori_n333_), .B(ori_ori_n329_), .C(ori_ori_n326_), .D(ori_ori_n321_), .Y(ori07));
  NOi31      o306(.An(n), .B(m), .C(b), .Y(ori_ori_n335_));
  NO3        o307(.A(n), .B(m), .C(h), .Y(ori_ori_n336_));
  NO2        o308(.A(ori_ori_n290_), .B(ori_ori_n145_), .Y(ori_ori_n337_));
  NO2        o309(.A(ori_ori_n292_), .B(ori_ori_n110_), .Y(ori_ori_n338_));
  INV        o310(.A(ori_ori_n337_), .Y(ori_ori_n339_));
  NO2        o311(.A(e), .B(c), .Y(ori_ori_n340_));
  NO2        o312(.A(ori_ori_n48_), .B(ori_ori_n78_), .Y(ori_ori_n341_));
  NA2        o313(.A(ori_ori_n341_), .B(ori_ori_n340_), .Y(ori_ori_n342_));
  INV        o314(.A(ori_ori_n342_), .Y(ori_ori_n343_));
  NA2        o315(.A(ori_ori_n214_), .B(ori_ori_n207_), .Y(ori_ori_n344_));
  INV        o316(.A(ori_ori_n344_), .Y(ori_ori_n345_));
  NO2        o317(.A(l), .B(k), .Y(ori_ori_n346_));
  NO3        o318(.A(ori_ori_n145_), .B(d), .C(c), .Y(ori_ori_n347_));
  NO2        o319(.A(ori_ori_n345_), .B(ori_ori_n343_), .Y(ori_ori_n348_));
  NOi31      o320(.An(m), .B(n), .C(b), .Y(ori_ori_n349_));
  NA2        o321(.A(ori_ori_n295_), .B(ori_ori_n159_), .Y(ori_ori_n350_));
  NO2        o322(.A(ori_ori_n350_), .B(ori_ori_n145_), .Y(ori_ori_n351_));
  NO2        o323(.A(ori_ori_n291_), .B(ori_ori_n351_), .Y(ori_ori_n352_));
  NA2        o324(.A(ori_ori_n336_), .B(ori_ori_n346_), .Y(ori_ori_n353_));
  INV        o325(.A(ori_ori_n353_), .Y(ori_ori_n354_));
  NA2        o326(.A(ori_ori_n300_), .B(ori_ori_n143_), .Y(ori_ori_n355_));
  INV        o327(.A(ori_ori_n355_), .Y(ori_ori_n356_));
  OR2        o328(.A(ori_ori_n356_), .B(ori_ori_n354_), .Y(ori_ori_n357_));
  NO2        o329(.A(ori_ori_n357_), .B(ori_ori_n298_), .Y(ori_ori_n358_));
  NA4        o330(.A(ori_ori_n358_), .B(ori_ori_n352_), .C(ori_ori_n348_), .D(ori_ori_n339_), .Y(ori_ori_n359_));
  NO2        o331(.A(ori_ori_n134_), .B(j), .Y(ori_ori_n360_));
  NA2        o332(.A(ori_ori_n360_), .B(ori_ori_n52_), .Y(ori_ori_n361_));
  INV        o333(.A(ori_ori_n361_), .Y(ori_ori_n362_));
  NO2        o334(.A(ori_ori_n362_), .B(ori_ori_n294_), .Y(ori_ori_n363_));
  INV        o335(.A(ori_ori_n32_), .Y(ori_ori_n364_));
  NA2        o336(.A(ori_ori_n364_), .B(ori_ori_n304_), .Y(ori_ori_n365_));
  INV        o337(.A(ori_ori_n365_), .Y(ori_ori_n366_));
  NO2        o338(.A(ori_ori_n82_), .B(ori_ori_n61_), .Y(ori_ori_n367_));
  NO2        o339(.A(ori_ori_n367_), .B(ori_ori_n366_), .Y(ori_ori_n368_));
  INV        o340(.A(a), .Y(ori_ori_n369_));
  NO2        o341(.A(ori_ori_n396_), .B(ori_ori_n369_), .Y(ori_ori_n370_));
  NO2        o342(.A(ori_ori_n331_), .B(ori_ori_n59_), .Y(ori_ori_n371_));
  NA2        o343(.A(h), .B(ori_ori_n371_), .Y(ori_ori_n372_));
  INV        o344(.A(ori_ori_n372_), .Y(ori_ori_n373_));
  NO2        o345(.A(ori_ori_n373_), .B(ori_ori_n370_), .Y(ori_ori_n374_));
  NA3        o346(.A(ori_ori_n374_), .B(ori_ori_n368_), .C(ori_ori_n363_), .Y(ori_ori_n375_));
  NA2        o347(.A(h), .B(ori_ori_n338_), .Y(ori_ori_n376_));
  NA2        o348(.A(ori_ori_n335_), .B(ori_ori_n246_), .Y(ori_ori_n377_));
  NO2        o349(.A(ori_ori_n287_), .B(ori_ori_n48_), .Y(ori_ori_n378_));
  NA2        o350(.A(ori_ori_n378_), .B(f), .Y(ori_ori_n379_));
  NA3        o351(.A(ori_ori_n379_), .B(ori_ori_n377_), .C(ori_ori_n376_), .Y(ori_ori_n380_));
  NA2        o352(.A(ori_ori_n299_), .B(ori_ori_n81_), .Y(ori_ori_n381_));
  INV        o353(.A(ori_ori_n349_), .Y(ori_ori_n382_));
  NA2        o354(.A(ori_ori_n382_), .B(ori_ori_n381_), .Y(ori_ori_n383_));
  NO2        o355(.A(ori_ori_n383_), .B(ori_ori_n380_), .Y(ori_ori_n384_));
  INV        o356(.A(ori_ori_n190_), .Y(ori_ori_n385_));
  BUFFER     o357(.A(ori_ori_n48_), .Y(ori_ori_n386_));
  OAI210     o358(.A0(ori_ori_n386_), .A1(f), .B0(ori_ori_n385_), .Y(ori_ori_n387_));
  INV        o359(.A(ori_ori_n387_), .Y(ori_ori_n388_));
  OR2        o360(.A(h), .B(ori_ori_n178_), .Y(ori_ori_n389_));
  NO2        o361(.A(ori_ori_n389_), .B(ori_ori_n59_), .Y(ori_ori_n390_));
  NO2        o362(.A(ori_ori_n390_), .B(ori_ori_n347_), .Y(ori_ori_n391_));
  NA3        o363(.A(ori_ori_n391_), .B(ori_ori_n388_), .C(ori_ori_n384_), .Y(ori_ori_n392_));
  OR3        o364(.A(ori_ori_n392_), .B(ori_ori_n375_), .C(ori_ori_n359_), .Y(ori04));
  INV        o365(.A(ori_ori_n43_), .Y(ori_ori_n396_));
  ZERO       o366(.Y(ori02));
  ZERO       o367(.Y(ori03));
  ZERO       o368(.Y(ori00));
  ZERO       o369(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO4        m0025(.A(mai_mai_n53_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n54_));
  AOI210     m0026(.A0(mai_mai_n54_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NA3        m0031(.A(g), .B(mai_mai_n59_), .C(a), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(h), .Y(mai_mai_n61_));
  NAi31      m0033(.An(i), .B(l), .C(j), .Y(mai_mai_n62_));
  OAI220     m0034(.A0(mai_mai_n62_), .A1(mai_mai_n49_), .B0(mai_mai_n61_), .B1(mai_mai_n44_), .Y(mai_mai_n63_));
  NAi31      m0035(.An(mai_mai_n60_), .B(mai_mai_n63_), .C(mai_mai_n58_), .Y(mai_mai_n64_));
  NAi41      m0036(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n65_));
  NA2        m0037(.A(g), .B(f), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi21      m0039(.An(i), .B(j), .Y(mai_mai_n68_));
  NAi32      m0040(.An(n), .Bn(k), .C(m), .Y(mai_mai_n69_));
  NO2        m0041(.A(mai_mai_n69_), .B(mai_mai_n68_), .Y(mai_mai_n70_));
  NAi31      m0042(.An(l), .B(m), .C(k), .Y(mai_mai_n71_));
  NAi21      m0043(.An(e), .B(h), .Y(mai_mai_n72_));
  NAi41      m0044(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n74_));
  INV        m0046(.A(m), .Y(mai_mai_n75_));
  NOi21      m0047(.An(k), .B(l), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n77_));
  AN4        m0049(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n78_));
  NOi31      m0050(.An(h), .B(g), .C(f), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  NAi32      m0052(.An(m), .Bn(k), .C(j), .Y(mai_mai_n81_));
  NOi32      m0053(.An(h), .Bn(g), .C(f), .Y(mai_mai_n82_));
  NA2        m0054(.A(mai_mai_n82_), .B(mai_mai_n78_), .Y(mai_mai_n83_));
  OA220      m0055(.A0(mai_mai_n83_), .A1(mai_mai_n81_), .B0(mai_mai_n80_), .B1(mai_mai_n77_), .Y(mai_mai_n84_));
  NA3        m0056(.A(mai_mai_n84_), .B(mai_mai_n74_), .C(mai_mai_n64_), .Y(mai_mai_n85_));
  INV        m0057(.A(n), .Y(mai_mai_n86_));
  NOi32      m0058(.An(e), .Bn(b), .C(d), .Y(mai_mai_n87_));
  NA2        m0059(.A(mai_mai_n87_), .B(mai_mai_n86_), .Y(mai_mai_n88_));
  INV        m0060(.A(j), .Y(mai_mai_n89_));
  AN3        m0061(.A(m), .B(k), .C(i), .Y(mai_mai_n90_));
  NA3        m0062(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(g), .Y(mai_mai_n91_));
  NO2        m0063(.A(mai_mai_n91_), .B(f), .Y(mai_mai_n92_));
  NAi32      m0064(.An(g), .Bn(f), .C(h), .Y(mai_mai_n93_));
  NAi31      m0065(.An(j), .B(m), .C(l), .Y(mai_mai_n94_));
  NO2        m0066(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n95_));
  NA2        m0067(.A(m), .B(l), .Y(mai_mai_n96_));
  NAi31      m0068(.An(k), .B(j), .C(g), .Y(mai_mai_n97_));
  NO3        m0069(.A(mai_mai_n97_), .B(mai_mai_n96_), .C(f), .Y(mai_mai_n98_));
  AN2        m0070(.A(j), .B(g), .Y(mai_mai_n99_));
  NOi21      m0071(.An(g), .B(i), .Y(mai_mai_n100_));
  NOi32      m0072(.An(m), .Bn(j), .C(k), .Y(mai_mai_n101_));
  AOI220     m0073(.A0(mai_mai_n101_), .A1(mai_mai_n100_), .B0(m), .B1(mai_mai_n99_), .Y(mai_mai_n102_));
  NO2        m0074(.A(mai_mai_n102_), .B(f), .Y(mai_mai_n103_));
  NO4        m0075(.A(mai_mai_n103_), .B(mai_mai_n98_), .C(mai_mai_n95_), .D(mai_mai_n92_), .Y(mai_mai_n104_));
  NAi41      m0076(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n105_));
  AN2        m0077(.A(e), .B(b), .Y(mai_mai_n106_));
  NOi31      m0078(.An(c), .B(h), .C(f), .Y(mai_mai_n107_));
  NA2        m0079(.A(mai_mai_n107_), .B(mai_mai_n106_), .Y(mai_mai_n108_));
  NO3        m0080(.A(mai_mai_n108_), .B(mai_mai_n105_), .C(g), .Y(mai_mai_n109_));
  NOi21      m0081(.An(i), .B(h), .Y(mai_mai_n110_));
  NA3        m0082(.A(mai_mai_n110_), .B(g), .C(mai_mai_n36_), .Y(mai_mai_n111_));
  INV        m0083(.A(a), .Y(mai_mai_n112_));
  NA2        m0084(.A(mai_mai_n106_), .B(mai_mai_n112_), .Y(mai_mai_n113_));
  INV        m0085(.A(l), .Y(mai_mai_n114_));
  NOi21      m0086(.An(m), .B(n), .Y(mai_mai_n115_));
  AN2        m0087(.A(k), .B(h), .Y(mai_mai_n116_));
  NO2        m0088(.A(mai_mai_n111_), .B(mai_mai_n88_), .Y(mai_mai_n117_));
  INV        m0089(.A(b), .Y(mai_mai_n118_));
  NA2        m0090(.A(l), .B(j), .Y(mai_mai_n119_));
  AN2        m0091(.A(k), .B(i), .Y(mai_mai_n120_));
  NA2        m0092(.A(g), .B(e), .Y(mai_mai_n121_));
  NOi32      m0093(.An(c), .Bn(a), .C(d), .Y(mai_mai_n122_));
  NA2        m0094(.A(mai_mai_n122_), .B(mai_mai_n115_), .Y(mai_mai_n123_));
  NO4        m0095(.A(mai_mai_n123_), .B(mai_mai_n121_), .C(mai_mai_n119_), .D(mai_mai_n118_), .Y(mai_mai_n124_));
  NO3        m0096(.A(mai_mai_n124_), .B(mai_mai_n117_), .C(mai_mai_n109_), .Y(mai_mai_n125_));
  OAI210     m0097(.A0(mai_mai_n104_), .A1(mai_mai_n88_), .B0(mai_mai_n125_), .Y(mai_mai_n126_));
  NOi31      m0098(.An(k), .B(m), .C(j), .Y(mai_mai_n127_));
  NA3        m0099(.A(mai_mai_n127_), .B(mai_mai_n79_), .C(mai_mai_n78_), .Y(mai_mai_n128_));
  NOi31      m0100(.An(k), .B(m), .C(i), .Y(mai_mai_n129_));
  NA3        m0101(.A(mai_mai_n129_), .B(mai_mai_n82_), .C(mai_mai_n78_), .Y(mai_mai_n130_));
  NA2        m0102(.A(mai_mai_n130_), .B(mai_mai_n128_), .Y(mai_mai_n131_));
  NOi32      m0103(.An(f), .Bn(b), .C(e), .Y(mai_mai_n132_));
  NAi21      m0104(.An(g), .B(h), .Y(mai_mai_n133_));
  NAi21      m0105(.An(m), .B(n), .Y(mai_mai_n134_));
  NAi21      m0106(.An(j), .B(k), .Y(mai_mai_n135_));
  NO3        m0107(.A(mai_mai_n135_), .B(mai_mai_n134_), .C(mai_mai_n133_), .Y(mai_mai_n136_));
  NAi41      m0108(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n137_));
  NAi31      m0109(.An(j), .B(k), .C(h), .Y(mai_mai_n138_));
  NO3        m0110(.A(mai_mai_n138_), .B(mai_mai_n137_), .C(mai_mai_n134_), .Y(mai_mai_n139_));
  AOI210     m0111(.A0(mai_mai_n136_), .A1(mai_mai_n132_), .B0(mai_mai_n139_), .Y(mai_mai_n140_));
  NO2        m0112(.A(k), .B(j), .Y(mai_mai_n141_));
  NO2        m0113(.A(mai_mai_n141_), .B(mai_mai_n134_), .Y(mai_mai_n142_));
  AN2        m0114(.A(k), .B(j), .Y(mai_mai_n143_));
  NAi21      m0115(.An(c), .B(b), .Y(mai_mai_n144_));
  NA2        m0116(.A(f), .B(d), .Y(mai_mai_n145_));
  NO4        m0117(.A(mai_mai_n145_), .B(mai_mai_n144_), .C(mai_mai_n143_), .D(mai_mai_n133_), .Y(mai_mai_n146_));
  NAi31      m0118(.An(f), .B(e), .C(b), .Y(mai_mai_n147_));
  NA2        m0119(.A(mai_mai_n146_), .B(mai_mai_n142_), .Y(mai_mai_n148_));
  NA2        m0120(.A(d), .B(b), .Y(mai_mai_n149_));
  NAi21      m0121(.An(e), .B(f), .Y(mai_mai_n150_));
  NO2        m0122(.A(mai_mai_n150_), .B(mai_mai_n149_), .Y(mai_mai_n151_));
  NA2        m0123(.A(b), .B(a), .Y(mai_mai_n152_));
  NAi21      m0124(.An(e), .B(g), .Y(mai_mai_n153_));
  NAi21      m0125(.An(c), .B(d), .Y(mai_mai_n154_));
  NAi31      m0126(.An(l), .B(k), .C(h), .Y(mai_mai_n155_));
  NO2        m0127(.A(mai_mai_n134_), .B(mai_mai_n155_), .Y(mai_mai_n156_));
  NA2        m0128(.A(mai_mai_n156_), .B(mai_mai_n151_), .Y(mai_mai_n157_));
  NAi41      m0129(.An(mai_mai_n131_), .B(mai_mai_n157_), .C(mai_mai_n148_), .D(mai_mai_n140_), .Y(mai_mai_n158_));
  NAi31      m0130(.An(e), .B(f), .C(b), .Y(mai_mai_n159_));
  NOi21      m0131(.An(g), .B(d), .Y(mai_mai_n160_));
  NO2        m0132(.A(mai_mai_n160_), .B(mai_mai_n159_), .Y(mai_mai_n161_));
  NOi21      m0133(.An(h), .B(i), .Y(mai_mai_n162_));
  NOi21      m0134(.An(k), .B(m), .Y(mai_mai_n163_));
  NA3        m0135(.A(mai_mai_n163_), .B(mai_mai_n162_), .C(n), .Y(mai_mai_n164_));
  NOi21      m0136(.An(mai_mai_n161_), .B(mai_mai_n164_), .Y(mai_mai_n165_));
  NO2        m0137(.A(mai_mai_n145_), .B(mai_mai_n144_), .Y(mai_mai_n166_));
  NA2        m0138(.A(mai_mai_n166_), .B(h), .Y(mai_mai_n167_));
  INV        m0139(.A(mai_mai_n49_), .Y(mai_mai_n168_));
  NA2        m0140(.A(mai_mai_n168_), .B(mai_mai_n67_), .Y(mai_mai_n169_));
  NOi32      m0141(.An(n), .Bn(k), .C(m), .Y(mai_mai_n170_));
  NA2        m0142(.A(l), .B(i), .Y(mai_mai_n171_));
  NA2        m0143(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  OAI210     m0144(.A0(mai_mai_n172_), .A1(mai_mai_n167_), .B0(mai_mai_n169_), .Y(mai_mai_n173_));
  NAi31      m0145(.An(d), .B(f), .C(c), .Y(mai_mai_n174_));
  NAi31      m0146(.An(e), .B(f), .C(c), .Y(mai_mai_n175_));
  NA2        m0147(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  NA2        m0148(.A(j), .B(h), .Y(mai_mai_n177_));
  OR3        m0149(.A(n), .B(m), .C(k), .Y(mai_mai_n178_));
  NO2        m0150(.A(mai_mai_n178_), .B(mai_mai_n177_), .Y(mai_mai_n179_));
  NAi32      m0151(.An(m), .Bn(k), .C(n), .Y(mai_mai_n180_));
  NO2        m0152(.A(mai_mai_n180_), .B(mai_mai_n177_), .Y(mai_mai_n181_));
  AOI220     m0153(.A0(mai_mai_n181_), .A1(mai_mai_n161_), .B0(mai_mai_n179_), .B1(mai_mai_n176_), .Y(mai_mai_n182_));
  NO2        m0154(.A(n), .B(m), .Y(mai_mai_n183_));
  NA2        m0155(.A(mai_mai_n183_), .B(mai_mai_n50_), .Y(mai_mai_n184_));
  NAi21      m0156(.An(f), .B(e), .Y(mai_mai_n185_));
  NA2        m0157(.A(d), .B(c), .Y(mai_mai_n186_));
  NO2        m0158(.A(mai_mai_n186_), .B(mai_mai_n185_), .Y(mai_mai_n187_));
  NOi21      m0159(.An(mai_mai_n187_), .B(mai_mai_n184_), .Y(mai_mai_n188_));
  NAi21      m0160(.An(d), .B(c), .Y(mai_mai_n189_));
  NAi31      m0161(.An(m), .B(n), .C(b), .Y(mai_mai_n190_));
  NA2        m0162(.A(k), .B(i), .Y(mai_mai_n191_));
  NAi21      m0163(.An(h), .B(f), .Y(mai_mai_n192_));
  NO2        m0164(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n193_));
  NO2        m0165(.A(mai_mai_n190_), .B(mai_mai_n154_), .Y(mai_mai_n194_));
  NA2        m0166(.A(mai_mai_n194_), .B(mai_mai_n193_), .Y(mai_mai_n195_));
  NOi32      m0167(.An(f), .Bn(c), .C(d), .Y(mai_mai_n196_));
  NOi32      m0168(.An(f), .Bn(c), .C(e), .Y(mai_mai_n197_));
  NO2        m0169(.A(mai_mai_n197_), .B(mai_mai_n196_), .Y(mai_mai_n198_));
  NO3        m0170(.A(n), .B(m), .C(j), .Y(mai_mai_n199_));
  NA2        m0171(.A(mai_mai_n199_), .B(mai_mai_n116_), .Y(mai_mai_n200_));
  AO210      m0172(.A0(mai_mai_n200_), .A1(mai_mai_n184_), .B0(mai_mai_n198_), .Y(mai_mai_n201_));
  NAi41      m0173(.An(mai_mai_n188_), .B(mai_mai_n201_), .C(mai_mai_n195_), .D(mai_mai_n182_), .Y(mai_mai_n202_));
  OR4        m0174(.A(mai_mai_n202_), .B(mai_mai_n173_), .C(mai_mai_n165_), .D(mai_mai_n158_), .Y(mai_mai_n203_));
  NO4        m0175(.A(mai_mai_n203_), .B(mai_mai_n126_), .C(mai_mai_n85_), .D(mai_mai_n55_), .Y(mai_mai_n204_));
  NAi31      m0176(.An(n), .B(h), .C(g), .Y(mai_mai_n205_));
  NO2        m0177(.A(mai_mai_n205_), .B(mai_mai_n1460_), .Y(mai_mai_n206_));
  NOi32      m0178(.An(m), .Bn(k), .C(l), .Y(mai_mai_n207_));
  NA3        m0179(.A(mai_mai_n207_), .B(mai_mai_n89_), .C(g), .Y(mai_mai_n208_));
  NO2        m0180(.A(mai_mai_n208_), .B(n), .Y(mai_mai_n209_));
  NOi21      m0181(.An(k), .B(j), .Y(mai_mai_n210_));
  NA4        m0182(.A(mai_mai_n210_), .B(mai_mai_n115_), .C(i), .D(g), .Y(mai_mai_n211_));
  AN2        m0183(.A(i), .B(g), .Y(mai_mai_n212_));
  NA3        m0184(.A(mai_mai_n76_), .B(mai_mai_n212_), .C(mai_mai_n115_), .Y(mai_mai_n213_));
  NA2        m0185(.A(mai_mai_n213_), .B(mai_mai_n211_), .Y(mai_mai_n214_));
  NO3        m0186(.A(mai_mai_n214_), .B(mai_mai_n209_), .C(mai_mai_n206_), .Y(mai_mai_n215_));
  NAi41      m0187(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n216_));
  INV        m0188(.A(mai_mai_n216_), .Y(mai_mai_n217_));
  INV        m0189(.A(f), .Y(mai_mai_n218_));
  INV        m0190(.A(g), .Y(mai_mai_n219_));
  NOi31      m0191(.An(i), .B(j), .C(h), .Y(mai_mai_n220_));
  NOi21      m0192(.An(l), .B(m), .Y(mai_mai_n221_));
  NA2        m0193(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n222_));
  NO3        m0194(.A(mai_mai_n222_), .B(mai_mai_n219_), .C(mai_mai_n218_), .Y(mai_mai_n223_));
  NA2        m0195(.A(mai_mai_n223_), .B(mai_mai_n217_), .Y(mai_mai_n224_));
  OAI210     m0196(.A0(mai_mai_n215_), .A1(mai_mai_n32_), .B0(mai_mai_n224_), .Y(mai_mai_n225_));
  NOi21      m0197(.An(n), .B(m), .Y(mai_mai_n226_));
  NOi32      m0198(.An(l), .Bn(i), .C(j), .Y(mai_mai_n227_));
  NA2        m0199(.A(mai_mai_n227_), .B(mai_mai_n226_), .Y(mai_mai_n228_));
  OA220      m0200(.A0(mai_mai_n228_), .A1(mai_mai_n108_), .B0(mai_mai_n81_), .B1(mai_mai_n80_), .Y(mai_mai_n229_));
  NAi21      m0201(.An(j), .B(h), .Y(mai_mai_n230_));
  XN2        m0202(.A(i), .B(h), .Y(mai_mai_n231_));
  NAi31      m0203(.An(f), .B(e), .C(c), .Y(mai_mai_n232_));
  NO4        m0204(.A(mai_mai_n232_), .B(mai_mai_n178_), .C(mai_mai_n177_), .D(mai_mai_n59_), .Y(mai_mai_n233_));
  NA4        m0205(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n234_));
  NAi32      m0206(.An(m), .Bn(i), .C(k), .Y(mai_mai_n235_));
  NO3        m0207(.A(mai_mai_n235_), .B(mai_mai_n93_), .C(mai_mai_n234_), .Y(mai_mai_n236_));
  NA2        m0208(.A(k), .B(h), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n236_), .B(mai_mai_n233_), .Y(mai_mai_n238_));
  NAi21      m0210(.An(n), .B(a), .Y(mai_mai_n239_));
  NO2        m0211(.A(mai_mai_n239_), .B(mai_mai_n149_), .Y(mai_mai_n240_));
  NAi41      m0212(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n241_), .B(e), .Y(mai_mai_n242_));
  NO3        m0214(.A(mai_mai_n150_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n243_));
  OAI210     m0215(.A0(mai_mai_n243_), .A1(mai_mai_n242_), .B0(mai_mai_n240_), .Y(mai_mai_n244_));
  AN3        m0216(.A(mai_mai_n244_), .B(mai_mai_n238_), .C(mai_mai_n229_), .Y(mai_mai_n245_));
  OR2        m0217(.A(h), .B(g), .Y(mai_mai_n246_));
  NO2        m0218(.A(mai_mai_n246_), .B(mai_mai_n105_), .Y(mai_mai_n247_));
  NAi41      m0219(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n248_));
  NO2        m0220(.A(mai_mai_n248_), .B(mai_mai_n218_), .Y(mai_mai_n249_));
  NA2        m0221(.A(mai_mai_n163_), .B(mai_mai_n110_), .Y(mai_mai_n250_));
  NAi21      m0222(.An(mai_mai_n250_), .B(mai_mai_n249_), .Y(mai_mai_n251_));
  NO2        m0223(.A(n), .B(a), .Y(mai_mai_n252_));
  NAi31      m0224(.An(mai_mai_n241_), .B(mai_mai_n252_), .C(mai_mai_n106_), .Y(mai_mai_n253_));
  AN2        m0225(.A(mai_mai_n253_), .B(mai_mai_n251_), .Y(mai_mai_n254_));
  NAi21      m0226(.An(h), .B(i), .Y(mai_mai_n255_));
  NA2        m0227(.A(mai_mai_n183_), .B(k), .Y(mai_mai_n256_));
  NO2        m0228(.A(mai_mai_n256_), .B(mai_mai_n255_), .Y(mai_mai_n257_));
  NA2        m0229(.A(mai_mai_n257_), .B(mai_mai_n196_), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n258_), .B(mai_mai_n254_), .Y(mai_mai_n259_));
  NOi21      m0231(.An(g), .B(e), .Y(mai_mai_n260_));
  NO2        m0232(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n261_));
  NO2        m0233(.A(mai_mai_n255_), .B(mai_mai_n44_), .Y(mai_mai_n262_));
  NAi21      m0234(.An(f), .B(g), .Y(mai_mai_n263_));
  NO2        m0235(.A(mai_mai_n263_), .B(mai_mai_n65_), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n69_), .B(mai_mai_n119_), .Y(mai_mai_n265_));
  AOI220     m0237(.A0(mai_mai_n265_), .A1(mai_mai_n264_), .B0(mai_mai_n262_), .B1(mai_mai_n67_), .Y(mai_mai_n266_));
  INV        m0238(.A(mai_mai_n266_), .Y(mai_mai_n267_));
  NO3        m0239(.A(mai_mai_n135_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n268_));
  NOi41      m0240(.An(mai_mai_n245_), .B(mai_mai_n267_), .C(mai_mai_n259_), .D(mai_mai_n225_), .Y(mai_mai_n269_));
  NO4        m0241(.A(mai_mai_n206_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n270_));
  NO2        m0242(.A(mai_mai_n270_), .B(mai_mai_n113_), .Y(mai_mai_n271_));
  NAi21      m0243(.An(h), .B(g), .Y(mai_mai_n272_));
  OR4        m0244(.A(mai_mai_n272_), .B(mai_mai_n1465_), .C(mai_mai_n228_), .D(e), .Y(mai_mai_n273_));
  NO2        m0245(.A(mai_mai_n250_), .B(mai_mai_n263_), .Y(mai_mai_n274_));
  NA2        m0246(.A(mai_mai_n274_), .B(mai_mai_n78_), .Y(mai_mai_n275_));
  NAi31      m0247(.An(g), .B(k), .C(h), .Y(mai_mai_n276_));
  NAi31      m0248(.An(e), .B(d), .C(a), .Y(mai_mai_n277_));
  NA2        m0249(.A(mai_mai_n275_), .B(mai_mai_n273_), .Y(mai_mai_n278_));
  NA4        m0250(.A(mai_mai_n163_), .B(mai_mai_n82_), .C(mai_mai_n78_), .D(mai_mai_n119_), .Y(mai_mai_n279_));
  NA3        m0251(.A(mai_mai_n163_), .B(mai_mai_n162_), .C(mai_mai_n86_), .Y(mai_mai_n280_));
  NO2        m0252(.A(mai_mai_n280_), .B(mai_mai_n198_), .Y(mai_mai_n281_));
  NA3        m0253(.A(e), .B(c), .C(b), .Y(mai_mai_n282_));
  NO2        m0254(.A(mai_mai_n60_), .B(mai_mai_n282_), .Y(mai_mai_n283_));
  NAi32      m0255(.An(k), .Bn(i), .C(j), .Y(mai_mai_n284_));
  INV        m0256(.A(mai_mai_n49_), .Y(mai_mai_n285_));
  OAI210     m0257(.A0(mai_mai_n264_), .A1(mai_mai_n283_), .B0(mai_mai_n285_), .Y(mai_mai_n286_));
  NAi21      m0258(.An(l), .B(k), .Y(mai_mai_n287_));
  NO2        m0259(.A(mai_mai_n287_), .B(mai_mai_n49_), .Y(mai_mai_n288_));
  NOi21      m0260(.An(l), .B(j), .Y(mai_mai_n289_));
  NA2        m0261(.A(h), .B(mai_mai_n289_), .Y(mai_mai_n290_));
  OR3        m0262(.A(mai_mai_n73_), .B(mai_mai_n75_), .C(e), .Y(mai_mai_n291_));
  NO2        m0263(.A(mai_mai_n290_), .B(mai_mai_n291_), .Y(mai_mai_n292_));
  INV        m0264(.A(mai_mai_n292_), .Y(mai_mai_n293_));
  NAi32      m0265(.An(j), .Bn(h), .C(i), .Y(mai_mai_n294_));
  NAi21      m0266(.An(m), .B(l), .Y(mai_mai_n295_));
  NO3        m0267(.A(mai_mai_n295_), .B(mai_mai_n294_), .C(mai_mai_n86_), .Y(mai_mai_n296_));
  NA2        m0268(.A(h), .B(g), .Y(mai_mai_n297_));
  NA2        m0269(.A(mai_mai_n170_), .B(mai_mai_n45_), .Y(mai_mai_n298_));
  NO2        m0270(.A(mai_mai_n298_), .B(mai_mai_n297_), .Y(mai_mai_n299_));
  OAI210     m0271(.A0(mai_mai_n299_), .A1(mai_mai_n296_), .B0(mai_mai_n166_), .Y(mai_mai_n300_));
  NA4        m0272(.A(mai_mai_n300_), .B(mai_mai_n293_), .C(mai_mai_n286_), .D(mai_mai_n279_), .Y(mai_mai_n301_));
  NO2        m0273(.A(mai_mai_n147_), .B(d), .Y(mai_mai_n302_));
  NA2        m0274(.A(mai_mai_n302_), .B(mai_mai_n53_), .Y(mai_mai_n303_));
  NO2        m0275(.A(mai_mai_n108_), .B(mai_mai_n105_), .Y(mai_mai_n304_));
  NAi32      m0276(.An(n), .Bn(m), .C(l), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n305_), .B(mai_mai_n294_), .Y(mai_mai_n306_));
  AOI220     m0278(.A0(mai_mai_n306_), .A1(mai_mai_n187_), .B0(mai_mai_n304_), .B1(mai_mai_n59_), .Y(mai_mai_n307_));
  NO2        m0279(.A(mai_mai_n123_), .B(mai_mai_n118_), .Y(mai_mai_n308_));
  INV        m0280(.A(mai_mai_n121_), .Y(mai_mai_n309_));
  NA2        m0281(.A(mai_mai_n309_), .B(mai_mai_n308_), .Y(mai_mai_n310_));
  NA3        m0282(.A(mai_mai_n310_), .B(mai_mai_n307_), .C(mai_mai_n303_), .Y(mai_mai_n311_));
  NO4        m0283(.A(mai_mai_n311_), .B(mai_mai_n301_), .C(mai_mai_n278_), .D(mai_mai_n271_), .Y(mai_mai_n312_));
  NAi21      m0284(.An(m), .B(k), .Y(mai_mai_n313_));
  NO2        m0285(.A(mai_mai_n231_), .B(mai_mai_n313_), .Y(mai_mai_n314_));
  NAi41      m0286(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n315_));
  NO2        m0287(.A(mai_mai_n315_), .B(mai_mai_n153_), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n316_), .B(mai_mai_n314_), .Y(mai_mai_n317_));
  NO4        m0289(.A(i), .B(mai_mai_n153_), .C(mai_mai_n73_), .D(mai_mai_n75_), .Y(mai_mai_n318_));
  NA2        m0290(.A(e), .B(c), .Y(mai_mai_n319_));
  NOi21      m0291(.An(f), .B(h), .Y(mai_mai_n320_));
  NA2        m0292(.A(mai_mai_n320_), .B(mai_mai_n120_), .Y(mai_mai_n321_));
  NO2        m0293(.A(mai_mai_n321_), .B(mai_mai_n219_), .Y(mai_mai_n322_));
  NAi31      m0294(.An(d), .B(e), .C(b), .Y(mai_mai_n323_));
  NO2        m0295(.A(mai_mai_n134_), .B(mai_mai_n323_), .Y(mai_mai_n324_));
  NA2        m0296(.A(mai_mai_n324_), .B(mai_mai_n322_), .Y(mai_mai_n325_));
  NAi31      m0297(.An(mai_mai_n318_), .B(mai_mai_n325_), .C(mai_mai_n317_), .Y(mai_mai_n326_));
  NO4        m0298(.A(mai_mai_n315_), .B(mai_mai_n81_), .C(mai_mai_n72_), .D(mai_mai_n219_), .Y(mai_mai_n327_));
  NA2        m0299(.A(mai_mai_n252_), .B(mai_mai_n106_), .Y(mai_mai_n328_));
  OR2        m0300(.A(mai_mai_n328_), .B(mai_mai_n208_), .Y(mai_mai_n329_));
  NOi31      m0301(.An(l), .B(n), .C(m), .Y(mai_mai_n330_));
  NA2        m0302(.A(mai_mai_n330_), .B(mai_mai_n220_), .Y(mai_mai_n331_));
  NAi21      m0303(.An(mai_mai_n327_), .B(mai_mai_n329_), .Y(mai_mai_n332_));
  NAi32      m0304(.An(m), .Bn(j), .C(k), .Y(mai_mai_n333_));
  NAi41      m0305(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n334_));
  OAI210     m0306(.A0(mai_mai_n216_), .A1(mai_mai_n333_), .B0(mai_mai_n334_), .Y(mai_mai_n335_));
  NOi31      m0307(.An(j), .B(m), .C(k), .Y(mai_mai_n336_));
  NO2        m0308(.A(mai_mai_n127_), .B(mai_mai_n336_), .Y(mai_mai_n337_));
  AN3        m0309(.A(h), .B(g), .C(f), .Y(mai_mai_n338_));
  NAi31      m0310(.An(mai_mai_n337_), .B(mai_mai_n338_), .C(mai_mai_n335_), .Y(mai_mai_n339_));
  NAi32      m0311(.An(mai_mai_n1459_), .Bn(mai_mai_n205_), .C(mai_mai_n302_), .Y(mai_mai_n340_));
  NO2        m0312(.A(mai_mai_n295_), .B(mai_mai_n294_), .Y(mai_mai_n341_));
  NO2        m0313(.A(mai_mai_n222_), .B(g), .Y(mai_mai_n342_));
  NO2        m0314(.A(mai_mai_n159_), .B(mai_mai_n86_), .Y(mai_mai_n343_));
  AOI220     m0315(.A0(mai_mai_n343_), .A1(mai_mai_n342_), .B0(mai_mai_n249_), .B1(mai_mai_n341_), .Y(mai_mai_n344_));
  NA2        m0316(.A(mai_mai_n235_), .B(mai_mai_n81_), .Y(mai_mai_n345_));
  NA3        m0317(.A(mai_mai_n345_), .B(mai_mai_n338_), .C(mai_mai_n217_), .Y(mai_mai_n346_));
  NA4        m0318(.A(mai_mai_n346_), .B(mai_mai_n344_), .C(mai_mai_n340_), .D(mai_mai_n339_), .Y(mai_mai_n347_));
  NA3        m0319(.A(h), .B(g), .C(f), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n348_), .B(mai_mai_n77_), .Y(mai_mai_n349_));
  NA2        m0321(.A(mai_mai_n334_), .B(mai_mai_n216_), .Y(mai_mai_n350_));
  NA2        m0322(.A(h), .B(e), .Y(mai_mai_n351_));
  NO2        m0323(.A(mai_mai_n351_), .B(mai_mai_n41_), .Y(mai_mai_n352_));
  AOI220     m0324(.A0(mai_mai_n352_), .A1(mai_mai_n308_), .B0(mai_mai_n350_), .B1(mai_mai_n349_), .Y(mai_mai_n353_));
  NOi32      m0325(.An(j), .Bn(g), .C(i), .Y(mai_mai_n354_));
  NA3        m0326(.A(mai_mai_n354_), .B(mai_mai_n287_), .C(mai_mai_n115_), .Y(mai_mai_n355_));
  AO210      m0327(.A0(mai_mai_n113_), .A1(mai_mai_n32_), .B0(mai_mai_n355_), .Y(mai_mai_n356_));
  NOi32      m0328(.An(e), .Bn(b), .C(a), .Y(mai_mai_n357_));
  AN2        m0329(.A(l), .B(j), .Y(mai_mai_n358_));
  INV        m0330(.A(mai_mai_n313_), .Y(mai_mai_n359_));
  NO3        m0331(.A(mai_mai_n315_), .B(mai_mai_n72_), .C(mai_mai_n219_), .Y(mai_mai_n360_));
  NA3        m0332(.A(mai_mai_n213_), .B(mai_mai_n211_), .C(mai_mai_n35_), .Y(mai_mai_n361_));
  AOI220     m0333(.A0(mai_mai_n361_), .A1(mai_mai_n357_), .B0(mai_mai_n360_), .B1(mai_mai_n359_), .Y(mai_mai_n362_));
  NO2        m0334(.A(mai_mai_n323_), .B(n), .Y(mai_mai_n363_));
  NA2        m0335(.A(mai_mai_n212_), .B(k), .Y(mai_mai_n364_));
  NA4        m0336(.A(mai_mai_n207_), .B(mai_mai_n89_), .C(g), .D(mai_mai_n218_), .Y(mai_mai_n365_));
  INV        m0337(.A(mai_mai_n365_), .Y(mai_mai_n366_));
  NAi41      m0338(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n367_));
  NA2        m0339(.A(mai_mai_n51_), .B(mai_mai_n115_), .Y(mai_mai_n368_));
  NO2        m0340(.A(mai_mai_n368_), .B(mai_mai_n367_), .Y(mai_mai_n369_));
  AOI220     m0341(.A0(mai_mai_n369_), .A1(b), .B0(mai_mai_n366_), .B1(mai_mai_n363_), .Y(mai_mai_n370_));
  NA4        m0342(.A(mai_mai_n370_), .B(mai_mai_n362_), .C(mai_mai_n356_), .D(mai_mai_n353_), .Y(mai_mai_n371_));
  NO4        m0343(.A(mai_mai_n371_), .B(mai_mai_n347_), .C(mai_mai_n332_), .D(mai_mai_n326_), .Y(mai_mai_n372_));
  NA4        m0344(.A(mai_mai_n372_), .B(mai_mai_n312_), .C(mai_mai_n269_), .D(mai_mai_n204_), .Y(mai10));
  NA3        m0345(.A(m), .B(k), .C(i), .Y(mai_mai_n374_));
  NO3        m0346(.A(mai_mai_n374_), .B(j), .C(mai_mai_n219_), .Y(mai_mai_n375_));
  NOi21      m0347(.An(e), .B(f), .Y(mai_mai_n376_));
  NO4        m0348(.A(mai_mai_n154_), .B(mai_mai_n376_), .C(n), .D(mai_mai_n112_), .Y(mai_mai_n377_));
  NAi31      m0349(.An(b), .B(f), .C(c), .Y(mai_mai_n378_));
  INV        m0350(.A(mai_mai_n378_), .Y(mai_mai_n379_));
  NOi32      m0351(.An(k), .Bn(h), .C(j), .Y(mai_mai_n380_));
  NA2        m0352(.A(mai_mai_n380_), .B(mai_mai_n226_), .Y(mai_mai_n381_));
  NA2        m0353(.A(mai_mai_n164_), .B(mai_mai_n381_), .Y(mai_mai_n382_));
  AOI220     m0354(.A0(mai_mai_n382_), .A1(mai_mai_n379_), .B0(mai_mai_n377_), .B1(mai_mai_n375_), .Y(mai_mai_n383_));
  AN2        m0355(.A(j), .B(h), .Y(mai_mai_n384_));
  OR2        m0356(.A(m), .B(k), .Y(mai_mai_n385_));
  NO2        m0357(.A(mai_mai_n177_), .B(mai_mai_n385_), .Y(mai_mai_n386_));
  NA4        m0358(.A(n), .B(f), .C(c), .D(mai_mai_n118_), .Y(mai_mai_n387_));
  NOi21      m0359(.An(mai_mai_n386_), .B(mai_mai_n387_), .Y(mai_mai_n388_));
  NOi32      m0360(.An(d), .Bn(a), .C(c), .Y(mai_mai_n389_));
  NA2        m0361(.A(mai_mai_n389_), .B(mai_mai_n185_), .Y(mai_mai_n390_));
  NAi21      m0362(.An(i), .B(g), .Y(mai_mai_n391_));
  NAi31      m0363(.An(k), .B(m), .C(j), .Y(mai_mai_n392_));
  NO3        m0364(.A(mai_mai_n392_), .B(mai_mai_n391_), .C(n), .Y(mai_mai_n393_));
  NOi21      m0365(.An(mai_mai_n393_), .B(mai_mai_n390_), .Y(mai_mai_n394_));
  NO2        m0366(.A(mai_mai_n394_), .B(mai_mai_n388_), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n387_), .B(mai_mai_n295_), .Y(mai_mai_n396_));
  NA2        m0368(.A(mai_mai_n396_), .B(mai_mai_n220_), .Y(mai_mai_n397_));
  NA3        m0369(.A(mai_mai_n397_), .B(mai_mai_n395_), .C(mai_mai_n383_), .Y(mai_mai_n398_));
  NO2        m0370(.A(mai_mai_n59_), .B(mai_mai_n118_), .Y(mai_mai_n399_));
  NA2        m0371(.A(mai_mai_n252_), .B(mai_mai_n399_), .Y(mai_mai_n400_));
  INV        m0372(.A(e), .Y(mai_mai_n401_));
  NA2        m0373(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n402_));
  OAI220     m0374(.A0(mai_mai_n402_), .A1(mai_mai_n1460_), .B0(mai_mai_n208_), .B1(mai_mai_n401_), .Y(mai_mai_n403_));
  AN2        m0375(.A(g), .B(e), .Y(mai_mai_n404_));
  NA3        m0376(.A(mai_mai_n404_), .B(mai_mai_n207_), .C(i), .Y(mai_mai_n405_));
  OAI210     m0377(.A0(mai_mai_n91_), .A1(mai_mai_n401_), .B0(mai_mai_n405_), .Y(mai_mai_n406_));
  NO2        m0378(.A(mai_mai_n102_), .B(mai_mai_n401_), .Y(mai_mai_n407_));
  NO3        m0379(.A(mai_mai_n407_), .B(mai_mai_n406_), .C(mai_mai_n403_), .Y(mai_mai_n408_));
  NOi32      m0380(.An(h), .Bn(e), .C(g), .Y(mai_mai_n409_));
  NA3        m0381(.A(mai_mai_n409_), .B(mai_mai_n289_), .C(m), .Y(mai_mai_n410_));
  NOi21      m0382(.An(g), .B(h), .Y(mai_mai_n411_));
  AN3        m0383(.A(m), .B(l), .C(i), .Y(mai_mai_n412_));
  NA3        m0384(.A(mai_mai_n412_), .B(mai_mai_n411_), .C(e), .Y(mai_mai_n413_));
  AN3        m0385(.A(h), .B(g), .C(e), .Y(mai_mai_n414_));
  NA2        m0386(.A(mai_mai_n414_), .B(m), .Y(mai_mai_n415_));
  AN3        m0387(.A(mai_mai_n415_), .B(mai_mai_n413_), .C(mai_mai_n410_), .Y(mai_mai_n416_));
  AOI210     m0388(.A0(mai_mai_n416_), .A1(mai_mai_n408_), .B0(mai_mai_n400_), .Y(mai_mai_n417_));
  NA3        m0389(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n418_));
  NO2        m0390(.A(mai_mai_n418_), .B(mai_mai_n400_), .Y(mai_mai_n419_));
  NA3        m0391(.A(mai_mai_n389_), .B(mai_mai_n185_), .C(mai_mai_n86_), .Y(mai_mai_n420_));
  NAi31      m0392(.An(b), .B(c), .C(a), .Y(mai_mai_n421_));
  NO2        m0393(.A(mai_mai_n421_), .B(n), .Y(mai_mai_n422_));
  OAI210     m0394(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n423_));
  NO2        m0395(.A(mai_mai_n423_), .B(mai_mai_n150_), .Y(mai_mai_n424_));
  NA2        m0396(.A(mai_mai_n424_), .B(mai_mai_n422_), .Y(mai_mai_n425_));
  INV        m0397(.A(mai_mai_n425_), .Y(mai_mai_n426_));
  NO4        m0398(.A(mai_mai_n426_), .B(mai_mai_n419_), .C(mai_mai_n417_), .D(mai_mai_n398_), .Y(mai_mai_n427_));
  NA2        m0399(.A(i), .B(g), .Y(mai_mai_n428_));
  NO3        m0400(.A(mai_mai_n277_), .B(mai_mai_n428_), .C(c), .Y(mai_mai_n429_));
  NOi21      m0401(.An(a), .B(n), .Y(mai_mai_n430_));
  NA2        m0402(.A(d), .B(mai_mai_n430_), .Y(mai_mai_n431_));
  NA3        m0403(.A(i), .B(g), .C(f), .Y(mai_mai_n432_));
  OR2        m0404(.A(mai_mai_n432_), .B(mai_mai_n71_), .Y(mai_mai_n433_));
  NA3        m0405(.A(mai_mai_n412_), .B(mai_mai_n411_), .C(mai_mai_n185_), .Y(mai_mai_n434_));
  AOI210     m0406(.A0(mai_mai_n434_), .A1(mai_mai_n433_), .B0(mai_mai_n431_), .Y(mai_mai_n435_));
  AOI210     m0407(.A0(mai_mai_n429_), .A1(mai_mai_n288_), .B0(mai_mai_n435_), .Y(mai_mai_n436_));
  OR2        m0408(.A(n), .B(m), .Y(mai_mai_n437_));
  NO2        m0409(.A(mai_mai_n437_), .B(mai_mai_n155_), .Y(mai_mai_n438_));
  NO2        m0410(.A(mai_mai_n186_), .B(mai_mai_n150_), .Y(mai_mai_n439_));
  OAI210     m0411(.A0(mai_mai_n438_), .A1(mai_mai_n179_), .B0(mai_mai_n439_), .Y(mai_mai_n440_));
  INV        m0412(.A(mai_mai_n368_), .Y(mai_mai_n441_));
  NA3        m0413(.A(mai_mai_n441_), .B(mai_mai_n357_), .C(d), .Y(mai_mai_n442_));
  NO2        m0414(.A(mai_mai_n421_), .B(mai_mai_n49_), .Y(mai_mai_n443_));
  NO3        m0415(.A(mai_mai_n66_), .B(mai_mai_n114_), .C(e), .Y(mai_mai_n444_));
  NAi21      m0416(.An(k), .B(j), .Y(mai_mai_n445_));
  NA3        m0417(.A(i), .B(mai_mai_n444_), .C(mai_mai_n443_), .Y(mai_mai_n446_));
  NAi21      m0418(.An(e), .B(d), .Y(mai_mai_n447_));
  NO2        m0419(.A(mai_mai_n256_), .B(mai_mai_n218_), .Y(mai_mai_n448_));
  NA3        m0420(.A(mai_mai_n446_), .B(mai_mai_n442_), .C(mai_mai_n440_), .Y(mai_mai_n449_));
  NO2        m0421(.A(mai_mai_n331_), .B(mai_mai_n218_), .Y(mai_mai_n450_));
  NA2        m0422(.A(mai_mai_n450_), .B(d), .Y(mai_mai_n451_));
  NOi31      m0423(.An(n), .B(m), .C(k), .Y(mai_mai_n452_));
  AOI220     m0424(.A0(mai_mai_n452_), .A1(mai_mai_n384_), .B0(mai_mai_n226_), .B1(mai_mai_n50_), .Y(mai_mai_n453_));
  NAi31      m0425(.An(g), .B(f), .C(c), .Y(mai_mai_n454_));
  NA2        m0426(.A(mai_mai_n451_), .B(mai_mai_n307_), .Y(mai_mai_n455_));
  NOi41      m0427(.An(mai_mai_n436_), .B(mai_mai_n455_), .C(mai_mai_n449_), .D(mai_mai_n267_), .Y(mai_mai_n456_));
  NOi32      m0428(.An(c), .Bn(a), .C(b), .Y(mai_mai_n457_));
  NA2        m0429(.A(mai_mai_n457_), .B(mai_mai_n115_), .Y(mai_mai_n458_));
  INV        m0430(.A(mai_mai_n276_), .Y(mai_mai_n459_));
  AN2        m0431(.A(e), .B(d), .Y(mai_mai_n460_));
  NA2        m0432(.A(mai_mai_n460_), .B(mai_mai_n459_), .Y(mai_mai_n461_));
  NO2        m0433(.A(mai_mai_n133_), .B(mai_mai_n41_), .Y(mai_mai_n462_));
  NO2        m0434(.A(mai_mai_n66_), .B(e), .Y(mai_mai_n463_));
  AOI210     m0435(.A0(mai_mai_n462_), .A1(f), .B0(mai_mai_n463_), .Y(mai_mai_n464_));
  AOI210     m0436(.A0(mai_mai_n464_), .A1(mai_mai_n461_), .B0(mai_mai_n458_), .Y(mai_mai_n465_));
  NO2        m0437(.A(mai_mai_n214_), .B(mai_mai_n209_), .Y(mai_mai_n466_));
  NOi21      m0438(.An(a), .B(b), .Y(mai_mai_n467_));
  NA3        m0439(.A(e), .B(d), .C(c), .Y(mai_mai_n468_));
  NAi21      m0440(.An(mai_mai_n468_), .B(mai_mai_n467_), .Y(mai_mai_n469_));
  NO2        m0441(.A(mai_mai_n420_), .B(mai_mai_n208_), .Y(mai_mai_n470_));
  NOi21      m0442(.An(mai_mai_n469_), .B(mai_mai_n470_), .Y(mai_mai_n471_));
  AOI210     m0443(.A0(mai_mai_n270_), .A1(mai_mai_n466_), .B0(mai_mai_n471_), .Y(mai_mai_n472_));
  NO4        m0444(.A(mai_mai_n192_), .B(mai_mai_n105_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n473_));
  NA2        m0445(.A(mai_mai_n379_), .B(mai_mai_n156_), .Y(mai_mai_n474_));
  OR2        m0446(.A(k), .B(j), .Y(mai_mai_n475_));
  NA2        m0447(.A(l), .B(k), .Y(mai_mai_n476_));
  NA3        m0448(.A(mai_mai_n476_), .B(mai_mai_n475_), .C(mai_mai_n226_), .Y(mai_mai_n477_));
  AOI210     m0449(.A0(mai_mai_n235_), .A1(mai_mai_n333_), .B0(mai_mai_n86_), .Y(mai_mai_n478_));
  NOi21      m0450(.An(mai_mai_n477_), .B(mai_mai_n478_), .Y(mai_mai_n479_));
  NA3        m0451(.A(mai_mai_n279_), .B(mai_mai_n130_), .C(mai_mai_n128_), .Y(mai_mai_n480_));
  NA2        m0452(.A(mai_mai_n389_), .B(mai_mai_n115_), .Y(mai_mai_n481_));
  NO4        m0453(.A(mai_mai_n481_), .B(mai_mai_n97_), .C(mai_mai_n114_), .D(e), .Y(mai_mai_n482_));
  NO3        m0454(.A(mai_mai_n420_), .B(mai_mai_n94_), .C(mai_mai_n133_), .Y(mai_mai_n483_));
  NO4        m0455(.A(mai_mai_n483_), .B(mai_mai_n482_), .C(mai_mai_n480_), .D(mai_mai_n318_), .Y(mai_mai_n484_));
  NA2        m0456(.A(mai_mai_n484_), .B(mai_mai_n474_), .Y(mai_mai_n485_));
  NO4        m0457(.A(mai_mai_n485_), .B(mai_mai_n473_), .C(mai_mai_n472_), .D(mai_mai_n465_), .Y(mai_mai_n486_));
  NA2        m0458(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n487_));
  NOi21      m0459(.An(d), .B(e), .Y(mai_mai_n488_));
  NO2        m0460(.A(mai_mai_n192_), .B(mai_mai_n56_), .Y(mai_mai_n489_));
  NAi31      m0461(.An(j), .B(l), .C(i), .Y(mai_mai_n490_));
  OAI210     m0462(.A0(mai_mai_n490_), .A1(mai_mai_n134_), .B0(mai_mai_n105_), .Y(mai_mai_n491_));
  NA4        m0463(.A(mai_mai_n491_), .B(mai_mai_n489_), .C(mai_mai_n488_), .D(b), .Y(mai_mai_n492_));
  NO3        m0464(.A(mai_mai_n390_), .B(mai_mai_n1459_), .C(mai_mai_n205_), .Y(mai_mai_n493_));
  NO2        m0465(.A(mai_mai_n390_), .B(mai_mai_n368_), .Y(mai_mai_n494_));
  NO4        m0466(.A(mai_mai_n494_), .B(mai_mai_n493_), .C(mai_mai_n188_), .D(mai_mai_n304_), .Y(mai_mai_n495_));
  NA4        m0467(.A(mai_mai_n495_), .B(mai_mai_n492_), .C(mai_mai_n487_), .D(mai_mai_n245_), .Y(mai_mai_n496_));
  OAI210     m0468(.A0(mai_mai_n129_), .A1(mai_mai_n127_), .B0(n), .Y(mai_mai_n497_));
  NO2        m0469(.A(mai_mai_n497_), .B(mai_mai_n133_), .Y(mai_mai_n498_));
  OA210      m0470(.A0(mai_mai_n296_), .A1(mai_mai_n498_), .B0(mai_mai_n197_), .Y(mai_mai_n499_));
  XO2        m0471(.A(i), .B(h), .Y(mai_mai_n500_));
  NA3        m0472(.A(mai_mai_n500_), .B(mai_mai_n163_), .C(n), .Y(mai_mai_n501_));
  NAi41      m0473(.An(mai_mai_n296_), .B(mai_mai_n501_), .C(mai_mai_n453_), .D(mai_mai_n381_), .Y(mai_mai_n502_));
  NOi32      m0474(.An(mai_mai_n502_), .Bn(mai_mai_n463_), .C(mai_mai_n1465_), .Y(mai_mai_n503_));
  NAi31      m0475(.An(c), .B(f), .C(d), .Y(mai_mai_n504_));
  AOI210     m0476(.A0(mai_mai_n280_), .A1(mai_mai_n200_), .B0(mai_mai_n504_), .Y(mai_mai_n505_));
  NA3        m0477(.A(mai_mai_n377_), .B(m), .C(mai_mai_n99_), .Y(mai_mai_n506_));
  NO2        m0478(.A(mai_mai_n184_), .B(mai_mai_n504_), .Y(mai_mai_n507_));
  AOI210     m0479(.A0(mai_mai_n355_), .A1(mai_mai_n35_), .B0(mai_mai_n469_), .Y(mai_mai_n508_));
  NOi31      m0480(.An(mai_mai_n506_), .B(mai_mai_n508_), .C(mai_mai_n507_), .Y(mai_mai_n509_));
  AO220      m0481(.A0(mai_mai_n285_), .A1(mai_mai_n264_), .B0(mai_mai_n168_), .B1(mai_mai_n67_), .Y(mai_mai_n510_));
  NA3        m0482(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n511_));
  NO2        m0483(.A(mai_mai_n511_), .B(mai_mai_n431_), .Y(mai_mai_n512_));
  NO2        m0484(.A(mai_mai_n512_), .B(mai_mai_n292_), .Y(mai_mai_n513_));
  NAi41      m0485(.An(mai_mai_n510_), .B(mai_mai_n513_), .C(mai_mai_n509_), .D(mai_mai_n84_), .Y(mai_mai_n514_));
  NO4        m0486(.A(mai_mai_n514_), .B(mai_mai_n503_), .C(mai_mai_n499_), .D(mai_mai_n496_), .Y(mai_mai_n515_));
  NA4        m0487(.A(mai_mai_n515_), .B(mai_mai_n486_), .C(mai_mai_n456_), .D(mai_mai_n427_), .Y(mai11));
  NO2        m0488(.A(mai_mai_n73_), .B(f), .Y(mai_mai_n517_));
  NA2        m0489(.A(j), .B(g), .Y(mai_mai_n518_));
  NAi31      m0490(.An(i), .B(m), .C(l), .Y(mai_mai_n519_));
  NA3        m0491(.A(m), .B(k), .C(j), .Y(mai_mai_n520_));
  OAI220     m0492(.A0(mai_mai_n520_), .A1(mai_mai_n133_), .B0(mai_mai_n519_), .B1(mai_mai_n518_), .Y(mai_mai_n521_));
  NA2        m0493(.A(mai_mai_n521_), .B(mai_mai_n517_), .Y(mai_mai_n522_));
  NOi32      m0494(.An(e), .Bn(b), .C(f), .Y(mai_mai_n523_));
  NA2        m0495(.A(j), .B(mai_mai_n115_), .Y(mai_mai_n524_));
  NA2        m0496(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n525_));
  OAI220     m0497(.A0(mai_mai_n525_), .A1(mai_mai_n298_), .B0(mai_mai_n524_), .B1(mai_mai_n219_), .Y(mai_mai_n526_));
  NAi31      m0498(.An(d), .B(e), .C(a), .Y(mai_mai_n527_));
  NO2        m0499(.A(mai_mai_n527_), .B(n), .Y(mai_mai_n528_));
  AOI220     m0500(.A0(mai_mai_n528_), .A1(mai_mai_n103_), .B0(mai_mai_n526_), .B1(mai_mai_n523_), .Y(mai_mai_n529_));
  NAi41      m0501(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n530_));
  AN2        m0502(.A(mai_mai_n530_), .B(mai_mai_n367_), .Y(mai_mai_n531_));
  AOI210     m0503(.A0(mai_mai_n531_), .A1(mai_mai_n390_), .B0(mai_mai_n272_), .Y(mai_mai_n532_));
  NA2        m0504(.A(j), .B(i), .Y(mai_mai_n533_));
  NAi31      m0505(.An(n), .B(m), .C(k), .Y(mai_mai_n534_));
  NO3        m0506(.A(mai_mai_n534_), .B(mai_mai_n533_), .C(mai_mai_n114_), .Y(mai_mai_n535_));
  NO4        m0507(.A(n), .B(d), .C(mai_mai_n118_), .D(a), .Y(mai_mai_n536_));
  OR2        m0508(.A(n), .B(c), .Y(mai_mai_n537_));
  NO2        m0509(.A(mai_mai_n537_), .B(mai_mai_n152_), .Y(mai_mai_n538_));
  NO2        m0510(.A(mai_mai_n538_), .B(mai_mai_n536_), .Y(mai_mai_n539_));
  NOi32      m0511(.An(g), .Bn(f), .C(i), .Y(mai_mai_n540_));
  AOI220     m0512(.A0(mai_mai_n540_), .A1(mai_mai_n101_), .B0(mai_mai_n521_), .B1(f), .Y(mai_mai_n541_));
  NO2        m0513(.A(mai_mai_n276_), .B(mai_mai_n49_), .Y(mai_mai_n542_));
  NO2        m0514(.A(mai_mai_n541_), .B(mai_mai_n539_), .Y(mai_mai_n543_));
  AOI210     m0515(.A0(mai_mai_n535_), .A1(mai_mai_n532_), .B0(mai_mai_n543_), .Y(mai_mai_n544_));
  NA2        m0516(.A(mai_mai_n143_), .B(mai_mai_n34_), .Y(mai_mai_n545_));
  OAI220     m0517(.A0(mai_mai_n545_), .A1(m), .B0(mai_mai_n525_), .B1(mai_mai_n235_), .Y(mai_mai_n546_));
  NOi41      m0518(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n547_));
  NAi32      m0519(.An(e), .Bn(b), .C(c), .Y(mai_mai_n548_));
  OR2        m0520(.A(mai_mai_n548_), .B(mai_mai_n86_), .Y(mai_mai_n549_));
  AN2        m0521(.A(mai_mai_n334_), .B(mai_mai_n315_), .Y(mai_mai_n550_));
  NA2        m0522(.A(mai_mai_n550_), .B(mai_mai_n549_), .Y(mai_mai_n551_));
  OA210      m0523(.A0(mai_mai_n551_), .A1(mai_mai_n547_), .B0(mai_mai_n546_), .Y(mai_mai_n552_));
  OAI220     m0524(.A0(mai_mai_n392_), .A1(mai_mai_n391_), .B0(mai_mai_n519_), .B1(mai_mai_n518_), .Y(mai_mai_n553_));
  NAi31      m0525(.An(d), .B(c), .C(a), .Y(mai_mai_n554_));
  NO2        m0526(.A(mai_mai_n554_), .B(n), .Y(mai_mai_n555_));
  NA3        m0527(.A(mai_mai_n555_), .B(mai_mai_n553_), .C(e), .Y(mai_mai_n556_));
  NO3        m0528(.A(mai_mai_n62_), .B(mai_mai_n49_), .C(mai_mai_n219_), .Y(mai_mai_n557_));
  NO2        m0529(.A(mai_mai_n232_), .B(mai_mai_n112_), .Y(mai_mai_n558_));
  OAI210     m0530(.A0(mai_mai_n557_), .A1(mai_mai_n393_), .B0(mai_mai_n558_), .Y(mai_mai_n559_));
  NA2        m0531(.A(mai_mai_n559_), .B(mai_mai_n556_), .Y(mai_mai_n560_));
  NO2        m0532(.A(mai_mai_n277_), .B(n), .Y(mai_mai_n561_));
  NO2        m0533(.A(mai_mai_n422_), .B(mai_mai_n561_), .Y(mai_mai_n562_));
  NA2        m0534(.A(mai_mai_n553_), .B(f), .Y(mai_mai_n563_));
  NAi32      m0535(.An(d), .Bn(a), .C(b), .Y(mai_mai_n564_));
  NO2        m0536(.A(mai_mai_n564_), .B(mai_mai_n49_), .Y(mai_mai_n565_));
  NA2        m0537(.A(h), .B(f), .Y(mai_mai_n566_));
  NO2        m0538(.A(mai_mai_n566_), .B(mai_mai_n97_), .Y(mai_mai_n567_));
  NO3        m0539(.A(mai_mai_n180_), .B(mai_mai_n177_), .C(g), .Y(mai_mai_n568_));
  AOI220     m0540(.A0(mai_mai_n568_), .A1(mai_mai_n58_), .B0(mai_mai_n567_), .B1(mai_mai_n565_), .Y(mai_mai_n569_));
  OAI210     m0541(.A0(mai_mai_n563_), .A1(mai_mai_n562_), .B0(mai_mai_n569_), .Y(mai_mai_n570_));
  AN3        m0542(.A(j), .B(h), .C(g), .Y(mai_mai_n571_));
  NO2        m0543(.A(mai_mai_n149_), .B(c), .Y(mai_mai_n572_));
  NA3        m0544(.A(mai_mai_n572_), .B(mai_mai_n571_), .C(mai_mai_n452_), .Y(mai_mai_n573_));
  NA3        m0545(.A(f), .B(d), .C(b), .Y(mai_mai_n574_));
  NO4        m0546(.A(mai_mai_n574_), .B(mai_mai_n180_), .C(mai_mai_n177_), .D(g), .Y(mai_mai_n575_));
  NAi21      m0547(.An(mai_mai_n575_), .B(mai_mai_n573_), .Y(mai_mai_n576_));
  NO4        m0548(.A(mai_mai_n576_), .B(mai_mai_n570_), .C(mai_mai_n560_), .D(mai_mai_n552_), .Y(mai_mai_n577_));
  AN4        m0549(.A(mai_mai_n577_), .B(mai_mai_n544_), .C(mai_mai_n529_), .D(mai_mai_n522_), .Y(mai_mai_n578_));
  INV        m0550(.A(k), .Y(mai_mai_n579_));
  NA4        m0551(.A(mai_mai_n389_), .B(mai_mai_n411_), .C(mai_mai_n185_), .D(mai_mai_n115_), .Y(mai_mai_n580_));
  NAi32      m0552(.An(h), .Bn(f), .C(g), .Y(mai_mai_n581_));
  NAi41      m0553(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n582_));
  OAI210     m0554(.A0(mai_mai_n527_), .A1(n), .B0(mai_mai_n582_), .Y(mai_mai_n583_));
  NA2        m0555(.A(mai_mai_n583_), .B(m), .Y(mai_mai_n584_));
  NAi31      m0556(.An(h), .B(g), .C(f), .Y(mai_mai_n585_));
  OR3        m0557(.A(mai_mai_n585_), .B(mai_mai_n277_), .C(mai_mai_n49_), .Y(mai_mai_n586_));
  NA4        m0558(.A(mai_mai_n411_), .B(mai_mai_n122_), .C(mai_mai_n115_), .D(e), .Y(mai_mai_n587_));
  AN2        m0559(.A(mai_mai_n587_), .B(mai_mai_n586_), .Y(mai_mai_n588_));
  OA210      m0560(.A0(mai_mai_n584_), .A1(mai_mai_n581_), .B0(mai_mai_n588_), .Y(mai_mai_n589_));
  NO3        m0561(.A(mai_mai_n581_), .B(mai_mai_n73_), .C(mai_mai_n75_), .Y(mai_mai_n590_));
  NO4        m0562(.A(mai_mai_n585_), .B(mai_mai_n537_), .C(mai_mai_n152_), .D(mai_mai_n75_), .Y(mai_mai_n591_));
  OR2        m0563(.A(mai_mai_n591_), .B(mai_mai_n590_), .Y(mai_mai_n592_));
  NAi31      m0564(.An(mai_mai_n592_), .B(mai_mai_n589_), .C(mai_mai_n580_), .Y(mai_mai_n593_));
  NAi31      m0565(.An(f), .B(h), .C(g), .Y(mai_mai_n594_));
  NO4        m0566(.A(k), .B(mai_mai_n594_), .C(mai_mai_n73_), .D(mai_mai_n75_), .Y(mai_mai_n595_));
  NOi41      m0567(.An(b), .B(mai_mai_n348_), .C(mai_mai_n69_), .D(mai_mai_n119_), .Y(mai_mai_n596_));
  OR2        m0568(.A(mai_mai_n596_), .B(mai_mai_n595_), .Y(mai_mai_n597_));
  NOi32      m0569(.An(d), .Bn(a), .C(e), .Y(mai_mai_n598_));
  NA2        m0570(.A(mai_mai_n598_), .B(mai_mai_n115_), .Y(mai_mai_n599_));
  NO2        m0571(.A(n), .B(c), .Y(mai_mai_n600_));
  NA3        m0572(.A(mai_mai_n600_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n601_));
  NAi32      m0573(.An(n), .Bn(f), .C(m), .Y(mai_mai_n602_));
  NA3        m0574(.A(mai_mai_n602_), .B(mai_mai_n601_), .C(mai_mai_n599_), .Y(mai_mai_n603_));
  NOi32      m0575(.An(e), .Bn(a), .C(d), .Y(mai_mai_n604_));
  AOI210     m0576(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n604_), .Y(mai_mai_n605_));
  AOI210     m0577(.A0(mai_mai_n605_), .A1(mai_mai_n218_), .B0(mai_mai_n545_), .Y(mai_mai_n606_));
  AOI210     m0578(.A0(mai_mai_n606_), .A1(mai_mai_n603_), .B0(mai_mai_n597_), .Y(mai_mai_n607_));
  OAI210     m0579(.A0(mai_mai_n251_), .A1(mai_mai_n89_), .B0(mai_mai_n607_), .Y(mai_mai_n608_));
  AOI210     m0580(.A0(mai_mai_n593_), .A1(mai_mai_n579_), .B0(mai_mai_n608_), .Y(mai_mai_n609_));
  NO3        m0581(.A(mai_mai_n313_), .B(mai_mai_n61_), .C(n), .Y(mai_mai_n610_));
  NA3        m0582(.A(mai_mai_n504_), .B(mai_mai_n175_), .C(mai_mai_n174_), .Y(mai_mai_n611_));
  NA2        m0583(.A(mai_mai_n454_), .B(mai_mai_n232_), .Y(mai_mai_n612_));
  OR2        m0584(.A(mai_mai_n612_), .B(mai_mai_n611_), .Y(mai_mai_n613_));
  NA2        m0585(.A(mai_mai_n76_), .B(mai_mai_n115_), .Y(mai_mai_n614_));
  AOI220     m0586(.A0(mai_mai_n115_), .A1(mai_mai_n532_), .B0(mai_mai_n613_), .B1(mai_mai_n610_), .Y(mai_mai_n615_));
  NO2        m0587(.A(mai_mai_n615_), .B(mai_mai_n89_), .Y(mai_mai_n616_));
  NA3        m0588(.A(mai_mai_n547_), .B(mai_mai_n336_), .C(mai_mai_n46_), .Y(mai_mai_n617_));
  NOi32      m0589(.An(e), .Bn(c), .C(f), .Y(mai_mai_n618_));
  INV        m0590(.A(mai_mai_n216_), .Y(mai_mai_n619_));
  AOI220     m0591(.A0(mai_mai_n619_), .A1(mai_mai_n386_), .B0(mai_mai_n618_), .B1(mai_mai_n179_), .Y(mai_mai_n620_));
  NA3        m0592(.A(mai_mai_n620_), .B(mai_mai_n617_), .C(mai_mai_n182_), .Y(mai_mai_n621_));
  AOI210     m0593(.A0(mai_mai_n531_), .A1(mai_mai_n390_), .B0(mai_mai_n297_), .Y(mai_mai_n622_));
  NA2        m0594(.A(mai_mai_n622_), .B(mai_mai_n265_), .Y(mai_mai_n623_));
  NAi21      m0595(.An(k), .B(h), .Y(mai_mai_n624_));
  NO2        m0596(.A(mai_mai_n624_), .B(mai_mai_n263_), .Y(mai_mai_n625_));
  NA2        m0597(.A(mai_mai_n625_), .B(j), .Y(mai_mai_n626_));
  OR2        m0598(.A(mai_mai_n626_), .B(mai_mai_n584_), .Y(mai_mai_n627_));
  NOi31      m0599(.An(m), .B(n), .C(k), .Y(mai_mai_n628_));
  NA2        m0600(.A(j), .B(mai_mai_n628_), .Y(mai_mai_n629_));
  AOI210     m0601(.A0(mai_mai_n390_), .A1(mai_mai_n367_), .B0(mai_mai_n297_), .Y(mai_mai_n630_));
  NAi21      m0602(.An(mai_mai_n629_), .B(mai_mai_n630_), .Y(mai_mai_n631_));
  NO2        m0603(.A(mai_mai_n277_), .B(mai_mai_n49_), .Y(mai_mai_n632_));
  NO2        m0604(.A(k), .B(mai_mai_n594_), .Y(mai_mai_n633_));
  NO2        m0605(.A(mai_mai_n527_), .B(mai_mai_n49_), .Y(mai_mai_n634_));
  AOI220     m0606(.A0(mai_mai_n634_), .A1(mai_mai_n633_), .B0(mai_mai_n632_), .B1(mai_mai_n567_), .Y(mai_mai_n635_));
  NA4        m0607(.A(mai_mai_n635_), .B(mai_mai_n631_), .C(mai_mai_n627_), .D(mai_mai_n623_), .Y(mai_mai_n636_));
  NA2        m0608(.A(mai_mai_n110_), .B(mai_mai_n36_), .Y(mai_mai_n637_));
  NO2        m0609(.A(k), .B(mai_mai_n219_), .Y(mai_mai_n638_));
  NO2        m0610(.A(mai_mai_n523_), .B(mai_mai_n357_), .Y(mai_mai_n639_));
  NO2        m0611(.A(mai_mai_n639_), .B(n), .Y(mai_mai_n640_));
  NAi31      m0612(.An(mai_mai_n637_), .B(mai_mai_n640_), .C(mai_mai_n638_), .Y(mai_mai_n641_));
  NO2        m0613(.A(mai_mai_n525_), .B(mai_mai_n180_), .Y(mai_mai_n642_));
  NA2        m0614(.A(mai_mai_n500_), .B(mai_mai_n163_), .Y(mai_mai_n643_));
  NO3        m0615(.A(mai_mai_n387_), .B(mai_mai_n643_), .C(mai_mai_n89_), .Y(mai_mai_n644_));
  AOI210     m0616(.A0(c), .A1(mai_mai_n642_), .B0(mai_mai_n644_), .Y(mai_mai_n645_));
  AN3        m0617(.A(f), .B(d), .C(b), .Y(mai_mai_n646_));
  NA3        m0618(.A(mai_mai_n500_), .B(mai_mai_n163_), .C(mai_mai_n219_), .Y(mai_mai_n647_));
  NO2        m0619(.A(mai_mai_n234_), .B(mai_mai_n647_), .Y(mai_mai_n648_));
  NAi31      m0620(.An(m), .B(n), .C(k), .Y(mai_mai_n649_));
  OR2        m0621(.A(mai_mai_n137_), .B(mai_mai_n61_), .Y(mai_mai_n650_));
  OAI210     m0622(.A0(mai_mai_n650_), .A1(mai_mai_n649_), .B0(mai_mai_n253_), .Y(mai_mai_n651_));
  OAI210     m0623(.A0(mai_mai_n651_), .A1(mai_mai_n648_), .B0(j), .Y(mai_mai_n652_));
  NA3        m0624(.A(mai_mai_n652_), .B(mai_mai_n645_), .C(mai_mai_n641_), .Y(mai_mai_n653_));
  NO4        m0625(.A(mai_mai_n653_), .B(mai_mai_n636_), .C(mai_mai_n621_), .D(mai_mai_n616_), .Y(mai_mai_n654_));
  NA2        m0626(.A(mai_mai_n377_), .B(h), .Y(mai_mai_n655_));
  NAi31      m0627(.An(g), .B(h), .C(f), .Y(mai_mai_n656_));
  OR3        m0628(.A(mai_mai_n656_), .B(mai_mai_n277_), .C(n), .Y(mai_mai_n657_));
  OA210      m0629(.A0(mai_mai_n527_), .A1(n), .B0(mai_mai_n582_), .Y(mai_mai_n658_));
  NA3        m0630(.A(mai_mai_n409_), .B(mai_mai_n122_), .C(mai_mai_n86_), .Y(mai_mai_n659_));
  OAI210     m0631(.A0(mai_mai_n658_), .A1(mai_mai_n93_), .B0(mai_mai_n659_), .Y(mai_mai_n660_));
  NOi21      m0632(.An(mai_mai_n657_), .B(mai_mai_n660_), .Y(mai_mai_n661_));
  AOI210     m0633(.A0(mai_mai_n661_), .A1(mai_mai_n655_), .B0(mai_mai_n520_), .Y(mai_mai_n662_));
  OR2        m0634(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n663_));
  NA2        m0635(.A(b), .B(mai_mai_n338_), .Y(mai_mai_n664_));
  OA220      m0636(.A0(mai_mai_n629_), .A1(mai_mai_n664_), .B0(mai_mai_n626_), .B1(mai_mai_n663_), .Y(mai_mai_n665_));
  NA3        m0637(.A(mai_mai_n517_), .B(mai_mai_n101_), .C(mai_mai_n100_), .Y(mai_mai_n666_));
  NA2        m0638(.A(h), .B(mai_mai_n37_), .Y(mai_mai_n667_));
  NA2        m0639(.A(mai_mai_n101_), .B(mai_mai_n46_), .Y(mai_mai_n668_));
  OAI220     m0640(.A0(mai_mai_n668_), .A1(mai_mai_n328_), .B0(mai_mai_n667_), .B1(mai_mai_n458_), .Y(mai_mai_n669_));
  AOI210     m0641(.A0(mai_mai_n564_), .A1(mai_mai_n421_), .B0(mai_mai_n49_), .Y(mai_mai_n670_));
  OAI220     m0642(.A0(mai_mai_n585_), .A1(k), .B0(mai_mai_n321_), .B1(mai_mai_n518_), .Y(mai_mai_n671_));
  AOI210     m0643(.A0(mai_mai_n671_), .A1(mai_mai_n670_), .B0(mai_mai_n669_), .Y(mai_mai_n672_));
  NA3        m0644(.A(mai_mai_n672_), .B(mai_mai_n666_), .C(mai_mai_n665_), .Y(mai_mai_n673_));
  NO2        m0645(.A(mai_mai_n255_), .B(f), .Y(mai_mai_n674_));
  INV        m0646(.A(mai_mai_n61_), .Y(mai_mai_n675_));
  NO3        m0647(.A(mai_mai_n675_), .B(mai_mai_n674_), .C(mai_mai_n34_), .Y(mai_mai_n676_));
  NA2        m0648(.A(mai_mai_n324_), .B(mai_mai_n143_), .Y(mai_mai_n677_));
  NA2        m0649(.A(mai_mai_n134_), .B(mai_mai_n49_), .Y(mai_mai_n678_));
  AOI220     m0650(.A0(mai_mai_n678_), .A1(mai_mai_n523_), .B0(mai_mai_n357_), .B1(mai_mai_n115_), .Y(mai_mai_n679_));
  OA220      m0651(.A0(mai_mai_n679_), .A1(mai_mai_n545_), .B0(mai_mai_n355_), .B1(mai_mai_n113_), .Y(mai_mai_n680_));
  OAI210     m0652(.A0(mai_mai_n677_), .A1(mai_mai_n676_), .B0(mai_mai_n680_), .Y(mai_mai_n681_));
  NA3        m0653(.A(mai_mai_n196_), .B(mai_mai_n257_), .C(j), .Y(mai_mai_n682_));
  NO3        m0654(.A(mai_mai_n454_), .B(mai_mai_n177_), .C(i), .Y(mai_mai_n683_));
  NA2        m0655(.A(mai_mai_n457_), .B(mai_mai_n86_), .Y(mai_mai_n684_));
  NO4        m0656(.A(mai_mai_n520_), .B(mai_mai_n684_), .C(mai_mai_n133_), .D(mai_mai_n218_), .Y(mai_mai_n685_));
  INV        m0657(.A(mai_mai_n685_), .Y(mai_mai_n686_));
  NA4        m0658(.A(mai_mai_n686_), .B(mai_mai_n682_), .C(mai_mai_n506_), .D(mai_mai_n395_), .Y(mai_mai_n687_));
  NO4        m0659(.A(mai_mai_n687_), .B(mai_mai_n681_), .C(mai_mai_n673_), .D(mai_mai_n662_), .Y(mai_mai_n688_));
  NA4        m0660(.A(mai_mai_n688_), .B(mai_mai_n654_), .C(mai_mai_n609_), .D(mai_mai_n578_), .Y(mai08));
  NO2        m0661(.A(k), .B(h), .Y(mai_mai_n690_));
  AO210      m0662(.A0(mai_mai_n255_), .A1(mai_mai_n445_), .B0(mai_mai_n690_), .Y(mai_mai_n691_));
  NO2        m0663(.A(mai_mai_n691_), .B(mai_mai_n295_), .Y(mai_mai_n692_));
  NA2        m0664(.A(mai_mai_n618_), .B(mai_mai_n86_), .Y(mai_mai_n693_));
  NA2        m0665(.A(mai_mai_n693_), .B(mai_mai_n454_), .Y(mai_mai_n694_));
  AOI210     m0666(.A0(mai_mai_n694_), .A1(mai_mai_n692_), .B0(mai_mai_n483_), .Y(mai_mai_n695_));
  NO2        m0667(.A(n), .B(mai_mai_n57_), .Y(mai_mai_n696_));
  NO4        m0668(.A(mai_mai_n374_), .B(mai_mai_n114_), .C(j), .D(mai_mai_n219_), .Y(mai_mai_n697_));
  OAI210     m0669(.A0(mai_mai_n574_), .A1(mai_mai_n86_), .B0(mai_mai_n234_), .Y(mai_mai_n698_));
  AOI220     m0670(.A0(mai_mai_n698_), .A1(mai_mai_n342_), .B0(mai_mai_n697_), .B1(mai_mai_n696_), .Y(mai_mai_n699_));
  AOI210     m0671(.A0(mai_mai_n574_), .A1(mai_mai_n159_), .B0(mai_mai_n86_), .Y(mai_mai_n700_));
  NA4        m0672(.A(mai_mai_n221_), .B(mai_mai_n143_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n701_));
  AN2        m0673(.A(l), .B(k), .Y(mai_mai_n702_));
  NA4        m0674(.A(mai_mai_n702_), .B(mai_mai_n110_), .C(mai_mai_n75_), .D(mai_mai_n219_), .Y(mai_mai_n703_));
  OAI210     m0675(.A0(mai_mai_n701_), .A1(g), .B0(mai_mai_n703_), .Y(mai_mai_n704_));
  NA2        m0676(.A(mai_mai_n704_), .B(mai_mai_n700_), .Y(mai_mai_n705_));
  NA4        m0677(.A(mai_mai_n705_), .B(mai_mai_n699_), .C(mai_mai_n695_), .D(mai_mai_n344_), .Y(mai_mai_n706_));
  AN2        m0678(.A(mai_mai_n528_), .B(mai_mai_n98_), .Y(mai_mai_n707_));
  NO4        m0679(.A(mai_mai_n177_), .B(mai_mai_n385_), .C(mai_mai_n114_), .D(g), .Y(mai_mai_n708_));
  AOI210     m0680(.A0(mai_mai_n708_), .A1(mai_mai_n698_), .B0(mai_mai_n512_), .Y(mai_mai_n709_));
  NO2        m0681(.A(mai_mai_n38_), .B(mai_mai_n218_), .Y(mai_mai_n710_));
  AOI220     m0682(.A0(mai_mai_n619_), .A1(mai_mai_n341_), .B0(mai_mai_n710_), .B1(mai_mai_n561_), .Y(mai_mai_n711_));
  NAi31      m0683(.An(mai_mai_n707_), .B(mai_mai_n711_), .C(mai_mai_n709_), .Y(mai_mai_n712_));
  NO2        m0684(.A(mai_mai_n531_), .B(mai_mai_n35_), .Y(mai_mai_n713_));
  OAI210     m0685(.A0(mai_mai_n548_), .A1(mai_mai_n47_), .B0(mai_mai_n650_), .Y(mai_mai_n714_));
  NO2        m0686(.A(mai_mai_n476_), .B(mai_mai_n134_), .Y(mai_mai_n715_));
  AOI210     m0687(.A0(mai_mai_n715_), .A1(mai_mai_n714_), .B0(mai_mai_n713_), .Y(mai_mai_n716_));
  NO3        m0688(.A(mai_mai_n313_), .B(mai_mai_n133_), .C(mai_mai_n41_), .Y(mai_mai_n717_));
  NAi21      m0689(.An(mai_mai_n717_), .B(mai_mai_n703_), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n718_), .B(mai_mai_n78_), .Y(mai_mai_n719_));
  OAI210     m0691(.A0(mai_mai_n716_), .A1(mai_mai_n89_), .B0(mai_mai_n719_), .Y(mai_mai_n720_));
  NA2        m0692(.A(mai_mai_n357_), .B(mai_mai_n43_), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n702_), .B(mai_mai_n226_), .Y(mai_mai_n722_));
  NO2        m0694(.A(mai_mai_n722_), .B(mai_mai_n323_), .Y(mai_mai_n723_));
  AOI210     m0695(.A0(mai_mai_n723_), .A1(mai_mai_n674_), .B0(mai_mai_n482_), .Y(mai_mai_n724_));
  NA3        m0696(.A(m), .B(l), .C(k), .Y(mai_mai_n725_));
  AOI210     m0697(.A0(mai_mai_n659_), .A1(mai_mai_n657_), .B0(mai_mai_n725_), .Y(mai_mai_n726_));
  NO2        m0698(.A(mai_mai_n530_), .B(mai_mai_n272_), .Y(mai_mai_n727_));
  NOi21      m0699(.An(mai_mai_n727_), .B(mai_mai_n524_), .Y(mai_mai_n728_));
  NA4        m0700(.A(mai_mai_n115_), .B(l), .C(k), .D(mai_mai_n89_), .Y(mai_mai_n729_));
  NA3        m0701(.A(mai_mai_n122_), .B(mai_mai_n404_), .C(i), .Y(mai_mai_n730_));
  NO2        m0702(.A(mai_mai_n730_), .B(mai_mai_n729_), .Y(mai_mai_n731_));
  NO3        m0703(.A(mai_mai_n731_), .B(mai_mai_n728_), .C(mai_mai_n726_), .Y(mai_mai_n732_));
  NA3        m0704(.A(mai_mai_n732_), .B(mai_mai_n724_), .C(mai_mai_n721_), .Y(mai_mai_n733_));
  NO4        m0705(.A(mai_mai_n733_), .B(mai_mai_n720_), .C(mai_mai_n712_), .D(mai_mai_n706_), .Y(mai_mai_n734_));
  NA2        m0706(.A(mai_mai_n619_), .B(mai_mai_n386_), .Y(mai_mai_n735_));
  NA2        m0707(.A(mai_mai_n634_), .B(g), .Y(mai_mai_n736_));
  AO210      m0708(.A0(mai_mai_n736_), .A1(mai_mai_n586_), .B0(mai_mai_n533_), .Y(mai_mai_n737_));
  NO3        m0709(.A(mai_mai_n390_), .B(mai_mai_n518_), .C(h), .Y(mai_mai_n738_));
  AOI210     m0710(.A0(mai_mai_n738_), .A1(mai_mai_n115_), .B0(mai_mai_n494_), .Y(mai_mai_n739_));
  NA4        m0711(.A(mai_mai_n739_), .B(mai_mai_n737_), .C(mai_mai_n735_), .D(mai_mai_n254_), .Y(mai_mai_n740_));
  NA2        m0712(.A(mai_mai_n702_), .B(mai_mai_n75_), .Y(mai_mai_n741_));
  NOi21      m0713(.An(h), .B(j), .Y(mai_mai_n742_));
  NA2        m0714(.A(mai_mai_n742_), .B(f), .Y(mai_mai_n743_));
  NO2        m0715(.A(mai_mai_n743_), .B(mai_mai_n248_), .Y(mai_mai_n744_));
  NO2        m0716(.A(mai_mai_n744_), .B(mai_mai_n683_), .Y(mai_mai_n745_));
  OAI220     m0717(.A0(mai_mai_n745_), .A1(mai_mai_n741_), .B0(mai_mai_n588_), .B1(mai_mai_n62_), .Y(mai_mai_n746_));
  AOI210     m0718(.A0(mai_mai_n740_), .A1(l), .B0(mai_mai_n746_), .Y(mai_mai_n747_));
  NO2        m0719(.A(j), .B(i), .Y(mai_mai_n748_));
  NA3        m0720(.A(mai_mai_n748_), .B(mai_mai_n82_), .C(l), .Y(mai_mai_n749_));
  NA2        m0721(.A(mai_mai_n748_), .B(mai_mai_n33_), .Y(mai_mai_n750_));
  NA2        m0722(.A(mai_mai_n414_), .B(mai_mai_n122_), .Y(mai_mai_n751_));
  OA220      m0723(.A0(mai_mai_n751_), .A1(mai_mai_n750_), .B0(mai_mai_n749_), .B1(mai_mai_n584_), .Y(mai_mai_n752_));
  NO3        m0724(.A(mai_mai_n154_), .B(mai_mai_n49_), .C(mai_mai_n112_), .Y(mai_mai_n753_));
  NO3        m0725(.A(mai_mai_n537_), .B(mai_mai_n152_), .C(mai_mai_n75_), .Y(mai_mai_n754_));
  NO3        m0726(.A(mai_mai_n476_), .B(mai_mai_n432_), .C(j), .Y(mai_mai_n755_));
  OAI210     m0727(.A0(mai_mai_n754_), .A1(mai_mai_n753_), .B0(mai_mai_n755_), .Y(mai_mai_n756_));
  OAI210     m0728(.A0(mai_mai_n736_), .A1(mai_mai_n62_), .B0(mai_mai_n756_), .Y(mai_mai_n757_));
  NA2        m0729(.A(k), .B(j), .Y(mai_mai_n758_));
  NO3        m0730(.A(mai_mai_n295_), .B(mai_mai_n758_), .C(mai_mai_n40_), .Y(mai_mai_n759_));
  AOI210     m0731(.A0(mai_mai_n523_), .A1(n), .B0(mai_mai_n547_), .Y(mai_mai_n760_));
  NA2        m0732(.A(mai_mai_n760_), .B(mai_mai_n550_), .Y(mai_mai_n761_));
  AN3        m0733(.A(mai_mai_n761_), .B(mai_mai_n759_), .C(mai_mai_n100_), .Y(mai_mai_n762_));
  NO3        m0734(.A(mai_mai_n177_), .B(mai_mai_n385_), .C(mai_mai_n114_), .Y(mai_mai_n763_));
  AOI220     m0735(.A0(mai_mai_n763_), .A1(mai_mai_n249_), .B0(mai_mai_n612_), .B1(mai_mai_n306_), .Y(mai_mai_n764_));
  NAi31      m0736(.An(mai_mai_n605_), .B(mai_mai_n95_), .C(mai_mai_n86_), .Y(mai_mai_n765_));
  NA2        m0737(.A(mai_mai_n765_), .B(mai_mai_n764_), .Y(mai_mai_n766_));
  NO2        m0738(.A(mai_mai_n295_), .B(mai_mai_n138_), .Y(mai_mai_n767_));
  AOI220     m0739(.A0(mai_mai_n767_), .A1(mai_mai_n619_), .B0(mai_mai_n717_), .B1(mai_mai_n700_), .Y(mai_mai_n768_));
  NO2        m0740(.A(mai_mai_n725_), .B(mai_mai_n93_), .Y(mai_mai_n769_));
  NA2        m0741(.A(mai_mai_n769_), .B(mai_mai_n583_), .Y(mai_mai_n770_));
  NO2        m0742(.A(mai_mai_n585_), .B(mai_mai_n119_), .Y(mai_mai_n771_));
  OAI210     m0743(.A0(mai_mai_n771_), .A1(mai_mai_n755_), .B0(mai_mai_n670_), .Y(mai_mai_n772_));
  NA3        m0744(.A(mai_mai_n772_), .B(mai_mai_n770_), .C(mai_mai_n768_), .Y(mai_mai_n773_));
  OR4        m0745(.A(mai_mai_n773_), .B(mai_mai_n766_), .C(mai_mai_n762_), .D(mai_mai_n757_), .Y(mai_mai_n774_));
  NA3        m0746(.A(mai_mai_n760_), .B(mai_mai_n550_), .C(mai_mai_n549_), .Y(mai_mai_n775_));
  NA4        m0747(.A(mai_mai_n775_), .B(mai_mai_n221_), .C(mai_mai_n445_), .D(mai_mai_n34_), .Y(mai_mai_n776_));
  NO4        m0748(.A(mai_mai_n476_), .B(mai_mai_n428_), .C(j), .D(f), .Y(mai_mai_n777_));
  OAI220     m0749(.A0(mai_mai_n701_), .A1(mai_mai_n693_), .B0(mai_mai_n328_), .B1(mai_mai_n38_), .Y(mai_mai_n778_));
  AOI210     m0750(.A0(mai_mai_n777_), .A1(mai_mai_n261_), .B0(mai_mai_n778_), .Y(mai_mai_n779_));
  NA3        m0751(.A(mai_mai_n540_), .B(mai_mai_n289_), .C(h), .Y(mai_mai_n780_));
  NOi21      m0752(.An(mai_mai_n670_), .B(mai_mai_n780_), .Y(mai_mai_n781_));
  NO2        m0753(.A(mai_mai_n94_), .B(mai_mai_n47_), .Y(mai_mai_n782_));
  OAI220     m0754(.A0(mai_mai_n780_), .A1(mai_mai_n601_), .B0(mai_mai_n749_), .B1(mai_mai_n663_), .Y(mai_mai_n783_));
  AOI210     m0755(.A0(mai_mai_n782_), .A1(mai_mai_n640_), .B0(mai_mai_n783_), .Y(mai_mai_n784_));
  NAi41      m0756(.An(mai_mai_n781_), .B(mai_mai_n784_), .C(mai_mai_n779_), .D(mai_mai_n776_), .Y(mai_mai_n785_));
  OR2        m0757(.A(mai_mai_n769_), .B(mai_mai_n98_), .Y(mai_mai_n786_));
  AOI220     m0758(.A0(mai_mai_n786_), .A1(mai_mai_n240_), .B0(mai_mai_n755_), .B1(mai_mai_n632_), .Y(mai_mai_n787_));
  NO2        m0759(.A(mai_mai_n658_), .B(mai_mai_n75_), .Y(mai_mai_n788_));
  NA2        m0760(.A(mai_mai_n777_), .B(mai_mai_n788_), .Y(mai_mai_n789_));
  OAI210     m0761(.A0(mai_mai_n725_), .A1(mai_mai_n656_), .B0(mai_mai_n511_), .Y(mai_mai_n790_));
  NA3        m0762(.A(mai_mai_n252_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n791_));
  AOI220     m0763(.A0(mai_mai_n600_), .A1(mai_mai_n29_), .B0(mai_mai_n457_), .B1(mai_mai_n86_), .Y(mai_mai_n792_));
  NA2        m0764(.A(mai_mai_n792_), .B(mai_mai_n791_), .Y(mai_mai_n793_));
  NO2        m0765(.A(mai_mai_n780_), .B(mai_mai_n481_), .Y(mai_mai_n794_));
  AOI210     m0766(.A0(mai_mai_n793_), .A1(mai_mai_n790_), .B0(mai_mai_n794_), .Y(mai_mai_n795_));
  NA3        m0767(.A(mai_mai_n795_), .B(mai_mai_n789_), .C(mai_mai_n787_), .Y(mai_mai_n796_));
  NOi41      m0768(.An(mai_mai_n752_), .B(mai_mai_n796_), .C(mai_mai_n785_), .D(mai_mai_n774_), .Y(mai_mai_n797_));
  OR3        m0769(.A(mai_mai_n701_), .B(mai_mai_n234_), .C(g), .Y(mai_mai_n798_));
  NO3        m0770(.A(mai_mai_n337_), .B(mai_mai_n297_), .C(mai_mai_n114_), .Y(mai_mai_n799_));
  NA2        m0771(.A(mai_mai_n799_), .B(mai_mai_n761_), .Y(mai_mai_n800_));
  INV        m0772(.A(mai_mai_n46_), .Y(mai_mai_n801_));
  NO3        m0773(.A(mai_mai_n801_), .B(mai_mai_n750_), .C(mai_mai_n277_), .Y(mai_mai_n802_));
  NO3        m0774(.A(mai_mai_n518_), .B(mai_mai_n96_), .C(h), .Y(mai_mai_n803_));
  AOI210     m0775(.A0(mai_mai_n803_), .A1(mai_mai_n696_), .B0(mai_mai_n802_), .Y(mai_mai_n804_));
  NA4        m0776(.A(mai_mai_n804_), .B(mai_mai_n800_), .C(mai_mai_n798_), .D(mai_mai_n397_), .Y(mai_mai_n805_));
  OR2        m0777(.A(mai_mai_n656_), .B(mai_mai_n94_), .Y(mai_mai_n806_));
  NO2        m0778(.A(mai_mai_n1464_), .B(n), .Y(mai_mai_n807_));
  NOi21      m0779(.An(mai_mai_n792_), .B(mai_mai_n807_), .Y(mai_mai_n808_));
  OAI220     m0780(.A0(mai_mai_n808_), .A1(mai_mai_n806_), .B0(mai_mai_n780_), .B1(mai_mai_n599_), .Y(mai_mai_n809_));
  NO2        m0781(.A(mai_mai_n323_), .B(mai_mai_n119_), .Y(mai_mai_n810_));
  NOi21      m0782(.An(mai_mai_n810_), .B(mai_mai_n164_), .Y(mai_mai_n811_));
  AOI210     m0783(.A0(mai_mai_n799_), .A1(c), .B0(mai_mai_n811_), .Y(mai_mai_n812_));
  OAI210     m0784(.A0(mai_mai_n701_), .A1(mai_mai_n387_), .B0(mai_mai_n812_), .Y(mai_mai_n813_));
  NA2        m0785(.A(mai_mai_n196_), .B(mai_mai_n692_), .Y(mai_mai_n814_));
  NO2        m0786(.A(mai_mai_n319_), .B(mai_mai_n239_), .Y(mai_mai_n815_));
  OAI210     m0787(.A0(mai_mai_n98_), .A1(mai_mai_n95_), .B0(mai_mai_n815_), .Y(mai_mai_n816_));
  NA2        m0788(.A(mai_mai_n122_), .B(mai_mai_n86_), .Y(mai_mai_n817_));
  AOI210     m0789(.A0(mai_mai_n418_), .A1(mai_mai_n410_), .B0(mai_mai_n817_), .Y(mai_mai_n818_));
  NAi21      m0790(.An(mai_mai_n818_), .B(mai_mai_n816_), .Y(mai_mai_n819_));
  NA2        m0791(.A(mai_mai_n723_), .B(mai_mai_n34_), .Y(mai_mai_n820_));
  NAi21      m0792(.An(mai_mai_n729_), .B(mai_mai_n429_), .Y(mai_mai_n821_));
  NO2        m0793(.A(mai_mai_n272_), .B(i), .Y(mai_mai_n822_));
  NA2        m0794(.A(mai_mai_n708_), .B(mai_mai_n343_), .Y(mai_mai_n823_));
  OAI210     m0795(.A0(mai_mai_n591_), .A1(mai_mai_n590_), .B0(mai_mai_n358_), .Y(mai_mai_n824_));
  AN3        m0796(.A(mai_mai_n824_), .B(mai_mai_n823_), .C(mai_mai_n821_), .Y(mai_mai_n825_));
  NAi41      m0797(.An(mai_mai_n819_), .B(mai_mai_n825_), .C(mai_mai_n820_), .D(mai_mai_n814_), .Y(mai_mai_n826_));
  NO4        m0798(.A(mai_mai_n826_), .B(mai_mai_n813_), .C(mai_mai_n809_), .D(mai_mai_n805_), .Y(mai_mai_n827_));
  NA4        m0799(.A(mai_mai_n827_), .B(mai_mai_n797_), .C(mai_mai_n747_), .D(mai_mai_n734_), .Y(mai09));
  INV        m0800(.A(mai_mai_n123_), .Y(mai_mai_n829_));
  NA2        m0801(.A(f), .B(e), .Y(mai_mai_n830_));
  NA2        m0802(.A(l), .B(g), .Y(mai_mai_n831_));
  NO2        m0803(.A(g), .B(mai_mai_n462_), .Y(mai_mai_n832_));
  AOI210     m0804(.A0(mai_mai_n832_), .A1(mai_mai_n831_), .B0(mai_mai_n830_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n833_), .B(mai_mai_n829_), .Y(mai_mai_n834_));
  NO2        m0806(.A(mai_mai_n208_), .B(mai_mai_n218_), .Y(mai_mai_n835_));
  NA3        m0807(.A(m), .B(l), .C(i), .Y(mai_mai_n836_));
  OAI220     m0808(.A0(mai_mai_n585_), .A1(mai_mai_n836_), .B0(mai_mai_n348_), .B1(mai_mai_n519_), .Y(mai_mai_n837_));
  NA4        m0809(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(g), .D(f), .Y(mai_mai_n838_));
  NAi31      m0810(.An(mai_mai_n837_), .B(mai_mai_n838_), .C(mai_mai_n433_), .Y(mai_mai_n839_));
  OA210      m0811(.A0(mai_mai_n839_), .A1(mai_mai_n835_), .B0(mai_mai_n561_), .Y(mai_mai_n840_));
  NA3        m0812(.A(mai_mai_n806_), .B(mai_mai_n563_), .C(mai_mai_n511_), .Y(mai_mai_n841_));
  OA210      m0813(.A0(mai_mai_n841_), .A1(mai_mai_n840_), .B0(mai_mai_n807_), .Y(mai_mai_n842_));
  INV        m0814(.A(mai_mai_n334_), .Y(mai_mai_n843_));
  NO2        m0815(.A(mai_mai_n129_), .B(mai_mai_n127_), .Y(mai_mai_n844_));
  NOi31      m0816(.An(k), .B(m), .C(l), .Y(mai_mai_n845_));
  NO2        m0817(.A(mai_mai_n336_), .B(mai_mai_n845_), .Y(mai_mai_n846_));
  AOI210     m0818(.A0(mai_mai_n846_), .A1(mai_mai_n844_), .B0(mai_mai_n594_), .Y(mai_mai_n847_));
  NA2        m0819(.A(mai_mai_n791_), .B(mai_mai_n328_), .Y(mai_mai_n848_));
  NA2        m0820(.A(mai_mai_n338_), .B(m), .Y(mai_mai_n849_));
  OAI210     m0821(.A0(mai_mai_n208_), .A1(mai_mai_n218_), .B0(mai_mai_n849_), .Y(mai_mai_n850_));
  AOI220     m0822(.A0(mai_mai_n850_), .A1(mai_mai_n848_), .B0(mai_mai_n847_), .B1(mai_mai_n843_), .Y(mai_mai_n851_));
  NA2        m0823(.A(mai_mai_n171_), .B(mai_mai_n116_), .Y(mai_mai_n852_));
  NA3        m0824(.A(mai_mai_n852_), .B(mai_mai_n691_), .C(mai_mai_n138_), .Y(mai_mai_n853_));
  NA3        m0825(.A(mai_mai_n853_), .B(mai_mai_n194_), .C(mai_mai_n31_), .Y(mai_mai_n854_));
  NA4        m0826(.A(mai_mai_n854_), .B(mai_mai_n851_), .C(mai_mai_n620_), .D(mai_mai_n84_), .Y(mai_mai_n855_));
  NO2        m0827(.A(mai_mai_n581_), .B(mai_mai_n490_), .Y(mai_mai_n856_));
  NA2        m0828(.A(mai_mai_n856_), .B(mai_mai_n194_), .Y(mai_mai_n857_));
  NOi21      m0829(.An(f), .B(d), .Y(mai_mai_n858_));
  NA2        m0830(.A(mai_mai_n858_), .B(m), .Y(mai_mai_n859_));
  NO2        m0831(.A(mai_mai_n859_), .B(mai_mai_n52_), .Y(mai_mai_n860_));
  NOi32      m0832(.An(g), .Bn(f), .C(d), .Y(mai_mai_n861_));
  NA4        m0833(.A(mai_mai_n861_), .B(mai_mai_n600_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n862_));
  INV        m0834(.A(mai_mai_n862_), .Y(mai_mai_n863_));
  AOI210     m0835(.A0(mai_mai_n860_), .A1(mai_mai_n538_), .B0(mai_mai_n863_), .Y(mai_mai_n864_));
  AN2        m0836(.A(f), .B(d), .Y(mai_mai_n865_));
  NA3        m0837(.A(mai_mai_n467_), .B(mai_mai_n865_), .C(mai_mai_n86_), .Y(mai_mai_n866_));
  NO3        m0838(.A(mai_mai_n866_), .B(mai_mai_n75_), .C(mai_mai_n219_), .Y(mai_mai_n867_));
  INV        m0839(.A(mai_mai_n867_), .Y(mai_mai_n868_));
  NAi41      m0840(.An(mai_mai_n480_), .B(mai_mai_n868_), .C(mai_mai_n864_), .D(mai_mai_n857_), .Y(mai_mai_n869_));
  NO3        m0841(.A(mai_mai_n134_), .B(mai_mai_n323_), .C(mai_mai_n155_), .Y(mai_mai_n870_));
  NO2        m0842(.A(mai_mai_n649_), .B(mai_mai_n323_), .Y(mai_mai_n871_));
  AN2        m0843(.A(mai_mai_n871_), .B(mai_mai_n674_), .Y(mai_mai_n872_));
  NO3        m0844(.A(mai_mai_n872_), .B(mai_mai_n870_), .C(mai_mai_n236_), .Y(mai_mai_n873_));
  NA2        m0845(.A(mai_mai_n598_), .B(mai_mai_n86_), .Y(mai_mai_n874_));
  OAI220     m0846(.A0(mai_mai_n849_), .A1(mai_mai_n874_), .B0(mai_mai_n791_), .B1(mai_mai_n433_), .Y(mai_mai_n875_));
  NA3        m0847(.A(mai_mai_n163_), .B(mai_mai_n110_), .C(g), .Y(mai_mai_n876_));
  OAI220     m0848(.A0(mai_mai_n866_), .A1(mai_mai_n423_), .B0(mai_mai_n334_), .B1(mai_mai_n876_), .Y(mai_mai_n877_));
  NOi41      m0849(.An(mai_mai_n229_), .B(mai_mai_n877_), .C(mai_mai_n875_), .D(mai_mai_n304_), .Y(mai_mai_n878_));
  NA2        m0850(.A(c), .B(mai_mai_n118_), .Y(mai_mai_n879_));
  NO2        m0851(.A(mai_mai_n879_), .B(mai_mai_n401_), .Y(mai_mai_n880_));
  NA3        m0852(.A(mai_mai_n880_), .B(mai_mai_n502_), .C(f), .Y(mai_mai_n881_));
  OR2        m0853(.A(mai_mai_n656_), .B(mai_mai_n534_), .Y(mai_mai_n882_));
  INV        m0854(.A(mai_mai_n882_), .Y(mai_mai_n883_));
  NA2        m0855(.A(b), .B(mai_mai_n883_), .Y(mai_mai_n884_));
  NA4        m0856(.A(mai_mai_n884_), .B(mai_mai_n881_), .C(mai_mai_n878_), .D(mai_mai_n873_), .Y(mai_mai_n885_));
  NO4        m0857(.A(mai_mai_n885_), .B(mai_mai_n869_), .C(mai_mai_n855_), .D(mai_mai_n842_), .Y(mai_mai_n886_));
  OR2        m0858(.A(mai_mai_n866_), .B(mai_mai_n75_), .Y(mai_mai_n887_));
  INV        m0859(.A(g), .Y(mai_mai_n888_));
  AOI210     m0860(.A0(mai_mai_n888_), .A1(mai_mai_n290_), .B0(mai_mai_n887_), .Y(mai_mai_n889_));
  AOI210     m0861(.A0(mai_mai_n791_), .A1(mai_mai_n328_), .B0(mai_mai_n838_), .Y(mai_mai_n890_));
  NO2        m0862(.A(mai_mai_n138_), .B(mai_mai_n134_), .Y(mai_mai_n891_));
  NA2        m0863(.A(mai_mai_n302_), .B(mai_mai_n891_), .Y(mai_mai_n892_));
  NO2        m0864(.A(mai_mai_n423_), .B(mai_mai_n830_), .Y(mai_mai_n893_));
  NA2        m0865(.A(mai_mai_n893_), .B(mai_mai_n555_), .Y(mai_mai_n894_));
  NA2        m0866(.A(mai_mai_n894_), .B(mai_mai_n892_), .Y(mai_mai_n895_));
  NA2        m0867(.A(e), .B(d), .Y(mai_mai_n896_));
  OAI220     m0868(.A0(mai_mai_n896_), .A1(c), .B0(mai_mai_n319_), .B1(d), .Y(mai_mai_n897_));
  NA3        m0869(.A(mai_mai_n897_), .B(mai_mai_n448_), .C(mai_mai_n500_), .Y(mai_mai_n898_));
  NO2        m0870(.A(mai_mai_n184_), .B(mai_mai_n232_), .Y(mai_mai_n899_));
  AOI210     m0871(.A0(mai_mai_n619_), .A1(mai_mai_n341_), .B0(mai_mai_n899_), .Y(mai_mai_n900_));
  NA2        m0872(.A(mai_mai_n867_), .B(j), .Y(mai_mai_n901_));
  NA3        m0873(.A(mai_mai_n170_), .B(mai_mai_n87_), .C(mai_mai_n34_), .Y(mai_mai_n902_));
  NA4        m0874(.A(mai_mai_n902_), .B(mai_mai_n901_), .C(mai_mai_n900_), .D(mai_mai_n898_), .Y(mai_mai_n903_));
  NO4        m0875(.A(mai_mai_n903_), .B(mai_mai_n895_), .C(mai_mai_n890_), .D(mai_mai_n889_), .Y(mai_mai_n904_));
  NA2        m0876(.A(mai_mai_n843_), .B(mai_mai_n31_), .Y(mai_mai_n905_));
  AO210      m0877(.A0(mai_mai_n905_), .A1(mai_mai_n693_), .B0(mai_mai_n222_), .Y(mai_mai_n906_));
  OAI210     m0878(.A0(mai_mai_n297_), .A1(j), .B0(mai_mai_n61_), .Y(mai_mai_n907_));
  AOI220     m0879(.A0(mai_mai_n907_), .A1(mai_mai_n871_), .B0(mai_mai_n610_), .B1(mai_mai_n618_), .Y(mai_mai_n908_));
  INV        m0880(.A(mai_mai_n908_), .Y(mai_mai_n909_));
  OAI210     m0881(.A0(l), .A1(j), .B0(mai_mai_n861_), .Y(mai_mai_n910_));
  NO2        m0882(.A(mai_mai_n910_), .B(mai_mai_n601_), .Y(mai_mai_n911_));
  INV        m0883(.A(mai_mai_n862_), .Y(mai_mai_n912_));
  AO210      m0884(.A0(mai_mai_n848_), .A1(mai_mai_n837_), .B0(mai_mai_n912_), .Y(mai_mai_n913_));
  NOi31      m0885(.An(mai_mai_n538_), .B(mai_mai_n859_), .C(mai_mai_n290_), .Y(mai_mai_n914_));
  NO4        m0886(.A(mai_mai_n914_), .B(mai_mai_n913_), .C(mai_mai_n911_), .D(mai_mai_n909_), .Y(mai_mai_n915_));
  AO220      m0887(.A0(mai_mai_n448_), .A1(mai_mai_n742_), .B0(mai_mai_n179_), .B1(f), .Y(mai_mai_n916_));
  NA2        m0888(.A(mai_mai_n916_), .B(mai_mai_n897_), .Y(mai_mai_n917_));
  NO2        m0889(.A(mai_mai_n432_), .B(mai_mai_n71_), .Y(mai_mai_n918_));
  OAI210     m0890(.A0(mai_mai_n841_), .A1(mai_mai_n918_), .B0(mai_mai_n696_), .Y(mai_mai_n919_));
  AN4        m0891(.A(mai_mai_n919_), .B(mai_mai_n917_), .C(mai_mai_n915_), .D(mai_mai_n906_), .Y(mai_mai_n920_));
  NA4        m0892(.A(mai_mai_n920_), .B(mai_mai_n904_), .C(mai_mai_n886_), .D(mai_mai_n834_), .Y(mai12));
  NO2        m0893(.A(mai_mai_n447_), .B(c), .Y(mai_mai_n922_));
  NO4        m0894(.A(mai_mai_n437_), .B(mai_mai_n255_), .C(mai_mai_n579_), .D(mai_mai_n219_), .Y(mai_mai_n923_));
  NA2        m0895(.A(mai_mai_n923_), .B(mai_mai_n922_), .Y(mai_mai_n924_));
  NA2        m0896(.A(mai_mai_n538_), .B(mai_mai_n918_), .Y(mai_mai_n925_));
  NO3        m0897(.A(mai_mai_n447_), .B(mai_mai_n86_), .C(mai_mai_n118_), .Y(mai_mai_n926_));
  NO2        m0898(.A(mai_mai_n844_), .B(mai_mai_n348_), .Y(mai_mai_n927_));
  NO2        m0899(.A(mai_mai_n656_), .B(mai_mai_n374_), .Y(mai_mai_n928_));
  AOI220     m0900(.A0(mai_mai_n928_), .A1(mai_mai_n536_), .B0(mai_mai_n927_), .B1(mai_mai_n926_), .Y(mai_mai_n929_));
  NA4        m0901(.A(mai_mai_n929_), .B(mai_mai_n925_), .C(mai_mai_n924_), .D(mai_mai_n436_), .Y(mai_mai_n930_));
  AOI210     m0902(.A0(mai_mai_n235_), .A1(mai_mai_n333_), .B0(mai_mai_n205_), .Y(mai_mai_n931_));
  NO2        m0903(.A(mai_mai_n637_), .B(mai_mai_n263_), .Y(mai_mai_n932_));
  NO2        m0904(.A(mai_mai_n585_), .B(mai_mai_n836_), .Y(mai_mai_n933_));
  AOI220     m0905(.A0(mai_mai_n933_), .A1(mai_mai_n561_), .B0(mai_mai_n815_), .B1(mai_mai_n932_), .Y(mai_mai_n934_));
  NO2        m0906(.A(mai_mai_n154_), .B(mai_mai_n239_), .Y(mai_mai_n935_));
  NA3        m0907(.A(mai_mai_n935_), .B(mai_mai_n242_), .C(i), .Y(mai_mai_n936_));
  NA2        m0908(.A(mai_mai_n936_), .B(mai_mai_n934_), .Y(mai_mai_n937_));
  OR2        m0909(.A(c), .B(mai_mai_n926_), .Y(mai_mai_n938_));
  NA2        m0910(.A(mai_mai_n938_), .B(mai_mai_n349_), .Y(mai_mai_n939_));
  NO3        m0911(.A(mai_mai_n134_), .B(mai_mai_n155_), .C(mai_mai_n219_), .Y(mai_mai_n940_));
  NA2        m0912(.A(mai_mai_n940_), .B(mai_mai_n523_), .Y(mai_mai_n941_));
  NA4        m0913(.A(mai_mai_n438_), .B(d), .C(mai_mai_n185_), .D(g), .Y(mai_mai_n942_));
  NA3        m0914(.A(mai_mai_n942_), .B(mai_mai_n941_), .C(mai_mai_n939_), .Y(mai_mai_n943_));
  NO3        m0915(.A(mai_mai_n661_), .B(mai_mai_n94_), .C(mai_mai_n45_), .Y(mai_mai_n944_));
  NO4        m0916(.A(mai_mai_n944_), .B(mai_mai_n943_), .C(mai_mai_n937_), .D(mai_mai_n930_), .Y(mai_mai_n945_));
  NO2        m0917(.A(mai_mai_n1462_), .B(mai_mai_n364_), .Y(mai_mai_n946_));
  NA2        m0918(.A(mai_mai_n582_), .B(mai_mai_n73_), .Y(mai_mai_n947_));
  NOi21      m0919(.An(mai_mai_n34_), .B(mai_mai_n649_), .Y(mai_mai_n948_));
  AOI220     m0920(.A0(mai_mai_n948_), .A1(c), .B0(mai_mai_n947_), .B1(mai_mai_n946_), .Y(mai_mai_n949_));
  OAI210     m0921(.A0(mai_mai_n253_), .A1(mai_mai_n45_), .B0(mai_mai_n949_), .Y(mai_mai_n950_));
  NA2        m0922(.A(mai_mai_n429_), .B(mai_mai_n265_), .Y(mai_mai_n951_));
  NO3        m0923(.A(mai_mai_n817_), .B(mai_mai_n91_), .C(mai_mai_n401_), .Y(mai_mai_n952_));
  NAi31      m0924(.An(mai_mai_n952_), .B(mai_mai_n951_), .C(mai_mai_n317_), .Y(mai_mai_n953_));
  NO2        m0925(.A(mai_mai_n497_), .B(mai_mai_n297_), .Y(mai_mai_n954_));
  NO2        m0926(.A(mai_mai_n954_), .B(mai_mai_n361_), .Y(mai_mai_n955_));
  NO2        m0927(.A(mai_mai_n955_), .B(mai_mai_n147_), .Y(mai_mai_n956_));
  INV        m0928(.A(mai_mai_n628_), .Y(mai_mai_n957_));
  OAI210     m0929(.A0(mai_mai_n730_), .A1(mai_mai_n957_), .B0(mai_mai_n362_), .Y(mai_mai_n958_));
  NO4        m0930(.A(mai_mai_n958_), .B(mai_mai_n956_), .C(mai_mai_n953_), .D(mai_mai_n950_), .Y(mai_mai_n959_));
  NA2        m0931(.A(mai_mai_n341_), .B(g), .Y(mai_mai_n960_));
  NA2        m0932(.A(h), .B(i), .Y(mai_mai_n961_));
  NA2        m0933(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n962_));
  OAI220     m0934(.A0(mai_mai_n962_), .A1(mai_mai_n1460_), .B0(mai_mai_n961_), .B1(mai_mai_n94_), .Y(mai_mai_n963_));
  AOI210     m0935(.A0(mai_mai_n412_), .A1(mai_mai_n37_), .B0(mai_mai_n963_), .Y(mai_mai_n964_));
  NO2        m0936(.A(mai_mai_n147_), .B(mai_mai_n86_), .Y(mai_mai_n965_));
  OR2        m0937(.A(mai_mai_n965_), .B(mai_mai_n547_), .Y(mai_mai_n966_));
  AOI210     m0938(.A0(c), .A1(n), .B0(mai_mai_n966_), .Y(mai_mai_n967_));
  OAI220     m0939(.A0(mai_mai_n967_), .A1(mai_mai_n960_), .B0(mai_mai_n964_), .B1(mai_mai_n328_), .Y(mai_mai_n968_));
  NO2        m0940(.A(mai_mai_n656_), .B(mai_mai_n490_), .Y(mai_mai_n969_));
  NA3        m0941(.A(mai_mai_n338_), .B(j), .C(i), .Y(mai_mai_n970_));
  OAI220     m0942(.A0(mai_mai_n1458_), .A1(mai_mai_n969_), .B0(mai_mai_n670_), .B1(mai_mai_n754_), .Y(mai_mai_n971_));
  NA2        m0943(.A(mai_mai_n604_), .B(mai_mai_n115_), .Y(mai_mai_n972_));
  NA3        m0944(.A(j), .B(mai_mai_n82_), .C(i), .Y(mai_mai_n973_));
  OA220      m0945(.A0(mai_mai_n973_), .A1(mai_mai_n972_), .B0(mai_mai_n428_), .B1(mai_mai_n584_), .Y(mai_mai_n974_));
  NA3        m0946(.A(mai_mai_n320_), .B(mai_mai_n120_), .C(g), .Y(mai_mai_n975_));
  AOI210     m0947(.A0(mai_mai_n667_), .A1(mai_mai_n975_), .B0(m), .Y(mai_mai_n976_));
  OAI210     m0948(.A0(mai_mai_n976_), .A1(mai_mai_n927_), .B0(c), .Y(mai_mai_n977_));
  NA2        m0949(.A(mai_mai_n684_), .B(mai_mai_n874_), .Y(mai_mai_n978_));
  NA2        m0950(.A(mai_mai_n838_), .B(mai_mai_n433_), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n227_), .B(mai_mai_n79_), .Y(mai_mai_n980_));
  NA3        m0952(.A(mai_mai_n980_), .B(mai_mai_n973_), .C(mai_mai_n428_), .Y(mai_mai_n981_));
  AOI220     m0953(.A0(mai_mai_n981_), .A1(mai_mai_n261_), .B0(mai_mai_n979_), .B1(mai_mai_n978_), .Y(mai_mai_n982_));
  NA4        m0954(.A(mai_mai_n982_), .B(mai_mai_n977_), .C(mai_mai_n974_), .D(mai_mai_n971_), .Y(mai_mai_n983_));
  NO2        m0955(.A(mai_mai_n374_), .B(mai_mai_n93_), .Y(mai_mai_n984_));
  OAI210     m0956(.A0(mai_mai_n984_), .A1(mai_mai_n932_), .B0(mai_mai_n240_), .Y(mai_mai_n985_));
  NA2        m0957(.A(mai_mai_n660_), .B(mai_mai_n90_), .Y(mai_mai_n986_));
  NO2        m0958(.A(mai_mai_n453_), .B(mai_mai_n219_), .Y(mai_mai_n987_));
  AOI220     m0959(.A0(mai_mai_n987_), .A1(mai_mai_n379_), .B0(mai_mai_n938_), .B1(mai_mai_n223_), .Y(mai_mai_n988_));
  AOI220     m0960(.A0(mai_mai_n928_), .A1(mai_mai_n935_), .B0(mai_mai_n583_), .B1(mai_mai_n92_), .Y(mai_mai_n989_));
  NA4        m0961(.A(mai_mai_n989_), .B(mai_mai_n988_), .C(mai_mai_n986_), .D(mai_mai_n985_), .Y(mai_mai_n990_));
  OAI210     m0962(.A0(mai_mai_n979_), .A1(mai_mai_n933_), .B0(mai_mai_n536_), .Y(mai_mai_n991_));
  AOI210     m0963(.A0(mai_mai_n413_), .A1(mai_mai_n405_), .B0(mai_mai_n817_), .Y(mai_mai_n992_));
  OAI210     m0964(.A0(mai_mai_n1462_), .A1(mai_mai_n364_), .B0(mai_mai_n111_), .Y(mai_mai_n993_));
  AOI210     m0965(.A0(mai_mai_n993_), .A1(mai_mai_n528_), .B0(mai_mai_n992_), .Y(mai_mai_n994_));
  NA2        m0966(.A(mai_mai_n976_), .B(mai_mai_n926_), .Y(mai_mai_n995_));
  NO2        m0967(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n996_));
  AOI220     m0968(.A0(mai_mai_n996_), .A1(mai_mai_n622_), .B0(mai_mai_n642_), .B1(mai_mai_n523_), .Y(mai_mai_n997_));
  NA4        m0969(.A(mai_mai_n997_), .B(mai_mai_n995_), .C(mai_mai_n994_), .D(mai_mai_n991_), .Y(mai_mai_n998_));
  NO4        m0970(.A(mai_mai_n998_), .B(mai_mai_n990_), .C(mai_mai_n983_), .D(mai_mai_n968_), .Y(mai_mai_n999_));
  NAi31      m0971(.An(mai_mai_n144_), .B(mai_mai_n414_), .C(n), .Y(mai_mai_n1000_));
  NO3        m0972(.A(mai_mai_n127_), .B(mai_mai_n336_), .C(mai_mai_n845_), .Y(mai_mai_n1001_));
  NO2        m0973(.A(mai_mai_n1001_), .B(mai_mai_n1000_), .Y(mai_mai_n1002_));
  NO3        m0974(.A(mai_mai_n272_), .B(mai_mai_n144_), .C(mai_mai_n401_), .Y(mai_mai_n1003_));
  AOI210     m0975(.A0(mai_mai_n1003_), .A1(mai_mai_n491_), .B0(mai_mai_n1002_), .Y(mai_mai_n1004_));
  NA2        m0976(.A(mai_mai_n483_), .B(i), .Y(mai_mai_n1005_));
  NA2        m0977(.A(mai_mai_n1005_), .B(mai_mai_n1004_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n232_), .B(mai_mai_n175_), .Y(mai_mai_n1007_));
  NO3        m0979(.A(mai_mai_n306_), .B(mai_mai_n438_), .C(mai_mai_n179_), .Y(mai_mai_n1008_));
  NOi31      m0980(.An(mai_mai_n1007_), .B(mai_mai_n1008_), .C(mai_mai_n219_), .Y(mai_mai_n1009_));
  NO3        m0981(.A(mai_mai_n432_), .B(k), .C(mai_mai_n75_), .Y(mai_mai_n1010_));
  NA2        m0982(.A(mai_mai_n1010_), .B(mai_mai_n430_), .Y(mai_mai_n1011_));
  INV        m0983(.A(mai_mai_n1011_), .Y(mai_mai_n1012_));
  OAI220     m0984(.A0(mai_mai_n1000_), .A1(mai_mai_n235_), .B0(mai_mai_n970_), .B1(mai_mai_n599_), .Y(mai_mai_n1013_));
  NO2        m0985(.A(mai_mai_n657_), .B(mai_mai_n374_), .Y(mai_mai_n1014_));
  NA2        m0986(.A(mai_mai_n931_), .B(mai_mai_n922_), .Y(mai_mai_n1015_));
  NO3        m0987(.A(mai_mai_n537_), .B(mai_mai_n152_), .C(mai_mai_n218_), .Y(mai_mai_n1016_));
  OAI210     m0988(.A0(mai_mai_n1016_), .A1(mai_mai_n517_), .B0(mai_mai_n375_), .Y(mai_mai_n1017_));
  OAI220     m0989(.A0(mai_mai_n928_), .A1(mai_mai_n933_), .B0(mai_mai_n538_), .B1(mai_mai_n422_), .Y(mai_mai_n1018_));
  NA4        m0990(.A(mai_mai_n1018_), .B(mai_mai_n1017_), .C(mai_mai_n1015_), .D(mai_mai_n617_), .Y(mai_mai_n1019_));
  OAI210     m0991(.A0(mai_mai_n931_), .A1(mai_mai_n923_), .B0(mai_mai_n1007_), .Y(mai_mai_n1020_));
  NA3        m0992(.A(c), .B(mai_mai_n478_), .C(mai_mai_n46_), .Y(mai_mai_n1021_));
  AOI210     m0993(.A0(mai_mai_n377_), .A1(mai_mai_n375_), .B0(mai_mai_n327_), .Y(mai_mai_n1022_));
  NA4        m0994(.A(mai_mai_n1022_), .B(mai_mai_n1021_), .C(mai_mai_n1020_), .D(mai_mai_n273_), .Y(mai_mai_n1023_));
  OR4        m0995(.A(mai_mai_n1023_), .B(mai_mai_n1019_), .C(mai_mai_n1014_), .D(mai_mai_n1013_), .Y(mai_mai_n1024_));
  NO4        m0996(.A(mai_mai_n1024_), .B(mai_mai_n1012_), .C(mai_mai_n1009_), .D(mai_mai_n1006_), .Y(mai_mai_n1025_));
  NA4        m0997(.A(mai_mai_n1025_), .B(mai_mai_n999_), .C(mai_mai_n959_), .D(mai_mai_n945_), .Y(mai13));
  AN2        m0998(.A(c), .B(b), .Y(mai_mai_n1027_));
  NA3        m0999(.A(mai_mai_n252_), .B(mai_mai_n1027_), .C(m), .Y(mai_mai_n1028_));
  NA2        m1000(.A(mai_mai_n488_), .B(f), .Y(mai_mai_n1029_));
  NO4        m1001(.A(mai_mai_n1029_), .B(mai_mai_n1028_), .C(j), .D(k), .Y(mai_mai_n1030_));
  INV        m1002(.A(mai_mai_n265_), .Y(mai_mai_n1031_));
  NO4        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1029_), .C(mai_mai_n961_), .D(a), .Y(mai_mai_n1032_));
  NAi32      m1004(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1033_));
  NA2        m1005(.A(mai_mai_n143_), .B(mai_mai_n45_), .Y(mai_mai_n1034_));
  NO4        m1006(.A(mai_mai_n1034_), .B(mai_mai_n1033_), .C(mai_mai_n585_), .D(mai_mai_n305_), .Y(mai_mai_n1035_));
  NA2        m1007(.A(mai_mai_n404_), .B(mai_mai_n218_), .Y(mai_mai_n1036_));
  AN2        m1008(.A(d), .B(c), .Y(mai_mai_n1037_));
  NA2        m1009(.A(mai_mai_n1037_), .B(mai_mai_n118_), .Y(mai_mai_n1038_));
  NO4        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1036_), .C(mai_mai_n180_), .D(mai_mai_n171_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n488_), .B(c), .Y(mai_mai_n1040_));
  NO4        m1012(.A(mai_mai_n1034_), .B(mai_mai_n581_), .C(mai_mai_n1040_), .D(mai_mai_n305_), .Y(mai_mai_n1041_));
  OR2        m1013(.A(mai_mai_n1039_), .B(mai_mai_n1041_), .Y(mai_mai_n1042_));
  OR4        m1014(.A(mai_mai_n1042_), .B(mai_mai_n1035_), .C(mai_mai_n1032_), .D(mai_mai_n1030_), .Y(mai_mai_n1043_));
  NAi32      m1015(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1044_));
  NO2        m1016(.A(mai_mai_n1044_), .B(mai_mai_n149_), .Y(mai_mai_n1045_));
  NA2        m1017(.A(mai_mai_n1045_), .B(g), .Y(mai_mai_n1046_));
  OR3        m1018(.A(mai_mai_n230_), .B(mai_mai_n180_), .C(mai_mai_n171_), .Y(mai_mai_n1047_));
  NO2        m1019(.A(mai_mai_n1047_), .B(mai_mai_n1046_), .Y(mai_mai_n1048_));
  NO2        m1020(.A(mai_mai_n1040_), .B(mai_mai_n305_), .Y(mai_mai_n1049_));
  NA2        m1021(.A(mai_mai_n625_), .B(mai_mai_n1461_), .Y(mai_mai_n1050_));
  NOi21      m1022(.An(mai_mai_n1049_), .B(mai_mai_n1050_), .Y(mai_mai_n1051_));
  NOi41      m1023(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1052_));
  NA2        m1024(.A(mai_mai_n1052_), .B(j), .Y(mai_mai_n1053_));
  NO2        m1025(.A(mai_mai_n1053_), .B(mai_mai_n1046_), .Y(mai_mai_n1054_));
  OR3        m1026(.A(e), .B(d), .C(c), .Y(mai_mai_n1055_));
  NA3        m1027(.A(k), .B(j), .C(i), .Y(mai_mai_n1056_));
  NO3        m1028(.A(mai_mai_n1056_), .B(mai_mai_n305_), .C(mai_mai_n93_), .Y(mai_mai_n1057_));
  NOi21      m1029(.An(mai_mai_n1057_), .B(mai_mai_n1055_), .Y(mai_mai_n1058_));
  OR4        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1054_), .C(mai_mai_n1051_), .D(mai_mai_n1048_), .Y(mai_mai_n1059_));
  NA3        m1031(.A(mai_mai_n460_), .B(mai_mai_n330_), .C(mai_mai_n56_), .Y(mai_mai_n1060_));
  NO2        m1032(.A(mai_mai_n1060_), .B(mai_mai_n1050_), .Y(mai_mai_n1061_));
  NO4        m1033(.A(mai_mai_n1060_), .B(mai_mai_n581_), .C(mai_mai_n445_), .D(mai_mai_n45_), .Y(mai_mai_n1062_));
  NO2        m1034(.A(f), .B(c), .Y(mai_mai_n1063_));
  NOi21      m1035(.An(mai_mai_n1063_), .B(mai_mai_n437_), .Y(mai_mai_n1064_));
  NA2        m1036(.A(mai_mai_n1064_), .B(mai_mai_n59_), .Y(mai_mai_n1065_));
  OR2        m1037(.A(k), .B(i), .Y(mai_mai_n1066_));
  NO3        m1038(.A(mai_mai_n1066_), .B(mai_mai_n246_), .C(l), .Y(mai_mai_n1067_));
  NOi31      m1039(.An(mai_mai_n1067_), .B(mai_mai_n1065_), .C(j), .Y(mai_mai_n1068_));
  OR3        m1040(.A(mai_mai_n1068_), .B(mai_mai_n1062_), .C(mai_mai_n1061_), .Y(mai_mai_n1069_));
  OR3        m1041(.A(mai_mai_n1069_), .B(mai_mai_n1059_), .C(mai_mai_n1043_), .Y(mai02));
  OR2        m1042(.A(l), .B(k), .Y(mai_mai_n1071_));
  OR3        m1043(.A(h), .B(g), .C(f), .Y(mai_mai_n1072_));
  OR3        m1044(.A(n), .B(m), .C(i), .Y(mai_mai_n1073_));
  NO4        m1045(.A(mai_mai_n1073_), .B(mai_mai_n1072_), .C(mai_mai_n1071_), .D(mai_mai_n1055_), .Y(mai_mai_n1074_));
  NOi31      m1046(.An(e), .B(d), .C(c), .Y(mai_mai_n1075_));
  AOI210     m1047(.A0(mai_mai_n1057_), .A1(mai_mai_n1075_), .B0(mai_mai_n1035_), .Y(mai_mai_n1076_));
  AN3        m1048(.A(g), .B(f), .C(c), .Y(mai_mai_n1077_));
  NA3        m1049(.A(mai_mai_n1077_), .B(mai_mai_n460_), .C(h), .Y(mai_mai_n1078_));
  OR2        m1050(.A(mai_mai_n305_), .B(mai_mai_n1078_), .Y(mai_mai_n1079_));
  NO3        m1051(.A(mai_mai_n1060_), .B(mai_mai_n1034_), .C(mai_mai_n581_), .Y(mai_mai_n1080_));
  NO2        m1052(.A(mai_mai_n1080_), .B(mai_mai_n1048_), .Y(mai_mai_n1081_));
  NA3        m1053(.A(l), .B(k), .C(j), .Y(mai_mai_n1082_));
  NA2        m1054(.A(i), .B(h), .Y(mai_mai_n1083_));
  NO3        m1055(.A(mai_mai_n1083_), .B(mai_mai_n1082_), .C(mai_mai_n134_), .Y(mai_mai_n1084_));
  NO3        m1056(.A(mai_mai_n145_), .B(mai_mai_n282_), .C(mai_mai_n219_), .Y(mai_mai_n1085_));
  AOI210     m1057(.A0(mai_mai_n1085_), .A1(mai_mai_n1084_), .B0(mai_mai_n1051_), .Y(mai_mai_n1086_));
  NA3        m1058(.A(c), .B(b), .C(a), .Y(mai_mai_n1087_));
  NO3        m1059(.A(mai_mai_n1087_), .B(mai_mai_n896_), .C(mai_mai_n218_), .Y(mai_mai_n1088_));
  NO4        m1060(.A(mai_mai_n1056_), .B(mai_mai_n297_), .C(mai_mai_n49_), .D(mai_mai_n114_), .Y(mai_mai_n1089_));
  AOI210     m1061(.A0(mai_mai_n1089_), .A1(mai_mai_n1088_), .B0(mai_mai_n1061_), .Y(mai_mai_n1090_));
  AN4        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1086_), .C(mai_mai_n1081_), .D(mai_mai_n1079_), .Y(mai_mai_n1091_));
  NO2        m1063(.A(mai_mai_n1038_), .B(mai_mai_n1036_), .Y(mai_mai_n1092_));
  NA2        m1064(.A(mai_mai_n1053_), .B(mai_mai_n1047_), .Y(mai_mai_n1093_));
  AOI210     m1065(.A0(mai_mai_n1093_), .A1(mai_mai_n1092_), .B0(mai_mai_n1030_), .Y(mai_mai_n1094_));
  NAi41      m1066(.An(mai_mai_n1074_), .B(mai_mai_n1094_), .C(mai_mai_n1091_), .D(mai_mai_n1076_), .Y(mai03));
  NO2        m1067(.A(mai_mai_n519_), .B(mai_mai_n594_), .Y(mai_mai_n1096_));
  NA4        m1068(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(g), .D(mai_mai_n218_), .Y(mai_mai_n1097_));
  NA4        m1069(.A(mai_mai_n571_), .B(m), .C(mai_mai_n114_), .D(mai_mai_n218_), .Y(mai_mai_n1098_));
  NA3        m1070(.A(mai_mai_n1098_), .B(mai_mai_n365_), .C(mai_mai_n1097_), .Y(mai_mai_n1099_));
  NO3        m1071(.A(mai_mai_n1099_), .B(mai_mai_n1096_), .C(mai_mai_n993_), .Y(mai_mai_n1100_));
  NOi41      m1072(.An(mai_mai_n806_), .B(mai_mai_n850_), .C(mai_mai_n839_), .D(mai_mai_n710_), .Y(mai_mai_n1101_));
  OAI220     m1073(.A0(mai_mai_n1101_), .A1(mai_mai_n684_), .B0(mai_mai_n1100_), .B1(mai_mai_n582_), .Y(mai_mai_n1102_));
  NA4        m1074(.A(i), .B(mai_mai_n1075_), .C(mai_mai_n338_), .D(mai_mai_n330_), .Y(mai_mai_n1103_));
  OAI210     m1075(.A0(mai_mai_n817_), .A1(mai_mai_n415_), .B0(mai_mai_n1103_), .Y(mai_mai_n1104_));
  NOi31      m1076(.An(m), .B(n), .C(f), .Y(mai_mai_n1105_));
  NA2        m1077(.A(mai_mai_n1105_), .B(mai_mai_n51_), .Y(mai_mai_n1106_));
  AN2        m1078(.A(e), .B(c), .Y(mai_mai_n1107_));
  NA2        m1079(.A(mai_mai_n1107_), .B(a), .Y(mai_mai_n1108_));
  OAI220     m1080(.A0(mai_mai_n1108_), .A1(mai_mai_n1106_), .B0(mai_mai_n882_), .B1(mai_mai_n421_), .Y(mai_mai_n1109_));
  NOi21      m1081(.An(mai_mai_n861_), .B(mai_mai_n1028_), .Y(mai_mai_n1110_));
  NO4        m1082(.A(mai_mai_n1110_), .B(mai_mai_n1109_), .C(mai_mai_n1104_), .D(mai_mai_n992_), .Y(mai_mai_n1111_));
  NO2        m1083(.A(mai_mai_n282_), .B(a), .Y(mai_mai_n1112_));
  INV        m1084(.A(mai_mai_n1035_), .Y(mai_mai_n1113_));
  NO2        m1085(.A(mai_mai_n1083_), .B(mai_mai_n476_), .Y(mai_mai_n1114_));
  NO2        m1086(.A(mai_mai_n89_), .B(g), .Y(mai_mai_n1115_));
  AOI210     m1087(.A0(mai_mai_n1115_), .A1(mai_mai_n1114_), .B0(mai_mai_n1067_), .Y(mai_mai_n1116_));
  OR2        m1088(.A(mai_mai_n1116_), .B(mai_mai_n1065_), .Y(mai_mai_n1117_));
  NA3        m1089(.A(mai_mai_n1117_), .B(mai_mai_n1113_), .C(mai_mai_n1111_), .Y(mai_mai_n1118_));
  NO4        m1090(.A(mai_mai_n1118_), .B(mai_mai_n1102_), .C(mai_mai_n819_), .D(mai_mai_n560_), .Y(mai_mai_n1119_));
  NA2        m1091(.A(c), .B(b), .Y(mai_mai_n1120_));
  NO2        m1092(.A(n), .B(mai_mai_n1120_), .Y(mai_mai_n1121_));
  OAI210     m1093(.A0(mai_mai_n859_), .A1(mai_mai_n832_), .B0(mai_mai_n408_), .Y(mai_mai_n1122_));
  OAI210     m1094(.A0(mai_mai_n1122_), .A1(mai_mai_n860_), .B0(mai_mai_n1121_), .Y(mai_mai_n1123_));
  NAi21      m1095(.An(mai_mai_n416_), .B(mai_mai_n1121_), .Y(mai_mai_n1124_));
  NA3        m1096(.A(mai_mai_n422_), .B(mai_mai_n553_), .C(f), .Y(mai_mai_n1125_));
  OAI210     m1097(.A0(mai_mai_n542_), .A1(mai_mai_n39_), .B0(mai_mai_n1112_), .Y(mai_mai_n1126_));
  NA3        m1098(.A(mai_mai_n1126_), .B(mai_mai_n1125_), .C(mai_mai_n1124_), .Y(mai_mai_n1127_));
  INV        m1099(.A(g), .Y(mai_mai_n1128_));
  NAi21      m1100(.An(f), .B(d), .Y(mai_mai_n1129_));
  NO2        m1101(.A(mai_mai_n1129_), .B(mai_mai_n1087_), .Y(mai_mai_n1130_));
  INV        m1102(.A(mai_mai_n1130_), .Y(mai_mai_n1131_));
  AOI210     m1103(.A0(mai_mai_n1128_), .A1(mai_mai_n290_), .B0(mai_mai_n1131_), .Y(mai_mai_n1132_));
  AOI210     m1104(.A0(mai_mai_n1132_), .A1(mai_mai_n115_), .B0(mai_mai_n1127_), .Y(mai_mai_n1133_));
  NA2        m1105(.A(mai_mai_n462_), .B(f), .Y(mai_mai_n1134_));
  NO2        m1106(.A(mai_mai_n186_), .B(mai_mai_n239_), .Y(mai_mai_n1135_));
  NA2        m1107(.A(mai_mai_n1135_), .B(m), .Y(mai_mai_n1136_));
  AOI210     m1108(.A0(mai_mai_n66_), .A1(mai_mai_n1134_), .B0(mai_mai_n1136_), .Y(mai_mai_n1137_));
  NA2        m1109(.A(mai_mai_n555_), .B(mai_mai_n403_), .Y(mai_mai_n1138_));
  NA2        m1110(.A(mai_mai_n441_), .B(mai_mai_n1130_), .Y(mai_mai_n1139_));
  NO2        m1111(.A(mai_mai_n368_), .B(mai_mai_n367_), .Y(mai_mai_n1140_));
  AOI210     m1112(.A0(mai_mai_n1135_), .A1(mai_mai_n424_), .B0(mai_mai_n952_), .Y(mai_mai_n1141_));
  NAi41      m1113(.An(mai_mai_n1140_), .B(mai_mai_n1141_), .C(mai_mai_n1139_), .D(mai_mai_n1138_), .Y(mai_mai_n1142_));
  NO2        m1114(.A(mai_mai_n1142_), .B(mai_mai_n1137_), .Y(mai_mai_n1143_));
  NA4        m1115(.A(mai_mai_n1143_), .B(mai_mai_n1133_), .C(mai_mai_n1123_), .D(mai_mai_n1119_), .Y(mai00));
  NA2        m1116(.A(mai_mai_n296_), .B(mai_mai_n219_), .Y(mai_mai_n1145_));
  NO2        m1117(.A(mai_mai_n1145_), .B(mai_mai_n574_), .Y(mai_mai_n1146_));
  AOI210     m1118(.A0(mai_mai_n893_), .A1(mai_mai_n935_), .B0(mai_mai_n1104_), .Y(mai_mai_n1147_));
  NO3        m1119(.A(mai_mai_n1080_), .B(mai_mai_n952_), .C(mai_mai_n707_), .Y(mai_mai_n1148_));
  NA3        m1120(.A(mai_mai_n1148_), .B(mai_mai_n1147_), .C(mai_mai_n994_), .Y(mai_mai_n1149_));
  NA2        m1121(.A(mai_mai_n502_), .B(f), .Y(mai_mai_n1150_));
  OAI210     m1122(.A0(mai_mai_n1001_), .A1(mai_mai_n40_), .B0(mai_mai_n643_), .Y(mai_mai_n1151_));
  NA3        m1123(.A(mai_mai_n1151_), .B(mai_mai_n260_), .C(n), .Y(mai_mai_n1152_));
  AOI210     m1124(.A0(mai_mai_n1152_), .A1(mai_mai_n1150_), .B0(mai_mai_n1038_), .Y(mai_mai_n1153_));
  NO4        m1125(.A(mai_mai_n1153_), .B(mai_mai_n1149_), .C(mai_mai_n1146_), .D(mai_mai_n1059_), .Y(mai_mai_n1154_));
  NA3        m1126(.A(mai_mai_n170_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(d), .B(b), .Y(mai_mai_n1156_));
  NOi31      m1128(.An(n), .B(m), .C(i), .Y(mai_mai_n1157_));
  NA3        m1129(.A(mai_mai_n1157_), .B(mai_mai_n646_), .C(mai_mai_n51_), .Y(mai_mai_n1158_));
  OAI210     m1130(.A0(mai_mai_n1156_), .A1(mai_mai_n1155_), .B0(mai_mai_n1158_), .Y(mai_mai_n1159_));
  INV        m1131(.A(mai_mai_n573_), .Y(mai_mai_n1160_));
  NO4        m1132(.A(mai_mai_n1160_), .B(mai_mai_n1159_), .C(mai_mai_n1140_), .D(mai_mai_n914_), .Y(mai_mai_n1161_));
  NO4        m1133(.A(mai_mai_n479_), .B(mai_mai_n351_), .C(mai_mai_n1120_), .D(mai_mai_n59_), .Y(mai_mai_n1162_));
  NA3        m1134(.A(mai_mai_n380_), .B(mai_mai_n226_), .C(g), .Y(mai_mai_n1163_));
  OA220      m1135(.A0(mai_mai_n1163_), .A1(mai_mai_n1156_), .B0(mai_mai_n381_), .B1(mai_mai_n137_), .Y(mai_mai_n1164_));
  NO2        m1136(.A(h), .B(g), .Y(mai_mai_n1165_));
  NA4        m1137(.A(mai_mai_n491_), .B(mai_mai_n460_), .C(mai_mai_n1165_), .D(mai_mai_n1027_), .Y(mai_mai_n1166_));
  OAI220     m1138(.A0(mai_mai_n519_), .A1(mai_mai_n594_), .B0(mai_mai_n94_), .B1(mai_mai_n93_), .Y(mai_mai_n1167_));
  AOI220     m1139(.A0(mai_mai_n1167_), .A1(mai_mai_n528_), .B0(mai_mai_n940_), .B1(mai_mai_n572_), .Y(mai_mai_n1168_));
  AOI220     m1140(.A0(mai_mai_n314_), .A1(mai_mai_n249_), .B0(mai_mai_n181_), .B1(mai_mai_n151_), .Y(mai_mai_n1169_));
  NA4        m1141(.A(mai_mai_n1169_), .B(mai_mai_n1168_), .C(mai_mai_n1166_), .D(mai_mai_n1164_), .Y(mai_mai_n1170_));
  NO3        m1142(.A(mai_mai_n1170_), .B(mai_mai_n1162_), .C(mai_mai_n267_), .Y(mai_mai_n1171_));
  INV        m1143(.A(mai_mai_n318_), .Y(mai_mai_n1172_));
  AOI210     m1144(.A0(mai_mai_n249_), .A1(mai_mai_n341_), .B0(mai_mai_n575_), .Y(mai_mai_n1173_));
  NA3        m1145(.A(mai_mai_n1173_), .B(mai_mai_n1172_), .C(mai_mai_n157_), .Y(mai_mai_n1174_));
  NO2        m1146(.A(mai_mai_n241_), .B(mai_mai_n185_), .Y(mai_mai_n1175_));
  NA2        m1147(.A(mai_mai_n1175_), .B(mai_mai_n422_), .Y(mai_mai_n1176_));
  NA3        m1148(.A(mai_mai_n183_), .B(mai_mai_n114_), .C(g), .Y(mai_mai_n1177_));
  NA3        m1149(.A(mai_mai_n460_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1178_));
  NOi31      m1150(.An(j), .B(mai_mai_n1178_), .C(mai_mai_n1177_), .Y(mai_mai_n1179_));
  NAi31      m1151(.An(mai_mai_n190_), .B(mai_mai_n856_), .C(mai_mai_n460_), .Y(mai_mai_n1180_));
  NAi31      m1152(.An(mai_mai_n1179_), .B(mai_mai_n1180_), .C(mai_mai_n1176_), .Y(mai_mai_n1181_));
  NO2        m1153(.A(mai_mai_n276_), .B(mai_mai_n75_), .Y(mai_mai_n1182_));
  NO3        m1154(.A(mai_mai_n421_), .B(mai_mai_n830_), .C(n), .Y(mai_mai_n1183_));
  AOI210     m1155(.A0(mai_mai_n1183_), .A1(mai_mai_n1182_), .B0(mai_mai_n1074_), .Y(mai_mai_n1184_));
  NAi31      m1156(.An(mai_mai_n1041_), .B(mai_mai_n1184_), .C(mai_mai_n74_), .Y(mai_mai_n1185_));
  NO4        m1157(.A(mai_mai_n1185_), .B(mai_mai_n1181_), .C(mai_mai_n1174_), .D(mai_mai_n510_), .Y(mai_mai_n1186_));
  AN3        m1158(.A(mai_mai_n1186_), .B(mai_mai_n1171_), .C(mai_mai_n1161_), .Y(mai_mai_n1187_));
  NA2        m1159(.A(mai_mai_n528_), .B(mai_mai_n103_), .Y(mai_mai_n1188_));
  NA3        m1160(.A(mai_mai_n1105_), .B(mai_mai_n604_), .C(mai_mai_n459_), .Y(mai_mai_n1189_));
  NA4        m1161(.A(mai_mai_n1189_), .B(mai_mai_n556_), .C(mai_mai_n1188_), .D(mai_mai_n244_), .Y(mai_mai_n1190_));
  NA2        m1162(.A(mai_mai_n1099_), .B(mai_mai_n528_), .Y(mai_mai_n1191_));
  NA4        m1163(.A(mai_mai_n646_), .B(mai_mai_n210_), .C(mai_mai_n226_), .D(h), .Y(mai_mai_n1192_));
  NA3        m1164(.A(mai_mai_n1192_), .B(mai_mai_n1191_), .C(mai_mai_n293_), .Y(mai_mai_n1193_));
  OAI210     m1165(.A0(mai_mai_n458_), .A1(mai_mai_n121_), .B0(mai_mai_n862_), .Y(mai_mai_n1194_));
  AOI210     m1166(.A0(mai_mai_n555_), .A1(mai_mai_n403_), .B0(mai_mai_n1194_), .Y(mai_mai_n1195_));
  OR4        m1167(.A(mai_mai_n1038_), .B(mai_mai_n272_), .C(mai_mai_n228_), .D(e), .Y(mai_mai_n1196_));
  NO2        m1168(.A(mai_mai_n222_), .B(mai_mai_n219_), .Y(mai_mai_n1197_));
  NA2        m1169(.A(n), .B(e), .Y(mai_mai_n1198_));
  NO2        m1170(.A(mai_mai_n1198_), .B(mai_mai_n149_), .Y(mai_mai_n1199_));
  AOI220     m1171(.A0(mai_mai_n1199_), .A1(mai_mai_n274_), .B0(mai_mai_n843_), .B1(mai_mai_n1197_), .Y(mai_mai_n1200_));
  OAI210     m1172(.A0(mai_mai_n352_), .A1(mai_mai_n309_), .B0(mai_mai_n443_), .Y(mai_mai_n1201_));
  NA4        m1173(.A(mai_mai_n1201_), .B(mai_mai_n1200_), .C(mai_mai_n1196_), .D(mai_mai_n1195_), .Y(mai_mai_n1202_));
  AOI210     m1174(.A0(mai_mai_n1199_), .A1(mai_mai_n847_), .B0(mai_mai_n818_), .Y(mai_mai_n1203_));
  AOI220     m1175(.A0(mai_mai_n948_), .A1(mai_mai_n572_), .B0(mai_mai_n646_), .B1(mai_mai_n247_), .Y(mai_mai_n1204_));
  NO2        m1176(.A(mai_mai_n68_), .B(h), .Y(mai_mai_n1205_));
  NO3        m1177(.A(mai_mai_n1038_), .B(mai_mai_n1036_), .C(mai_mai_n722_), .Y(mai_mai_n1206_));
  OAI210     m1178(.A0(mai_mai_n1085_), .A1(mai_mai_n1206_), .B0(mai_mai_n1205_), .Y(mai_mai_n1207_));
  NA4        m1179(.A(mai_mai_n1207_), .B(mai_mai_n1204_), .C(mai_mai_n1203_), .D(mai_mai_n864_), .Y(mai_mai_n1208_));
  NO4        m1180(.A(mai_mai_n1208_), .B(mai_mai_n1202_), .C(mai_mai_n1193_), .D(mai_mai_n1190_), .Y(mai_mai_n1209_));
  NA2        m1181(.A(mai_mai_n833_), .B(mai_mai_n753_), .Y(mai_mai_n1210_));
  NA4        m1182(.A(mai_mai_n1210_), .B(mai_mai_n1209_), .C(mai_mai_n1187_), .D(mai_mai_n1154_), .Y(mai01));
  AN2        m1183(.A(mai_mai_n1017_), .B(mai_mai_n1015_), .Y(mai_mai_n1212_));
  NO4        m1184(.A(mai_mai_n802_), .B(mai_mai_n794_), .C(mai_mai_n470_), .D(mai_mai_n281_), .Y(mai_mai_n1213_));
  NA3        m1185(.A(mai_mai_n587_), .B(mai_mai_n1213_), .C(mai_mai_n1212_), .Y(mai_mai_n1214_));
  NA2        m1186(.A(mai_mai_n583_), .B(mai_mai_n92_), .Y(mai_mai_n1215_));
  NA2        m1187(.A(mai_mai_n954_), .B(c), .Y(mai_mai_n1216_));
  NA4        m1188(.A(mai_mai_n1216_), .B(mai_mai_n1215_), .C(mai_mai_n908_), .D(mai_mai_n329_), .Y(mai_mai_n1217_));
  NA2        m1189(.A(mai_mai_n702_), .B(mai_mai_n99_), .Y(mai_mai_n1218_));
  OAI220     m1190(.A0(mai_mai_n1218_), .A1(mai_mai_n1455_), .B0(mai_mai_n348_), .B1(mai_mai_n284_), .Y(mai_mai_n1219_));
  OAI210     m1191(.A0(mai_mai_n780_), .A1(mai_mai_n599_), .B0(mai_mai_n1192_), .Y(mai_mai_n1220_));
  AOI210     m1192(.A0(mai_mai_n1219_), .A1(mai_mai_n632_), .B0(mai_mai_n1220_), .Y(mai_mai_n1221_));
  OA220      m1193(.A0(mai_mai_n1457_), .A1(mai_mai_n580_), .B0(mai_mai_n658_), .B1(mai_mai_n365_), .Y(mai_mai_n1222_));
  NAi41      m1194(.An(mai_mai_n165_), .B(mai_mai_n1222_), .C(mai_mai_n1221_), .D(mai_mai_n892_), .Y(mai_mai_n1223_));
  NO3        m1195(.A(mai_mai_n781_), .B(mai_mai_n669_), .C(mai_mai_n505_), .Y(mai_mai_n1224_));
  NA4        m1196(.A(mai_mai_n702_), .B(mai_mai_n99_), .C(mai_mai_n45_), .D(mai_mai_n218_), .Y(mai_mai_n1225_));
  OA220      m1197(.A0(mai_mai_n1225_), .A1(mai_mai_n663_), .B0(mai_mai_n200_), .B1(mai_mai_n198_), .Y(mai_mai_n1226_));
  NA3        m1198(.A(mai_mai_n1226_), .B(mai_mai_n1224_), .C(mai_mai_n140_), .Y(mai_mai_n1227_));
  NO4        m1199(.A(mai_mai_n1227_), .B(mai_mai_n1223_), .C(mai_mai_n1217_), .D(mai_mai_n1214_), .Y(mai_mai_n1228_));
  NA2        m1200(.A(mai_mai_n1163_), .B(mai_mai_n211_), .Y(mai_mai_n1229_));
  OAI210     m1201(.A0(mai_mai_n1229_), .A1(mai_mai_n299_), .B0(mai_mai_n523_), .Y(mai_mai_n1230_));
  NA2        m1202(.A(mai_mai_n531_), .B(mai_mai_n390_), .Y(mai_mai_n1231_));
  AOI210     m1203(.A0(mai_mai_n586_), .A1(mai_mai_n580_), .B0(mai_mai_n1456_), .Y(mai_mai_n1232_));
  AOI210     m1204(.A0(mai_mai_n557_), .A1(mai_mai_n1231_), .B0(mai_mai_n1232_), .Y(mai_mai_n1233_));
  AOI210     m1205(.A0(mai_mai_n208_), .A1(mai_mai_n91_), .B0(mai_mai_n218_), .Y(mai_mai_n1234_));
  OAI210     m1206(.A0(mai_mai_n807_), .A1(mai_mai_n422_), .B0(mai_mai_n1234_), .Y(mai_mai_n1235_));
  AN3        m1207(.A(m), .B(l), .C(k), .Y(mai_mai_n1236_));
  OAI210     m1208(.A0(mai_mai_n354_), .A1(mai_mai_n34_), .B0(mai_mai_n1236_), .Y(mai_mai_n1237_));
  NA2        m1209(.A(mai_mai_n207_), .B(mai_mai_n34_), .Y(mai_mai_n1238_));
  AO210      m1210(.A0(mai_mai_n1238_), .A1(mai_mai_n1237_), .B0(mai_mai_n328_), .Y(mai_mai_n1239_));
  NA4        m1211(.A(mai_mai_n1239_), .B(mai_mai_n1235_), .C(mai_mai_n1233_), .D(mai_mai_n1230_), .Y(mai_mai_n1240_));
  AOI210     m1212(.A0(mai_mai_n592_), .A1(mai_mai_n120_), .B0(mai_mai_n597_), .Y(mai_mai_n1241_));
  OAI210     m1213(.A0(mai_mai_n1457_), .A1(mai_mai_n589_), .B0(mai_mai_n1241_), .Y(mai_mai_n1242_));
  NO3        m1214(.A(mai_mai_n817_), .B(mai_mai_n208_), .C(mai_mai_n401_), .Y(mai_mai_n1243_));
  NO2        m1215(.A(mai_mai_n1243_), .B(mai_mai_n952_), .Y(mai_mai_n1244_));
  OAI210     m1216(.A0(mai_mai_n1219_), .A1(mai_mai_n322_), .B0(mai_mai_n670_), .Y(mai_mai_n1245_));
  NA3        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1244_), .C(mai_mai_n784_), .Y(mai_mai_n1246_));
  NO3        m1218(.A(mai_mai_n1246_), .B(mai_mai_n1242_), .C(mai_mai_n1240_), .Y(mai_mai_n1247_));
  NA3        m1219(.A(mai_mai_n600_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1248_));
  NO2        m1220(.A(mai_mai_n1248_), .B(mai_mai_n208_), .Y(mai_mai_n1249_));
  AOI210     m1221(.A0(mai_mai_n498_), .A1(mai_mai_n58_), .B0(mai_mai_n1249_), .Y(mai_mai_n1250_));
  OR3        m1222(.A(mai_mai_n1218_), .B(mai_mai_n601_), .C(mai_mai_n1455_), .Y(mai_mai_n1251_));
  NA3        m1223(.A(g), .B(mai_mai_n76_), .C(i), .Y(mai_mai_n1252_));
  AOI210     m1224(.A0(mai_mai_n1252_), .A1(mai_mai_n1225_), .B0(mai_mai_n972_), .Y(mai_mai_n1253_));
  NO2        m1225(.A(mai_mai_n211_), .B(mai_mai_n113_), .Y(mai_mai_n1254_));
  NO3        m1226(.A(mai_mai_n1254_), .B(mai_mai_n1253_), .C(mai_mai_n1159_), .Y(mai_mai_n1255_));
  NA4        m1227(.A(mai_mai_n1255_), .B(mai_mai_n1251_), .C(mai_mai_n1250_), .D(mai_mai_n752_), .Y(mai_mai_n1256_));
  NO2        m1228(.A(mai_mai_n961_), .B(mai_mai_n234_), .Y(mai_mai_n1257_));
  NO2        m1229(.A(mai_mai_n962_), .B(mai_mai_n550_), .Y(mai_mai_n1258_));
  OAI210     m1230(.A0(mai_mai_n1258_), .A1(mai_mai_n1257_), .B0(mai_mai_n336_), .Y(mai_mai_n1259_));
  NA2        m1231(.A(mai_mai_n567_), .B(mai_mai_n565_), .Y(mai_mai_n1260_));
  NO3        m1232(.A(mai_mai_n81_), .B(mai_mai_n297_), .C(mai_mai_n45_), .Y(mai_mai_n1261_));
  NA2        m1233(.A(mai_mai_n1261_), .B(mai_mai_n547_), .Y(mai_mai_n1262_));
  NA3        m1234(.A(mai_mai_n1262_), .B(mai_mai_n1260_), .C(mai_mai_n665_), .Y(mai_mai_n1263_));
  OR2        m1235(.A(mai_mai_n1163_), .B(mai_mai_n1156_), .Y(mai_mai_n1264_));
  NO2        m1236(.A(mai_mai_n365_), .B(mai_mai_n73_), .Y(mai_mai_n1265_));
  AOI210     m1237(.A0(mai_mai_n727_), .A1(mai_mai_n115_), .B0(mai_mai_n1265_), .Y(mai_mai_n1266_));
  NA2        m1238(.A(mai_mai_n1261_), .B(c), .Y(mai_mai_n1267_));
  NA4        m1239(.A(mai_mai_n1267_), .B(mai_mai_n1266_), .C(mai_mai_n1264_), .D(mai_mai_n383_), .Y(mai_mai_n1268_));
  NOi41      m1240(.An(mai_mai_n1259_), .B(mai_mai_n1268_), .C(mai_mai_n1263_), .D(mai_mai_n1256_), .Y(mai_mai_n1269_));
  NO2        m1241(.A(mai_mai_n133_), .B(mai_mai_n45_), .Y(mai_mai_n1270_));
  NO2        m1242(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1271_));
  AO220      m1243(.A0(mai_mai_n1271_), .A1(mai_mai_n619_), .B0(mai_mai_n1270_), .B1(mai_mai_n700_), .Y(mai_mai_n1272_));
  NA2        m1244(.A(mai_mai_n1272_), .B(mai_mai_n336_), .Y(mai_mai_n1273_));
  NA2        m1245(.A(mai_mai_n454_), .B(mai_mai_n137_), .Y(mai_mai_n1274_));
  NO3        m1246(.A(mai_mai_n1083_), .B(mai_mai_n180_), .C(mai_mai_n89_), .Y(mai_mai_n1275_));
  AOI220     m1247(.A0(mai_mai_n1275_), .A1(mai_mai_n1274_), .B0(mai_mai_n1261_), .B1(mai_mai_n965_), .Y(mai_mai_n1276_));
  NA2        m1248(.A(mai_mai_n1276_), .B(mai_mai_n1273_), .Y(mai_mai_n1277_));
  NO2        m1249(.A(mai_mai_n612_), .B(mai_mai_n611_), .Y(mai_mai_n1278_));
  NO4        m1250(.A(mai_mai_n1083_), .B(mai_mai_n1278_), .C(mai_mai_n178_), .D(mai_mai_n89_), .Y(mai_mai_n1279_));
  NO3        m1251(.A(mai_mai_n1279_), .B(mai_mai_n1277_), .C(mai_mai_n636_), .Y(mai_mai_n1280_));
  NA4        m1252(.A(mai_mai_n1280_), .B(mai_mai_n1269_), .C(mai_mai_n1247_), .D(mai_mai_n1228_), .Y(mai06));
  NO2        m1253(.A(mai_mai_n402_), .B(mai_mai_n554_), .Y(mai_mai_n1282_));
  OAI210     m1254(.A0(mai_mai_n115_), .A1(mai_mai_n268_), .B0(mai_mai_n1282_), .Y(mai_mai_n1283_));
  OR2        m1255(.A(mai_mai_n1463_), .B(mai_mai_n882_), .Y(mai_mai_n1284_));
  NA3        m1256(.A(mai_mai_n1284_), .B(mai_mai_n1283_), .C(mai_mai_n1259_), .Y(mai_mai_n1285_));
  NO3        m1257(.A(mai_mai_n1285_), .B(mai_mai_n1263_), .C(mai_mai_n259_), .Y(mai_mai_n1286_));
  NO2        m1258(.A(mai_mai_n297_), .B(mai_mai_n45_), .Y(mai_mai_n1287_));
  AOI210     m1259(.A0(mai_mai_n1287_), .A1(mai_mai_n966_), .B0(mai_mai_n1257_), .Y(mai_mai_n1288_));
  AOI210     m1260(.A0(mai_mai_n1287_), .A1(mai_mai_n551_), .B0(mai_mai_n1272_), .Y(mai_mai_n1289_));
  AOI210     m1261(.A0(mai_mai_n1289_), .A1(mai_mai_n1288_), .B0(mai_mai_n333_), .Y(mai_mai_n1290_));
  OAI210     m1262(.A0(mai_mai_n91_), .A1(mai_mai_n40_), .B0(mai_mai_n668_), .Y(mai_mai_n1291_));
  NA2        m1263(.A(mai_mai_n1291_), .B(mai_mai_n640_), .Y(mai_mai_n1292_));
  NO2        m1264(.A(mai_mai_n605_), .B(mai_mai_n1106_), .Y(mai_mai_n1293_));
  OAI210     m1265(.A0(mai_mai_n454_), .A1(mai_mai_n250_), .B0(mai_mai_n902_), .Y(mai_mai_n1294_));
  NO3        m1266(.A(mai_mai_n1294_), .B(mai_mai_n1293_), .C(mai_mai_n139_), .Y(mai_mai_n1295_));
  OR2        m1267(.A(mai_mai_n596_), .B(mai_mai_n595_), .Y(mai_mai_n1296_));
  NO2        m1268(.A(mai_mai_n1462_), .B(mai_mai_n138_), .Y(mai_mai_n1297_));
  AOI210     m1269(.A0(mai_mai_n1297_), .A1(mai_mai_n583_), .B0(mai_mai_n1296_), .Y(mai_mai_n1298_));
  NA3        m1270(.A(mai_mai_n1298_), .B(mai_mai_n1295_), .C(mai_mai_n1292_), .Y(mai_mai_n1299_));
  NO2        m1271(.A(mai_mai_n743_), .B(mai_mai_n364_), .Y(mai_mai_n1300_));
  NO3        m1272(.A(mai_mai_n670_), .B(mai_mai_n754_), .C(mai_mai_n632_), .Y(mai_mai_n1301_));
  NOi21      m1273(.An(mai_mai_n1300_), .B(mai_mai_n1301_), .Y(mai_mai_n1302_));
  AN2        m1274(.A(mai_mai_n948_), .B(c), .Y(mai_mai_n1303_));
  NO4        m1275(.A(mai_mai_n1303_), .B(mai_mai_n1302_), .C(mai_mai_n1299_), .D(mai_mai_n1290_), .Y(mai_mai_n1304_));
  NO2        m1276(.A(mai_mai_n801_), .B(mai_mai_n277_), .Y(mai_mai_n1305_));
  OAI220     m1277(.A0(mai_mai_n729_), .A1(mai_mai_n47_), .B0(mai_mai_n230_), .B1(mai_mai_n614_), .Y(mai_mai_n1306_));
  OAI210     m1278(.A0(mai_mai_n277_), .A1(c), .B0(mai_mai_n639_), .Y(mai_mai_n1307_));
  AOI220     m1279(.A0(mai_mai_n1307_), .A1(mai_mai_n1306_), .B0(mai_mai_n1305_), .B1(mai_mai_n268_), .Y(mai_mai_n1308_));
  NO3        m1280(.A(mai_mai_n246_), .B(mai_mai_n105_), .C(mai_mai_n282_), .Y(mai_mai_n1309_));
  NO2        m1281(.A(mai_mai_n693_), .B(mai_mai_n250_), .Y(mai_mai_n1310_));
  NO2        m1282(.A(mai_mai_n594_), .B(j), .Y(mai_mai_n1311_));
  NOi21      m1283(.An(mai_mai_n1311_), .B(mai_mai_n663_), .Y(mai_mai_n1312_));
  NO4        m1284(.A(mai_mai_n1312_), .B(mai_mai_n1310_), .C(mai_mai_n1309_), .D(mai_mai_n1109_), .Y(mai_mai_n1313_));
  NA4        m1285(.A(mai_mai_n792_), .B(mai_mai_n791_), .C(mai_mai_n431_), .D(mai_mai_n874_), .Y(mai_mai_n1314_));
  NAi31      m1286(.An(mai_mai_n743_), .B(mai_mai_n1314_), .C(mai_mai_n207_), .Y(mai_mai_n1315_));
  NA4        m1287(.A(mai_mai_n1315_), .B(mai_mai_n1313_), .C(mai_mai_n1308_), .D(mai_mai_n1204_), .Y(mai_mai_n1316_));
  OR2        m1288(.A(mai_mai_n780_), .B(mai_mai_n534_), .Y(mai_mai_n1317_));
  OR3        m1289(.A(mai_mai_n367_), .B(mai_mai_n230_), .C(mai_mai_n614_), .Y(mai_mai_n1318_));
  AOI210     m1290(.A0(mai_mai_n567_), .A1(mai_mai_n443_), .B0(mai_mai_n369_), .Y(mai_mai_n1319_));
  NA2        m1291(.A(mai_mai_n1311_), .B(mai_mai_n788_), .Y(mai_mai_n1320_));
  NA4        m1292(.A(mai_mai_n1320_), .B(mai_mai_n1319_), .C(mai_mai_n1318_), .D(mai_mai_n1317_), .Y(mai_mai_n1321_));
  AOI220     m1293(.A0(mai_mai_n1300_), .A1(mai_mai_n753_), .B0(mai_mai_n1297_), .B1(mai_mai_n240_), .Y(mai_mai_n1322_));
  AN2        m1294(.A(mai_mai_n923_), .B(mai_mai_n922_), .Y(mai_mai_n1323_));
  NO3        m1295(.A(mai_mai_n1323_), .B(mai_mai_n872_), .C(mai_mai_n494_), .Y(mai_mai_n1324_));
  NA3        m1296(.A(mai_mai_n1324_), .B(mai_mai_n1322_), .C(mai_mai_n1267_), .Y(mai_mai_n1325_));
  NAi21      m1297(.An(j), .B(i), .Y(mai_mai_n1326_));
  NO4        m1298(.A(mai_mai_n1278_), .B(mai_mai_n1326_), .C(mai_mai_n437_), .D(mai_mai_n237_), .Y(mai_mai_n1327_));
  NO4        m1299(.A(mai_mai_n1327_), .B(mai_mai_n1325_), .C(mai_mai_n1321_), .D(mai_mai_n1316_), .Y(mai_mai_n1328_));
  NA4        m1300(.A(mai_mai_n1328_), .B(mai_mai_n1304_), .C(mai_mai_n1286_), .D(mai_mai_n1280_), .Y(mai07));
  NAi32      m1301(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1330_));
  NO3        m1302(.A(mai_mai_n1330_), .B(g), .C(f), .Y(mai_mai_n1331_));
  OAI210     m1303(.A0(i), .A1(mai_mai_n475_), .B0(mai_mai_n1331_), .Y(mai_mai_n1332_));
  NAi21      m1304(.An(f), .B(c), .Y(mai_mai_n1333_));
  OR2        m1305(.A(e), .B(d), .Y(mai_mai_n1334_));
  OAI220     m1306(.A0(mai_mai_n1334_), .A1(mai_mai_n1333_), .B0(mai_mai_n624_), .B1(mai_mai_n319_), .Y(mai_mai_n1335_));
  NA3        m1307(.A(mai_mai_n1335_), .B(mai_mai_n1461_), .C(mai_mai_n183_), .Y(mai_mai_n1336_));
  NOi31      m1308(.An(n), .B(m), .C(b), .Y(mai_mai_n1337_));
  NO3        m1309(.A(mai_mai_n134_), .B(mai_mai_n445_), .C(h), .Y(mai_mai_n1338_));
  NA2        m1310(.A(mai_mai_n1336_), .B(mai_mai_n1332_), .Y(mai_mai_n1339_));
  NOi41      m1311(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1340_));
  NO2        m1312(.A(k), .B(i), .Y(mai_mai_n1341_));
  NA2        m1313(.A(mai_mai_n89_), .B(mai_mai_n45_), .Y(mai_mai_n1342_));
  NO2        m1314(.A(mai_mai_n1044_), .B(mai_mai_n437_), .Y(mai_mai_n1343_));
  NA3        m1315(.A(mai_mai_n1343_), .B(mai_mai_n1342_), .C(mai_mai_n219_), .Y(mai_mai_n1344_));
  NO2        m1316(.A(mai_mai_n1056_), .B(mai_mai_n305_), .Y(mai_mai_n1345_));
  NA2        m1317(.A(mai_mai_n535_), .B(mai_mai_n82_), .Y(mai_mai_n1346_));
  NA2        m1318(.A(mai_mai_n1346_), .B(mai_mai_n1344_), .Y(mai_mai_n1347_));
  NO2        m1319(.A(mai_mai_n1347_), .B(mai_mai_n1339_), .Y(mai_mai_n1348_));
  NO3        m1320(.A(e), .B(d), .C(c), .Y(mai_mai_n1349_));
  OAI210     m1321(.A0(mai_mai_n134_), .A1(mai_mai_n219_), .B0(mai_mai_n602_), .Y(mai_mai_n1350_));
  NA2        m1322(.A(mai_mai_n1350_), .B(mai_mai_n1349_), .Y(mai_mai_n1351_));
  NO2        m1323(.A(mai_mai_n1351_), .B(mai_mai_n219_), .Y(mai_mai_n1352_));
  NA3        m1324(.A(mai_mai_n690_), .B(mai_mai_n678_), .C(mai_mai_n114_), .Y(mai_mai_n1353_));
  NO2        m1325(.A(mai_mai_n1353_), .B(mai_mai_n45_), .Y(mai_mai_n1354_));
  NO2        m1326(.A(l), .B(k), .Y(mai_mai_n1355_));
  NO3        m1327(.A(mai_mai_n437_), .B(d), .C(c), .Y(mai_mai_n1356_));
  NO2        m1328(.A(mai_mai_n1354_), .B(mai_mai_n1352_), .Y(mai_mai_n1357_));
  NO2        m1329(.A(mai_mai_n150_), .B(h), .Y(mai_mai_n1358_));
  NO2        m1330(.A(g), .B(c), .Y(mai_mai_n1359_));
  NO2        m1331(.A(i), .B(h), .Y(mai_mai_n1360_));
  NA2        m1332(.A(mai_mai_n1129_), .B(h), .Y(mai_mai_n1361_));
  NA2        m1333(.A(mai_mai_n141_), .B(mai_mai_n226_), .Y(mai_mai_n1362_));
  NO2        m1334(.A(mai_mai_n1362_), .B(mai_mai_n1361_), .Y(mai_mai_n1363_));
  NOi31      m1335(.An(m), .B(n), .C(b), .Y(mai_mai_n1364_));
  NOi31      m1336(.An(f), .B(d), .C(c), .Y(mai_mai_n1365_));
  NA2        m1337(.A(mai_mai_n1365_), .B(mai_mai_n1364_), .Y(mai_mai_n1366_));
  INV        m1338(.A(mai_mai_n1366_), .Y(mai_mai_n1367_));
  NO2        m1339(.A(mai_mai_n1367_), .B(mai_mai_n1363_), .Y(mai_mai_n1368_));
  NA2        m1340(.A(mai_mai_n1077_), .B(mai_mai_n460_), .Y(mai_mai_n1369_));
  OAI210     m1341(.A0(mai_mai_n186_), .A1(mai_mai_n518_), .B0(mai_mai_n1052_), .Y(mai_mai_n1370_));
  AN2        m1342(.A(mai_mai_n1370_), .B(mai_mai_n1368_), .Y(mai_mai_n1371_));
  NA2        m1343(.A(mai_mai_n1356_), .B(mai_mai_n220_), .Y(mai_mai_n1372_));
  NA2        m1344(.A(mai_mai_n1084_), .B(mai_mai_n1369_), .Y(mai_mai_n1373_));
  NA2        m1345(.A(mai_mai_n1373_), .B(mai_mai_n1372_), .Y(mai_mai_n1374_));
  NO4        m1346(.A(mai_mai_n134_), .B(g), .C(f), .D(e), .Y(mai_mai_n1375_));
  NA2        m1347(.A(mai_mai_n1341_), .B(h), .Y(mai_mai_n1376_));
  OR2        m1348(.A(e), .B(a), .Y(mai_mai_n1377_));
  NA2        m1349(.A(mai_mai_n30_), .B(h), .Y(mai_mai_n1378_));
  NO2        m1350(.A(mai_mai_n1378_), .B(mai_mai_n1073_), .Y(mai_mai_n1379_));
  NA2        m1351(.A(mai_mai_n1340_), .B(mai_mai_n1355_), .Y(mai_mai_n1380_));
  INV        m1352(.A(mai_mai_n1380_), .Y(mai_mai_n1381_));
  OR3        m1353(.A(mai_mai_n534_), .B(mai_mai_n533_), .C(mai_mai_n114_), .Y(mai_mai_n1382_));
  NA2        m1354(.A(mai_mai_n1105_), .B(mai_mai_n401_), .Y(mai_mai_n1383_));
  NO3        m1355(.A(mai_mai_n1381_), .B(mai_mai_n1379_), .C(mai_mai_n1374_), .Y(mai_mai_n1384_));
  NA4        m1356(.A(mai_mai_n1384_), .B(mai_mai_n1371_), .C(mai_mai_n1357_), .D(mai_mai_n1348_), .Y(mai_mai_n1385_));
  NO2        m1357(.A(mai_mai_n385_), .B(j), .Y(mai_mai_n1386_));
  NAi41      m1358(.An(mai_mai_n1360_), .B(mai_mai_n1064_), .C(mai_mai_n171_), .D(mai_mai_n153_), .Y(mai_mai_n1387_));
  INV        m1359(.A(mai_mai_n1387_), .Y(mai_mai_n1388_));
  NA3        m1360(.A(g), .B(mai_mai_n1386_), .C(mai_mai_n162_), .Y(mai_mai_n1389_));
  INV        m1361(.A(mai_mai_n1389_), .Y(mai_mai_n1390_));
  NO3        m1362(.A(mai_mai_n743_), .B(mai_mai_n178_), .C(mai_mai_n404_), .Y(mai_mai_n1391_));
  NO3        m1363(.A(mai_mai_n1391_), .B(mai_mai_n1390_), .C(mai_mai_n1388_), .Y(mai_mai_n1392_));
  OR2        m1364(.A(n), .B(i), .Y(mai_mai_n1393_));
  OAI210     m1365(.A0(mai_mai_n1393_), .A1(mai_mai_n1063_), .B0(mai_mai_n49_), .Y(mai_mai_n1394_));
  AOI220     m1366(.A0(mai_mai_n1394_), .A1(mai_mai_n1165_), .B0(mai_mai_n822_), .B1(mai_mai_n199_), .Y(mai_mai_n1395_));
  NO2        m1367(.A(mai_mai_n1073_), .B(h), .Y(mai_mai_n1396_));
  NA2        m1368(.A(mai_mai_n183_), .B(mai_mai_n114_), .Y(mai_mai_n1397_));
  NOi21      m1369(.An(d), .B(f), .Y(mai_mai_n1398_));
  NA2        m1370(.A(mai_mai_n1395_), .B(mai_mai_n1392_), .Y(mai_mai_n1399_));
  NO3        m1371(.A(mai_mai_n1077_), .B(mai_mai_n1063_), .C(mai_mai_n40_), .Y(mai_mai_n1400_));
  NA2        m1372(.A(mai_mai_n1400_), .B(mai_mai_n1345_), .Y(mai_mai_n1401_));
  OAI210     m1373(.A0(mai_mai_n1375_), .A1(mai_mai_n1337_), .B0(mai_mai_n879_), .Y(mai_mai_n1402_));
  NA2        m1374(.A(mai_mai_n1402_), .B(mai_mai_n1401_), .Y(mai_mai_n1403_));
  NA2        m1375(.A(mai_mai_n1359_), .B(mai_mai_n1398_), .Y(mai_mai_n1404_));
  NO2        m1376(.A(mai_mai_n1404_), .B(m), .Y(mai_mai_n1405_));
  OAI220     m1377(.A0(mai_mai_n154_), .A1(mai_mai_n185_), .B0(mai_mai_n445_), .B1(g), .Y(mai_mai_n1406_));
  OAI210     m1378(.A0(mai_mai_n1406_), .A1(mai_mai_n112_), .B0(mai_mai_n1364_), .Y(mai_mai_n1407_));
  INV        m1379(.A(mai_mai_n1407_), .Y(mai_mai_n1408_));
  NO3        m1380(.A(mai_mai_n1408_), .B(mai_mai_n1405_), .C(mai_mai_n1403_), .Y(mai_mai_n1409_));
  NO2        m1381(.A(mai_mai_n1333_), .B(e), .Y(mai_mai_n1410_));
  NA2        m1382(.A(mai_mai_n1115_), .B(mai_mai_n628_), .Y(mai_mai_n1411_));
  NO2        m1383(.A(mai_mai_n1411_), .B(mai_mai_n439_), .Y(mai_mai_n1412_));
  NO3        m1384(.A(mai_mai_n1382_), .B(mai_mai_n348_), .C(a), .Y(mai_mai_n1413_));
  NO2        m1385(.A(mai_mai_n1413_), .B(mai_mai_n1412_), .Y(mai_mai_n1414_));
  NO2        m1386(.A(mai_mai_n185_), .B(c), .Y(mai_mai_n1415_));
  OAI210     m1387(.A0(mai_mai_n1415_), .A1(mai_mai_n1410_), .B0(mai_mai_n183_), .Y(mai_mai_n1416_));
  AOI220     m1388(.A0(mai_mai_n1416_), .A1(mai_mai_n1065_), .B0(mai_mai_n525_), .B1(mai_mai_n364_), .Y(mai_mai_n1417_));
  NA2        m1389(.A(mai_mai_n533_), .B(g), .Y(mai_mai_n1418_));
  NA2        m1390(.A(mai_mai_n1418_), .B(mai_mai_n1356_), .Y(mai_mai_n1419_));
  NO2        m1391(.A(mai_mai_n1377_), .B(f), .Y(mai_mai_n1420_));
  NO2        m1392(.A(mai_mai_n1419_), .B(mai_mai_n218_), .Y(mai_mai_n1421_));
  AOI210     m1393(.A0(mai_mai_n896_), .A1(mai_mai_n411_), .B0(mai_mai_n107_), .Y(mai_mai_n1422_));
  OR2        m1394(.A(mai_mai_n1422_), .B(mai_mai_n533_), .Y(mai_mai_n1423_));
  NA2        m1395(.A(mai_mai_n1420_), .B(mai_mai_n1342_), .Y(mai_mai_n1424_));
  OAI220     m1396(.A0(mai_mai_n1424_), .A1(mai_mai_n49_), .B0(mai_mai_n1423_), .B1(mai_mai_n178_), .Y(mai_mai_n1425_));
  NA2        m1397(.A(mai_mai_n1338_), .B(mai_mai_n186_), .Y(mai_mai_n1426_));
  NO2        m1398(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1427_));
  OAI210     m1399(.A0(mai_mai_n1377_), .A1(mai_mai_n858_), .B0(mai_mai_n475_), .Y(mai_mai_n1428_));
  OAI210     m1400(.A0(mai_mai_n1428_), .A1(mai_mai_n1088_), .B0(mai_mai_n1427_), .Y(mai_mai_n1429_));
  NO2        m1401(.A(m), .B(i), .Y(mai_mai_n1430_));
  NA2        m1402(.A(mai_mai_n1430_), .B(mai_mai_n1358_), .Y(mai_mai_n1431_));
  NA3        m1403(.A(mai_mai_n1431_), .B(mai_mai_n1429_), .C(mai_mai_n1426_), .Y(mai_mai_n1432_));
  NO4        m1404(.A(mai_mai_n1432_), .B(mai_mai_n1425_), .C(mai_mai_n1421_), .D(mai_mai_n1417_), .Y(mai_mai_n1433_));
  NA3        m1405(.A(mai_mai_n1433_), .B(mai_mai_n1414_), .C(mai_mai_n1409_), .Y(mai_mai_n1434_));
  OAI210     m1406(.A0(mai_mai_n579_), .A1(g), .B0(mai_mai_n189_), .Y(mai_mai_n1435_));
  NA2        m1407(.A(mai_mai_n1435_), .B(mai_mai_n1396_), .Y(mai_mai_n1436_));
  AOI210     m1408(.A0(mai_mai_n160_), .A1(mai_mai_n56_), .B0(mai_mai_n1410_), .Y(mai_mai_n1437_));
  NO2        m1409(.A(mai_mai_n1437_), .B(mai_mai_n1397_), .Y(mai_mai_n1438_));
  INV        m1410(.A(mai_mai_n1438_), .Y(mai_mai_n1439_));
  NA2        m1411(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1440_));
  NO2        m1412(.A(mai_mai_n1383_), .B(mai_mai_n1440_), .Y(mai_mai_n1441_));
  INV        m1413(.A(mai_mai_n1441_), .Y(mai_mai_n1442_));
  NA3        m1414(.A(mai_mai_n1442_), .B(mai_mai_n1439_), .C(mai_mai_n1436_), .Y(mai_mai_n1443_));
  OR4        m1415(.A(mai_mai_n1443_), .B(mai_mai_n1434_), .C(mai_mai_n1399_), .D(mai_mai_n1385_), .Y(mai04));
  NOi31      m1416(.An(mai_mai_n1375_), .B(mai_mai_n1376_), .C(mai_mai_n1038_), .Y(mai_mai_n1445_));
  NO4        m1417(.A(mai_mai_n272_), .B(mai_mai_n1028_), .C(mai_mai_n476_), .D(j), .Y(mai_mai_n1446_));
  OR3        m1418(.A(mai_mai_n1446_), .B(mai_mai_n1445_), .C(mai_mai_n1054_), .Y(mai_mai_n1447_));
  NO3        m1419(.A(mai_mai_n1342_), .B(mai_mai_n93_), .C(k), .Y(mai_mai_n1448_));
  AOI210     m1420(.A0(mai_mai_n1448_), .A1(mai_mai_n1049_), .B0(mai_mai_n1179_), .Y(mai_mai_n1449_));
  NA2        m1421(.A(mai_mai_n1449_), .B(mai_mai_n1207_), .Y(mai_mai_n1450_));
  NO4        m1422(.A(mai_mai_n1450_), .B(mai_mai_n1447_), .C(mai_mai_n1062_), .D(mai_mai_n1043_), .Y(mai_mai_n1451_));
  NA4        m1423(.A(mai_mai_n1451_), .B(mai_mai_n1117_), .C(mai_mai_n1103_), .D(mai_mai_n1091_), .Y(mai05));
  INV        m1424(.A(f), .Y(mai_mai_n1455_));
  INV        m1425(.A(k), .Y(mai_mai_n1456_));
  INV        m1426(.A(k), .Y(mai_mai_n1457_));
  INV        m1427(.A(mai_mai_n432_), .Y(mai_mai_n1458_));
  INV        m1428(.A(m), .Y(mai_mai_n1459_));
  INV        m1429(.A(m), .Y(mai_mai_n1460_));
  INV        m1430(.A(j), .Y(mai_mai_n1461_));
  INV        m1431(.A(m), .Y(mai_mai_n1462_));
  INV        m1432(.A(b), .Y(mai_mai_n1463_));
  INV        m1433(.A(b), .Y(mai_mai_n1464_));
  INV        m1434(.A(c), .Y(mai_mai_n1465_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NAi21      u0031(.An(i), .B(h), .Y(men_men_n60_));
  NAi31      u0032(.An(i), .B(l), .C(j), .Y(men_men_n61_));
  OAI220     u0033(.A0(men_men_n61_), .A1(men_men_n49_), .B0(men_men_n60_), .B1(men_men_n44_), .Y(men_men_n62_));
  NAi31      u0034(.An(d), .B(men_men_n62_), .C(men_men_n58_), .Y(men_men_n63_));
  NAi41      u0035(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n64_));
  NA2        u0036(.A(g), .B(f), .Y(men_men_n65_));
  NO2        u0037(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NAi21      u0038(.An(i), .B(j), .Y(men_men_n67_));
  NAi32      u0039(.An(n), .Bn(k), .C(m), .Y(men_men_n68_));
  NO2        u0040(.A(men_men_n68_), .B(men_men_n67_), .Y(men_men_n69_));
  NAi31      u0041(.An(l), .B(m), .C(k), .Y(men_men_n70_));
  NAi21      u0042(.An(e), .B(h), .Y(men_men_n71_));
  NAi41      u0043(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n73_));
  INV        u0045(.A(m), .Y(men_men_n74_));
  NOi21      u0046(.An(k), .B(l), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  AN4        u0048(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n77_));
  NOi31      u0049(.An(h), .B(g), .C(f), .Y(men_men_n78_));
  NA2        u0050(.A(men_men_n78_), .B(men_men_n77_), .Y(men_men_n79_));
  NAi32      u0051(.An(m), .Bn(k), .C(j), .Y(men_men_n80_));
  NOi32      u0052(.An(h), .Bn(g), .C(f), .Y(men_men_n81_));
  NA2        u0053(.A(men_men_n81_), .B(men_men_n77_), .Y(men_men_n82_));
  OA220      u0054(.A0(men_men_n82_), .A1(men_men_n80_), .B0(men_men_n79_), .B1(men_men_n76_), .Y(men_men_n83_));
  NA3        u0055(.A(men_men_n83_), .B(men_men_n73_), .C(men_men_n63_), .Y(men_men_n84_));
  INV        u0056(.A(n), .Y(men_men_n85_));
  NOi32      u0057(.An(e), .Bn(b), .C(d), .Y(men_men_n86_));
  NA2        u0058(.A(men_men_n86_), .B(men_men_n85_), .Y(men_men_n87_));
  INV        u0059(.A(j), .Y(men_men_n88_));
  AN3        u0060(.A(m), .B(k), .C(i), .Y(men_men_n89_));
  NA3        u0061(.A(men_men_n89_), .B(men_men_n88_), .C(g), .Y(men_men_n90_));
  NO2        u0062(.A(men_men_n90_), .B(f), .Y(men_men_n91_));
  NAi32      u0063(.An(g), .Bn(f), .C(h), .Y(men_men_n92_));
  NAi31      u0064(.An(j), .B(m), .C(l), .Y(men_men_n93_));
  NO2        u0065(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  NA2        u0066(.A(m), .B(l), .Y(men_men_n95_));
  NAi31      u0067(.An(k), .B(j), .C(g), .Y(men_men_n96_));
  NO3        u0068(.A(men_men_n96_), .B(men_men_n95_), .C(f), .Y(men_men_n97_));
  AN2        u0069(.A(j), .B(g), .Y(men_men_n98_));
  NOi32      u0070(.An(m), .Bn(l), .C(i), .Y(men_men_n99_));
  NOi21      u0071(.An(g), .B(i), .Y(men_men_n100_));
  NOi32      u0072(.An(m), .Bn(j), .C(k), .Y(men_men_n101_));
  AOI220     u0073(.A0(men_men_n101_), .A1(men_men_n100_), .B0(men_men_n99_), .B1(men_men_n98_), .Y(men_men_n102_));
  NO2        u0074(.A(men_men_n102_), .B(f), .Y(men_men_n103_));
  NO4        u0075(.A(men_men_n103_), .B(men_men_n97_), .C(men_men_n94_), .D(men_men_n91_), .Y(men_men_n104_));
  NAi41      u0076(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n105_));
  AN2        u0077(.A(e), .B(b), .Y(men_men_n106_));
  NOi31      u0078(.An(c), .B(h), .C(f), .Y(men_men_n107_));
  NA2        u0079(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NO3        u0080(.A(men_men_n108_), .B(men_men_n105_), .C(g), .Y(men_men_n109_));
  NOi21      u0081(.An(g), .B(f), .Y(men_men_n110_));
  NOi21      u0082(.An(i), .B(h), .Y(men_men_n111_));
  NA3        u0083(.A(men_men_n111_), .B(men_men_n110_), .C(men_men_n36_), .Y(men_men_n112_));
  INV        u0084(.A(a), .Y(men_men_n113_));
  NA2        u0085(.A(men_men_n106_), .B(men_men_n113_), .Y(men_men_n114_));
  INV        u0086(.A(l), .Y(men_men_n115_));
  NOi21      u0087(.An(m), .B(n), .Y(men_men_n116_));
  AN2        u0088(.A(k), .B(h), .Y(men_men_n117_));
  NO2        u0089(.A(men_men_n112_), .B(men_men_n87_), .Y(men_men_n118_));
  INV        u0090(.A(b), .Y(men_men_n119_));
  NA2        u0091(.A(l), .B(j), .Y(men_men_n120_));
  AN2        u0092(.A(k), .B(i), .Y(men_men_n121_));
  NA2        u0093(.A(men_men_n121_), .B(men_men_n120_), .Y(men_men_n122_));
  NA2        u0094(.A(g), .B(e), .Y(men_men_n123_));
  NOi32      u0095(.An(c), .Bn(a), .C(d), .Y(men_men_n124_));
  NA2        u0096(.A(men_men_n124_), .B(men_men_n116_), .Y(men_men_n125_));
  NO4        u0097(.A(men_men_n125_), .B(men_men_n123_), .C(men_men_n122_), .D(men_men_n119_), .Y(men_men_n126_));
  NO3        u0098(.A(men_men_n126_), .B(men_men_n118_), .C(men_men_n109_), .Y(men_men_n127_));
  OAI210     u0099(.A0(men_men_n104_), .A1(men_men_n87_), .B0(men_men_n127_), .Y(men_men_n128_));
  NOi31      u0100(.An(k), .B(m), .C(j), .Y(men_men_n129_));
  NA3        u0101(.A(men_men_n129_), .B(men_men_n78_), .C(men_men_n77_), .Y(men_men_n130_));
  NOi31      u0102(.An(k), .B(m), .C(i), .Y(men_men_n131_));
  NA3        u0103(.A(men_men_n131_), .B(men_men_n81_), .C(men_men_n77_), .Y(men_men_n132_));
  NA2        u0104(.A(men_men_n132_), .B(men_men_n130_), .Y(men_men_n133_));
  NOi32      u0105(.An(f), .Bn(b), .C(e), .Y(men_men_n134_));
  NAi21      u0106(.An(g), .B(h), .Y(men_men_n135_));
  NAi21      u0107(.An(m), .B(n), .Y(men_men_n136_));
  NAi21      u0108(.An(j), .B(k), .Y(men_men_n137_));
  NO3        u0109(.A(men_men_n137_), .B(men_men_n136_), .C(men_men_n135_), .Y(men_men_n138_));
  NAi41      u0110(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n139_));
  NAi31      u0111(.An(j), .B(k), .C(h), .Y(men_men_n140_));
  NO3        u0112(.A(men_men_n140_), .B(men_men_n139_), .C(men_men_n136_), .Y(men_men_n141_));
  AOI210     u0113(.A0(men_men_n138_), .A1(men_men_n134_), .B0(men_men_n141_), .Y(men_men_n142_));
  NO2        u0114(.A(k), .B(j), .Y(men_men_n143_));
  INV        u0115(.A(men_men_n136_), .Y(men_men_n144_));
  AN2        u0116(.A(k), .B(j), .Y(men_men_n145_));
  NAi21      u0117(.An(c), .B(b), .Y(men_men_n146_));
  NA2        u0118(.A(f), .B(d), .Y(men_men_n147_));
  NO4        u0119(.A(men_men_n147_), .B(men_men_n146_), .C(men_men_n145_), .D(men_men_n135_), .Y(men_men_n148_));
  NA2        u0120(.A(h), .B(c), .Y(men_men_n149_));
  NAi31      u0121(.An(f), .B(e), .C(b), .Y(men_men_n150_));
  NA2        u0122(.A(men_men_n148_), .B(men_men_n144_), .Y(men_men_n151_));
  NA2        u0123(.A(d), .B(b), .Y(men_men_n152_));
  NAi21      u0124(.An(e), .B(f), .Y(men_men_n153_));
  NO2        u0125(.A(men_men_n153_), .B(men_men_n152_), .Y(men_men_n154_));
  NA2        u0126(.A(b), .B(a), .Y(men_men_n155_));
  NAi21      u0127(.An(e), .B(g), .Y(men_men_n156_));
  NAi21      u0128(.An(c), .B(d), .Y(men_men_n157_));
  NAi31      u0129(.An(l), .B(k), .C(h), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n136_), .B(men_men_n158_), .Y(men_men_n159_));
  NA2        u0131(.A(men_men_n159_), .B(men_men_n154_), .Y(men_men_n160_));
  NAi41      u0132(.An(men_men_n133_), .B(men_men_n160_), .C(men_men_n151_), .D(men_men_n142_), .Y(men_men_n161_));
  NAi31      u0133(.An(e), .B(f), .C(b), .Y(men_men_n162_));
  NOi21      u0134(.An(g), .B(d), .Y(men_men_n163_));
  NO2        u0135(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  NOi21      u0136(.An(h), .B(i), .Y(men_men_n165_));
  NOi21      u0137(.An(k), .B(m), .Y(men_men_n166_));
  NA3        u0138(.A(men_men_n166_), .B(men_men_n165_), .C(n), .Y(men_men_n167_));
  NOi21      u0139(.An(men_men_n164_), .B(men_men_n167_), .Y(men_men_n168_));
  NOi21      u0140(.An(h), .B(g), .Y(men_men_n169_));
  NO2        u0141(.A(men_men_n147_), .B(men_men_n146_), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n169_), .Y(men_men_n171_));
  NAi31      u0143(.An(l), .B(j), .C(h), .Y(men_men_n172_));
  NO2        u0144(.A(men_men_n172_), .B(men_men_n49_), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n66_), .Y(men_men_n174_));
  NOi32      u0146(.An(n), .Bn(k), .C(m), .Y(men_men_n175_));
  NA2        u0147(.A(l), .B(i), .Y(men_men_n176_));
  NA2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  OAI210     u0149(.A0(men_men_n177_), .A1(men_men_n171_), .B0(men_men_n174_), .Y(men_men_n178_));
  NAi31      u0150(.An(d), .B(f), .C(c), .Y(men_men_n179_));
  NAi31      u0151(.An(e), .B(f), .C(c), .Y(men_men_n180_));
  NA2        u0152(.A(j), .B(h), .Y(men_men_n181_));
  OR3        u0153(.A(n), .B(m), .C(k), .Y(men_men_n182_));
  NAi32      u0154(.An(m), .Bn(k), .C(n), .Y(men_men_n183_));
  NO2        u0155(.A(men_men_n183_), .B(men_men_n181_), .Y(men_men_n184_));
  NA2        u0156(.A(men_men_n184_), .B(men_men_n164_), .Y(men_men_n185_));
  NO2        u0157(.A(n), .B(m), .Y(men_men_n186_));
  NA2        u0158(.A(men_men_n186_), .B(men_men_n50_), .Y(men_men_n187_));
  NAi21      u0159(.An(f), .B(e), .Y(men_men_n188_));
  NA2        u0160(.A(d), .B(c), .Y(men_men_n189_));
  NO2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NOi21      u0162(.An(men_men_n190_), .B(men_men_n187_), .Y(men_men_n191_));
  NAi31      u0163(.An(m), .B(n), .C(b), .Y(men_men_n192_));
  NA2        u0164(.A(k), .B(i), .Y(men_men_n193_));
  NAi21      u0165(.An(h), .B(f), .Y(men_men_n194_));
  NO2        u0166(.A(men_men_n194_), .B(men_men_n193_), .Y(men_men_n195_));
  NO2        u0167(.A(men_men_n192_), .B(men_men_n157_), .Y(men_men_n196_));
  NA2        u0168(.A(men_men_n196_), .B(men_men_n195_), .Y(men_men_n197_));
  NOi32      u0169(.An(f), .Bn(c), .C(d), .Y(men_men_n198_));
  NOi32      u0170(.An(f), .Bn(c), .C(e), .Y(men_men_n199_));
  NO2        u0171(.A(men_men_n199_), .B(men_men_n198_), .Y(men_men_n200_));
  NO3        u0172(.A(n), .B(m), .C(j), .Y(men_men_n201_));
  NA2        u0173(.A(men_men_n201_), .B(men_men_n117_), .Y(men_men_n202_));
  NAi31      u0174(.An(men_men_n191_), .B(men_men_n197_), .C(men_men_n185_), .Y(men_men_n203_));
  OR4        u0175(.A(men_men_n203_), .B(men_men_n178_), .C(men_men_n168_), .D(men_men_n161_), .Y(men_men_n204_));
  NO4        u0176(.A(men_men_n204_), .B(men_men_n128_), .C(men_men_n84_), .D(men_men_n55_), .Y(men_men_n205_));
  NA3        u0177(.A(m), .B(men_men_n115_), .C(j), .Y(men_men_n206_));
  NAi31      u0178(.An(n), .B(h), .C(g), .Y(men_men_n207_));
  NO2        u0179(.A(men_men_n207_), .B(men_men_n206_), .Y(men_men_n208_));
  NOi32      u0180(.An(m), .Bn(k), .C(l), .Y(men_men_n209_));
  NA3        u0181(.A(men_men_n209_), .B(men_men_n88_), .C(g), .Y(men_men_n210_));
  NO2        u0182(.A(men_men_n210_), .B(n), .Y(men_men_n211_));
  NOi21      u0183(.An(k), .B(j), .Y(men_men_n212_));
  NA4        u0184(.A(men_men_n212_), .B(men_men_n116_), .C(i), .D(g), .Y(men_men_n213_));
  AN2        u0185(.A(i), .B(g), .Y(men_men_n214_));
  NA3        u0186(.A(men_men_n75_), .B(men_men_n214_), .C(men_men_n116_), .Y(men_men_n215_));
  NA2        u0187(.A(men_men_n215_), .B(men_men_n213_), .Y(men_men_n216_));
  NO3        u0188(.A(men_men_n216_), .B(men_men_n211_), .C(men_men_n208_), .Y(men_men_n217_));
  NAi41      u0189(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n218_));
  INV        u0190(.A(men_men_n218_), .Y(men_men_n219_));
  INV        u0191(.A(f), .Y(men_men_n220_));
  INV        u0192(.A(g), .Y(men_men_n221_));
  NOi31      u0193(.An(i), .B(j), .C(h), .Y(men_men_n222_));
  NOi21      u0194(.An(l), .B(m), .Y(men_men_n223_));
  NA2        u0195(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n224_));
  NO3        u0196(.A(men_men_n224_), .B(men_men_n221_), .C(men_men_n220_), .Y(men_men_n225_));
  NA2        u0197(.A(men_men_n225_), .B(men_men_n219_), .Y(men_men_n226_));
  OAI210     u0198(.A0(men_men_n217_), .A1(men_men_n32_), .B0(men_men_n226_), .Y(men_men_n227_));
  NOi21      u0199(.An(n), .B(m), .Y(men_men_n228_));
  NA2        u0200(.A(i), .B(men_men_n228_), .Y(men_men_n229_));
  OA220      u0201(.A0(men_men_n229_), .A1(men_men_n108_), .B0(men_men_n80_), .B1(men_men_n79_), .Y(men_men_n230_));
  NAi21      u0202(.An(j), .B(h), .Y(men_men_n231_));
  XN2        u0203(.A(i), .B(h), .Y(men_men_n232_));
  NA2        u0204(.A(men_men_n232_), .B(men_men_n231_), .Y(men_men_n233_));
  NOi31      u0205(.An(k), .B(n), .C(m), .Y(men_men_n234_));
  NOi31      u0206(.An(men_men_n234_), .B(men_men_n189_), .C(men_men_n188_), .Y(men_men_n235_));
  NA2        u0207(.A(men_men_n235_), .B(men_men_n233_), .Y(men_men_n236_));
  NAi31      u0208(.An(f), .B(e), .C(c), .Y(men_men_n237_));
  NA4        u0209(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n238_));
  NAi32      u0210(.An(m), .Bn(i), .C(k), .Y(men_men_n239_));
  NO3        u0211(.A(men_men_n239_), .B(men_men_n92_), .C(men_men_n238_), .Y(men_men_n240_));
  INV        u0212(.A(men_men_n240_), .Y(men_men_n241_));
  NAi21      u0213(.An(n), .B(a), .Y(men_men_n242_));
  NO2        u0214(.A(men_men_n242_), .B(men_men_n152_), .Y(men_men_n243_));
  NAi41      u0215(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n244_));
  NO2        u0216(.A(men_men_n244_), .B(e), .Y(men_men_n245_));
  NO3        u0217(.A(men_men_n153_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n246_));
  OAI210     u0218(.A0(men_men_n246_), .A1(men_men_n245_), .B0(men_men_n243_), .Y(men_men_n247_));
  AN4        u0219(.A(men_men_n247_), .B(men_men_n241_), .C(men_men_n236_), .D(men_men_n230_), .Y(men_men_n248_));
  OR2        u0220(.A(h), .B(g), .Y(men_men_n249_));
  NO2        u0221(.A(men_men_n249_), .B(men_men_n105_), .Y(men_men_n250_));
  NA2        u0222(.A(men_men_n250_), .B(men_men_n134_), .Y(men_men_n251_));
  NAi41      u0223(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n252_));
  NO2        u0224(.A(men_men_n252_), .B(men_men_n220_), .Y(men_men_n253_));
  NA2        u0225(.A(men_men_n166_), .B(men_men_n111_), .Y(men_men_n254_));
  NAi21      u0226(.An(men_men_n254_), .B(men_men_n253_), .Y(men_men_n255_));
  NO2        u0227(.A(n), .B(a), .Y(men_men_n256_));
  NAi31      u0228(.An(men_men_n244_), .B(men_men_n256_), .C(men_men_n106_), .Y(men_men_n257_));
  AN2        u0229(.A(men_men_n257_), .B(men_men_n255_), .Y(men_men_n258_));
  NAi21      u0230(.An(h), .B(i), .Y(men_men_n259_));
  NA2        u0231(.A(men_men_n186_), .B(k), .Y(men_men_n260_));
  NO2        u0232(.A(men_men_n260_), .B(men_men_n259_), .Y(men_men_n261_));
  NA2        u0233(.A(men_men_n258_), .B(men_men_n251_), .Y(men_men_n262_));
  NOi21      u0234(.An(g), .B(e), .Y(men_men_n263_));
  NO2        u0235(.A(men_men_n72_), .B(men_men_n74_), .Y(men_men_n264_));
  NA2        u0236(.A(men_men_n264_), .B(men_men_n263_), .Y(men_men_n265_));
  NOi32      u0237(.An(l), .Bn(j), .C(i), .Y(men_men_n266_));
  AOI210     u0238(.A0(men_men_n75_), .A1(men_men_n88_), .B0(men_men_n266_), .Y(men_men_n267_));
  NO2        u0239(.A(men_men_n259_), .B(men_men_n44_), .Y(men_men_n268_));
  NAi21      u0240(.An(f), .B(g), .Y(men_men_n269_));
  NO2        u0241(.A(men_men_n269_), .B(men_men_n64_), .Y(men_men_n270_));
  NO2        u0242(.A(men_men_n68_), .B(men_men_n120_), .Y(men_men_n271_));
  AOI220     u0243(.A0(men_men_n271_), .A1(men_men_n270_), .B0(men_men_n268_), .B1(men_men_n66_), .Y(men_men_n272_));
  OAI210     u0244(.A0(men_men_n267_), .A1(men_men_n265_), .B0(men_men_n272_), .Y(men_men_n273_));
  NO3        u0245(.A(men_men_n137_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n274_));
  NOi41      u0246(.An(men_men_n248_), .B(men_men_n273_), .C(men_men_n262_), .D(men_men_n227_), .Y(men_men_n275_));
  NO4        u0247(.A(men_men_n208_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n276_));
  NO2        u0248(.A(men_men_n276_), .B(men_men_n114_), .Y(men_men_n277_));
  NA3        u0249(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n278_));
  NAi21      u0250(.An(h), .B(g), .Y(men_men_n279_));
  OR4        u0251(.A(men_men_n279_), .B(men_men_n278_), .C(men_men_n229_), .D(e), .Y(men_men_n280_));
  NO2        u0252(.A(men_men_n254_), .B(men_men_n269_), .Y(men_men_n281_));
  NA2        u0253(.A(men_men_n281_), .B(men_men_n77_), .Y(men_men_n282_));
  NAi31      u0254(.An(g), .B(k), .C(h), .Y(men_men_n283_));
  NO3        u0255(.A(men_men_n136_), .B(men_men_n283_), .C(l), .Y(men_men_n284_));
  NAi31      u0256(.An(e), .B(d), .C(a), .Y(men_men_n285_));
  NA2        u0257(.A(men_men_n284_), .B(men_men_n134_), .Y(men_men_n286_));
  NA3        u0258(.A(men_men_n286_), .B(men_men_n282_), .C(men_men_n280_), .Y(men_men_n287_));
  NA4        u0259(.A(men_men_n166_), .B(men_men_n81_), .C(men_men_n77_), .D(men_men_n120_), .Y(men_men_n288_));
  NA3        u0260(.A(men_men_n166_), .B(men_men_n165_), .C(men_men_n85_), .Y(men_men_n289_));
  NO2        u0261(.A(men_men_n289_), .B(men_men_n200_), .Y(men_men_n290_));
  NOi21      u0262(.An(men_men_n288_), .B(men_men_n290_), .Y(men_men_n291_));
  NA3        u0263(.A(e), .B(c), .C(b), .Y(men_men_n292_));
  NO2        u0264(.A(d), .B(men_men_n292_), .Y(men_men_n293_));
  NAi32      u0265(.An(k), .Bn(i), .C(j), .Y(men_men_n294_));
  NAi31      u0266(.An(h), .B(l), .C(i), .Y(men_men_n295_));
  NA3        u0267(.A(men_men_n295_), .B(men_men_n294_), .C(men_men_n172_), .Y(men_men_n296_));
  NOi21      u0268(.An(men_men_n296_), .B(men_men_n49_), .Y(men_men_n297_));
  OAI210     u0269(.A0(men_men_n270_), .A1(men_men_n293_), .B0(men_men_n297_), .Y(men_men_n298_));
  NAi21      u0270(.An(l), .B(k), .Y(men_men_n299_));
  NO2        u0271(.A(men_men_n299_), .B(men_men_n49_), .Y(men_men_n300_));
  NOi21      u0272(.An(l), .B(j), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n169_), .B(men_men_n301_), .Y(men_men_n302_));
  NA3        u0274(.A(men_men_n121_), .B(men_men_n120_), .C(g), .Y(men_men_n303_));
  OR3        u0275(.A(men_men_n72_), .B(men_men_n74_), .C(e), .Y(men_men_n304_));
  AOI210     u0276(.A0(men_men_n303_), .A1(men_men_n302_), .B0(men_men_n304_), .Y(men_men_n305_));
  INV        u0277(.A(men_men_n305_), .Y(men_men_n306_));
  NAi32      u0278(.An(j), .Bn(h), .C(i), .Y(men_men_n307_));
  NAi21      u0279(.An(m), .B(l), .Y(men_men_n308_));
  NO3        u0280(.A(men_men_n308_), .B(men_men_n307_), .C(men_men_n85_), .Y(men_men_n309_));
  NA2        u0281(.A(h), .B(g), .Y(men_men_n310_));
  NA2        u0282(.A(men_men_n175_), .B(men_men_n45_), .Y(men_men_n311_));
  NO2        u0283(.A(men_men_n311_), .B(men_men_n310_), .Y(men_men_n312_));
  OAI210     u0284(.A0(men_men_n312_), .A1(men_men_n309_), .B0(men_men_n170_), .Y(men_men_n313_));
  NA4        u0285(.A(men_men_n313_), .B(men_men_n306_), .C(men_men_n298_), .D(men_men_n291_), .Y(men_men_n314_));
  NO2        u0286(.A(men_men_n150_), .B(d), .Y(men_men_n315_));
  NA2        u0287(.A(men_men_n315_), .B(men_men_n53_), .Y(men_men_n316_));
  NO2        u0288(.A(men_men_n108_), .B(men_men_n105_), .Y(men_men_n317_));
  NAi32      u0289(.An(n), .Bn(m), .C(l), .Y(men_men_n318_));
  NO2        u0290(.A(men_men_n318_), .B(men_men_n307_), .Y(men_men_n319_));
  AOI220     u0291(.A0(men_men_n319_), .A1(men_men_n190_), .B0(men_men_n317_), .B1(men_men_n59_), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n125_), .B(men_men_n119_), .Y(men_men_n321_));
  NAi31      u0293(.An(k), .B(l), .C(j), .Y(men_men_n322_));
  OAI210     u0294(.A0(men_men_n299_), .A1(j), .B0(men_men_n322_), .Y(men_men_n323_));
  NOi21      u0295(.An(men_men_n323_), .B(men_men_n123_), .Y(men_men_n324_));
  NA2        u0296(.A(men_men_n324_), .B(men_men_n321_), .Y(men_men_n325_));
  NA3        u0297(.A(men_men_n325_), .B(men_men_n320_), .C(men_men_n316_), .Y(men_men_n326_));
  NO4        u0298(.A(men_men_n326_), .B(men_men_n314_), .C(men_men_n287_), .D(men_men_n277_), .Y(men_men_n327_));
  NA2        u0299(.A(men_men_n261_), .B(men_men_n199_), .Y(men_men_n328_));
  NAi21      u0300(.An(m), .B(k), .Y(men_men_n329_));
  NO2        u0301(.A(men_men_n232_), .B(men_men_n329_), .Y(men_men_n330_));
  NAi41      u0302(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n331_));
  NO2        u0303(.A(men_men_n331_), .B(men_men_n156_), .Y(men_men_n332_));
  NA2        u0304(.A(men_men_n332_), .B(men_men_n330_), .Y(men_men_n333_));
  NAi31      u0305(.An(i), .B(l), .C(h), .Y(men_men_n334_));
  NO4        u0306(.A(men_men_n334_), .B(men_men_n156_), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n335_));
  NA2        u0307(.A(e), .B(c), .Y(men_men_n336_));
  NO3        u0308(.A(men_men_n336_), .B(n), .C(d), .Y(men_men_n337_));
  NOi21      u0309(.An(f), .B(h), .Y(men_men_n338_));
  NA2        u0310(.A(men_men_n338_), .B(men_men_n121_), .Y(men_men_n339_));
  NO2        u0311(.A(men_men_n339_), .B(men_men_n221_), .Y(men_men_n340_));
  NAi31      u0312(.An(d), .B(e), .C(b), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n136_), .B(men_men_n341_), .Y(men_men_n342_));
  NA2        u0314(.A(men_men_n342_), .B(men_men_n340_), .Y(men_men_n343_));
  NAi41      u0315(.An(men_men_n335_), .B(men_men_n343_), .C(men_men_n333_), .D(men_men_n328_), .Y(men_men_n344_));
  NO4        u0316(.A(men_men_n331_), .B(men_men_n80_), .C(men_men_n71_), .D(men_men_n221_), .Y(men_men_n345_));
  NA2        u0317(.A(men_men_n256_), .B(men_men_n106_), .Y(men_men_n346_));
  OR2        u0318(.A(men_men_n346_), .B(men_men_n210_), .Y(men_men_n347_));
  NOi31      u0319(.An(l), .B(n), .C(m), .Y(men_men_n348_));
  NA2        u0320(.A(men_men_n348_), .B(men_men_n222_), .Y(men_men_n349_));
  NO2        u0321(.A(men_men_n349_), .B(men_men_n200_), .Y(men_men_n350_));
  NAi32      u0322(.An(men_men_n350_), .Bn(men_men_n345_), .C(men_men_n347_), .Y(men_men_n351_));
  NAi32      u0323(.An(m), .Bn(j), .C(k), .Y(men_men_n352_));
  NAi41      u0324(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n353_));
  OAI210     u0325(.A0(men_men_n218_), .A1(men_men_n352_), .B0(men_men_n353_), .Y(men_men_n354_));
  NOi31      u0326(.An(j), .B(m), .C(k), .Y(men_men_n355_));
  NO2        u0327(.A(men_men_n129_), .B(men_men_n355_), .Y(men_men_n356_));
  AN3        u0328(.A(h), .B(g), .C(f), .Y(men_men_n357_));
  NAi31      u0329(.An(men_men_n356_), .B(men_men_n357_), .C(men_men_n354_), .Y(men_men_n358_));
  NOi32      u0330(.An(m), .Bn(j), .C(l), .Y(men_men_n359_));
  NO2        u0331(.A(men_men_n359_), .B(men_men_n99_), .Y(men_men_n360_));
  NAi32      u0332(.An(men_men_n360_), .Bn(men_men_n207_), .C(men_men_n315_), .Y(men_men_n361_));
  NO2        u0333(.A(men_men_n308_), .B(men_men_n307_), .Y(men_men_n362_));
  NO2        u0334(.A(men_men_n224_), .B(g), .Y(men_men_n363_));
  NO2        u0335(.A(men_men_n162_), .B(men_men_n85_), .Y(men_men_n364_));
  AOI220     u0336(.A0(men_men_n364_), .A1(men_men_n363_), .B0(men_men_n253_), .B1(men_men_n362_), .Y(men_men_n365_));
  NA2        u0337(.A(men_men_n239_), .B(men_men_n80_), .Y(men_men_n366_));
  NA3        u0338(.A(men_men_n366_), .B(men_men_n357_), .C(men_men_n219_), .Y(men_men_n367_));
  NA4        u0339(.A(men_men_n367_), .B(men_men_n365_), .C(men_men_n361_), .D(men_men_n358_), .Y(men_men_n368_));
  NA3        u0340(.A(h), .B(g), .C(f), .Y(men_men_n369_));
  NO2        u0341(.A(men_men_n369_), .B(men_men_n76_), .Y(men_men_n370_));
  NA2        u0342(.A(men_men_n353_), .B(men_men_n218_), .Y(men_men_n371_));
  NA2        u0343(.A(men_men_n169_), .B(e), .Y(men_men_n372_));
  NO2        u0344(.A(men_men_n372_), .B(men_men_n41_), .Y(men_men_n373_));
  AOI220     u0345(.A0(men_men_n373_), .A1(men_men_n321_), .B0(men_men_n371_), .B1(men_men_n370_), .Y(men_men_n374_));
  NOi32      u0346(.An(j), .Bn(g), .C(i), .Y(men_men_n375_));
  NA3        u0347(.A(men_men_n375_), .B(men_men_n299_), .C(men_men_n116_), .Y(men_men_n376_));
  AO210      u0348(.A0(men_men_n114_), .A1(men_men_n32_), .B0(men_men_n376_), .Y(men_men_n377_));
  NOi32      u0349(.An(e), .Bn(b), .C(a), .Y(men_men_n378_));
  AN2        u0350(.A(l), .B(j), .Y(men_men_n379_));
  NO2        u0351(.A(men_men_n329_), .B(men_men_n379_), .Y(men_men_n380_));
  NO3        u0352(.A(men_men_n331_), .B(men_men_n71_), .C(men_men_n221_), .Y(men_men_n381_));
  NA3        u0353(.A(men_men_n215_), .B(men_men_n213_), .C(men_men_n35_), .Y(men_men_n382_));
  AOI220     u0354(.A0(men_men_n382_), .A1(men_men_n378_), .B0(men_men_n381_), .B1(men_men_n380_), .Y(men_men_n383_));
  NO2        u0355(.A(men_men_n341_), .B(n), .Y(men_men_n384_));
  NA2        u0356(.A(men_men_n214_), .B(k), .Y(men_men_n385_));
  NA3        u0357(.A(m), .B(men_men_n115_), .C(men_men_n220_), .Y(men_men_n386_));
  NA4        u0358(.A(men_men_n209_), .B(men_men_n88_), .C(g), .D(men_men_n220_), .Y(men_men_n387_));
  OAI210     u0359(.A0(men_men_n386_), .A1(men_men_n385_), .B0(men_men_n387_), .Y(men_men_n388_));
  NAi41      u0360(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n389_));
  NA2        u0361(.A(men_men_n51_), .B(men_men_n116_), .Y(men_men_n390_));
  NO2        u0362(.A(men_men_n390_), .B(men_men_n389_), .Y(men_men_n391_));
  AOI220     u0363(.A0(men_men_n391_), .A1(b), .B0(men_men_n388_), .B1(men_men_n384_), .Y(men_men_n392_));
  NA4        u0364(.A(men_men_n392_), .B(men_men_n383_), .C(men_men_n377_), .D(men_men_n374_), .Y(men_men_n393_));
  NO4        u0365(.A(men_men_n393_), .B(men_men_n368_), .C(men_men_n351_), .D(men_men_n344_), .Y(men_men_n394_));
  NA4        u0366(.A(men_men_n394_), .B(men_men_n327_), .C(men_men_n275_), .D(men_men_n205_), .Y(men10));
  NA3        u0367(.A(m), .B(k), .C(i), .Y(men_men_n396_));
  NO3        u0368(.A(men_men_n396_), .B(j), .C(men_men_n221_), .Y(men_men_n397_));
  NOi21      u0369(.An(e), .B(f), .Y(men_men_n398_));
  NO4        u0370(.A(men_men_n157_), .B(men_men_n398_), .C(n), .D(men_men_n113_), .Y(men_men_n399_));
  NAi31      u0371(.An(b), .B(f), .C(c), .Y(men_men_n400_));
  INV        u0372(.A(men_men_n400_), .Y(men_men_n401_));
  NOi32      u0373(.An(k), .Bn(h), .C(j), .Y(men_men_n402_));
  NA2        u0374(.A(men_men_n402_), .B(men_men_n228_), .Y(men_men_n403_));
  INV        u0375(.A(men_men_n403_), .Y(men_men_n404_));
  AOI220     u0376(.A0(men_men_n404_), .A1(men_men_n401_), .B0(men_men_n399_), .B1(men_men_n397_), .Y(men_men_n405_));
  AN2        u0377(.A(j), .B(h), .Y(men_men_n406_));
  NO3        u0378(.A(n), .B(m), .C(k), .Y(men_men_n407_));
  NA2        u0379(.A(men_men_n407_), .B(men_men_n406_), .Y(men_men_n408_));
  NO3        u0380(.A(men_men_n408_), .B(men_men_n157_), .C(men_men_n220_), .Y(men_men_n409_));
  OR2        u0381(.A(m), .B(k), .Y(men_men_n410_));
  NO2        u0382(.A(men_men_n181_), .B(men_men_n410_), .Y(men_men_n411_));
  NA4        u0383(.A(n), .B(f), .C(c), .D(men_men_n119_), .Y(men_men_n412_));
  NOi32      u0384(.An(d), .Bn(a), .C(c), .Y(men_men_n413_));
  NA2        u0385(.A(men_men_n413_), .B(men_men_n188_), .Y(men_men_n414_));
  NAi21      u0386(.An(i), .B(g), .Y(men_men_n415_));
  NAi31      u0387(.An(k), .B(m), .C(j), .Y(men_men_n416_));
  NO3        u0388(.A(men_men_n416_), .B(men_men_n415_), .C(n), .Y(men_men_n417_));
  NOi21      u0389(.An(men_men_n417_), .B(men_men_n414_), .Y(men_men_n418_));
  NO2        u0390(.A(men_men_n418_), .B(men_men_n409_), .Y(men_men_n419_));
  NO2        u0391(.A(men_men_n412_), .B(men_men_n308_), .Y(men_men_n420_));
  NOi32      u0392(.An(f), .Bn(d), .C(c), .Y(men_men_n421_));
  AOI220     u0393(.A0(men_men_n421_), .A1(men_men_n319_), .B0(men_men_n420_), .B1(men_men_n222_), .Y(men_men_n422_));
  NA3        u0394(.A(men_men_n422_), .B(men_men_n419_), .C(men_men_n405_), .Y(men_men_n423_));
  NO2        u0395(.A(men_men_n59_), .B(men_men_n119_), .Y(men_men_n424_));
  NA2        u0396(.A(men_men_n256_), .B(men_men_n424_), .Y(men_men_n425_));
  INV        u0397(.A(e), .Y(men_men_n426_));
  NA2        u0398(.A(men_men_n46_), .B(e), .Y(men_men_n427_));
  OAI220     u0399(.A0(men_men_n427_), .A1(men_men_n206_), .B0(men_men_n210_), .B1(men_men_n426_), .Y(men_men_n428_));
  AN2        u0400(.A(g), .B(e), .Y(men_men_n429_));
  NA3        u0401(.A(men_men_n429_), .B(men_men_n209_), .C(i), .Y(men_men_n430_));
  OAI210     u0402(.A0(men_men_n90_), .A1(men_men_n426_), .B0(men_men_n430_), .Y(men_men_n431_));
  NO2        u0403(.A(men_men_n102_), .B(men_men_n426_), .Y(men_men_n432_));
  NO3        u0404(.A(men_men_n432_), .B(men_men_n431_), .C(men_men_n428_), .Y(men_men_n433_));
  NOi32      u0405(.An(h), .Bn(e), .C(g), .Y(men_men_n434_));
  NA3        u0406(.A(men_men_n434_), .B(men_men_n301_), .C(m), .Y(men_men_n435_));
  NOi21      u0407(.An(g), .B(h), .Y(men_men_n436_));
  AN3        u0408(.A(m), .B(l), .C(i), .Y(men_men_n437_));
  NA3        u0409(.A(men_men_n437_), .B(men_men_n436_), .C(e), .Y(men_men_n438_));
  AN3        u0410(.A(h), .B(g), .C(e), .Y(men_men_n439_));
  NA2        u0411(.A(men_men_n439_), .B(men_men_n99_), .Y(men_men_n440_));
  AN3        u0412(.A(men_men_n440_), .B(men_men_n438_), .C(men_men_n435_), .Y(men_men_n441_));
  AOI210     u0413(.A0(men_men_n441_), .A1(men_men_n433_), .B0(men_men_n425_), .Y(men_men_n442_));
  NA3        u0414(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n443_));
  NO2        u0415(.A(men_men_n443_), .B(men_men_n425_), .Y(men_men_n444_));
  NA3        u0416(.A(men_men_n413_), .B(men_men_n188_), .C(men_men_n85_), .Y(men_men_n445_));
  NAi31      u0417(.An(b), .B(c), .C(a), .Y(men_men_n446_));
  NO2        u0418(.A(men_men_n446_), .B(n), .Y(men_men_n447_));
  OAI210     u0419(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n448_));
  NO2        u0420(.A(men_men_n448_), .B(men_men_n153_), .Y(men_men_n449_));
  NA2        u0421(.A(men_men_n449_), .B(men_men_n447_), .Y(men_men_n450_));
  INV        u0422(.A(men_men_n450_), .Y(men_men_n451_));
  NO4        u0423(.A(men_men_n451_), .B(men_men_n444_), .C(men_men_n442_), .D(men_men_n423_), .Y(men_men_n452_));
  NA2        u0424(.A(i), .B(g), .Y(men_men_n453_));
  NO3        u0425(.A(men_men_n285_), .B(men_men_n453_), .C(c), .Y(men_men_n454_));
  NOi21      u0426(.An(a), .B(n), .Y(men_men_n455_));
  NOi21      u0427(.An(d), .B(c), .Y(men_men_n456_));
  NA2        u0428(.A(men_men_n456_), .B(men_men_n455_), .Y(men_men_n457_));
  NA3        u0429(.A(i), .B(g), .C(f), .Y(men_men_n458_));
  OR2        u0430(.A(men_men_n458_), .B(men_men_n70_), .Y(men_men_n459_));
  NA3        u0431(.A(men_men_n437_), .B(men_men_n436_), .C(men_men_n188_), .Y(men_men_n460_));
  AOI210     u0432(.A0(men_men_n460_), .A1(men_men_n459_), .B0(men_men_n457_), .Y(men_men_n461_));
  AOI210     u0433(.A0(men_men_n454_), .A1(men_men_n300_), .B0(men_men_n461_), .Y(men_men_n462_));
  OR2        u0434(.A(n), .B(m), .Y(men_men_n463_));
  NO2        u0435(.A(men_men_n463_), .B(men_men_n158_), .Y(men_men_n464_));
  NO2        u0436(.A(men_men_n189_), .B(men_men_n153_), .Y(men_men_n465_));
  NA2        u0437(.A(men_men_n464_), .B(men_men_n465_), .Y(men_men_n466_));
  INV        u0438(.A(men_men_n390_), .Y(men_men_n467_));
  NA3        u0439(.A(men_men_n467_), .B(men_men_n378_), .C(d), .Y(men_men_n468_));
  NO2        u0440(.A(men_men_n446_), .B(men_men_n49_), .Y(men_men_n469_));
  NO3        u0441(.A(men_men_n65_), .B(men_men_n115_), .C(e), .Y(men_men_n470_));
  NAi21      u0442(.An(k), .B(j), .Y(men_men_n471_));
  NA2        u0443(.A(men_men_n259_), .B(men_men_n471_), .Y(men_men_n472_));
  NA3        u0444(.A(men_men_n472_), .B(men_men_n470_), .C(men_men_n469_), .Y(men_men_n473_));
  NAi21      u0445(.An(e), .B(d), .Y(men_men_n474_));
  NO2        u0446(.A(men_men_n474_), .B(men_men_n56_), .Y(men_men_n475_));
  NO2        u0447(.A(men_men_n260_), .B(men_men_n220_), .Y(men_men_n476_));
  NA3        u0448(.A(men_men_n476_), .B(men_men_n475_), .C(men_men_n233_), .Y(men_men_n477_));
  NA4        u0449(.A(men_men_n477_), .B(men_men_n473_), .C(men_men_n468_), .D(men_men_n466_), .Y(men_men_n478_));
  NO2        u0450(.A(men_men_n349_), .B(men_men_n220_), .Y(men_men_n479_));
  NA2        u0451(.A(men_men_n479_), .B(men_men_n475_), .Y(men_men_n480_));
  NOi31      u0452(.An(n), .B(m), .C(k), .Y(men_men_n481_));
  AOI220     u0453(.A0(men_men_n481_), .A1(men_men_n406_), .B0(men_men_n228_), .B1(men_men_n50_), .Y(men_men_n482_));
  NAi31      u0454(.An(g), .B(f), .C(c), .Y(men_men_n483_));
  OR3        u0455(.A(men_men_n483_), .B(men_men_n482_), .C(e), .Y(men_men_n484_));
  NA3        u0456(.A(men_men_n484_), .B(men_men_n480_), .C(men_men_n320_), .Y(men_men_n485_));
  NOi41      u0457(.An(men_men_n462_), .B(men_men_n485_), .C(men_men_n478_), .D(men_men_n273_), .Y(men_men_n486_));
  NOi32      u0458(.An(c), .Bn(a), .C(b), .Y(men_men_n487_));
  NA2        u0459(.A(men_men_n487_), .B(men_men_n116_), .Y(men_men_n488_));
  NA2        u0460(.A(men_men_n283_), .B(men_men_n158_), .Y(men_men_n489_));
  AN2        u0461(.A(e), .B(d), .Y(men_men_n490_));
  NA2        u0462(.A(men_men_n490_), .B(men_men_n489_), .Y(men_men_n491_));
  INV        u0463(.A(men_men_n153_), .Y(men_men_n492_));
  NO2        u0464(.A(men_men_n135_), .B(men_men_n41_), .Y(men_men_n493_));
  NO2        u0465(.A(men_men_n65_), .B(e), .Y(men_men_n494_));
  NOi31      u0466(.An(j), .B(k), .C(i), .Y(men_men_n495_));
  NOi21      u0467(.An(men_men_n172_), .B(men_men_n495_), .Y(men_men_n496_));
  NA4        u0468(.A(men_men_n334_), .B(men_men_n496_), .C(men_men_n267_), .D(men_men_n122_), .Y(men_men_n497_));
  AOI220     u0469(.A0(men_men_n497_), .A1(men_men_n494_), .B0(men_men_n493_), .B1(men_men_n492_), .Y(men_men_n498_));
  AOI210     u0470(.A0(men_men_n498_), .A1(men_men_n491_), .B0(men_men_n488_), .Y(men_men_n499_));
  NO2        u0471(.A(men_men_n216_), .B(men_men_n211_), .Y(men_men_n500_));
  NOi21      u0472(.An(a), .B(b), .Y(men_men_n501_));
  NA3        u0473(.A(e), .B(d), .C(c), .Y(men_men_n502_));
  NAi21      u0474(.An(men_men_n502_), .B(men_men_n501_), .Y(men_men_n503_));
  NO2        u0475(.A(men_men_n445_), .B(men_men_n210_), .Y(men_men_n504_));
  NOi21      u0476(.An(men_men_n503_), .B(men_men_n504_), .Y(men_men_n505_));
  AOI210     u0477(.A0(men_men_n276_), .A1(men_men_n500_), .B0(men_men_n505_), .Y(men_men_n506_));
  NA2        u0478(.A(men_men_n401_), .B(men_men_n159_), .Y(men_men_n507_));
  OR2        u0479(.A(k), .B(j), .Y(men_men_n508_));
  NA2        u0480(.A(l), .B(k), .Y(men_men_n509_));
  NA3        u0481(.A(men_men_n509_), .B(men_men_n508_), .C(men_men_n228_), .Y(men_men_n510_));
  AOI210     u0482(.A0(men_men_n239_), .A1(men_men_n352_), .B0(men_men_n85_), .Y(men_men_n511_));
  NOi21      u0483(.An(men_men_n510_), .B(men_men_n511_), .Y(men_men_n512_));
  NA3        u0484(.A(men_men_n288_), .B(men_men_n132_), .C(men_men_n130_), .Y(men_men_n513_));
  NA2        u0485(.A(men_men_n413_), .B(men_men_n116_), .Y(men_men_n514_));
  NO4        u0486(.A(men_men_n514_), .B(men_men_n96_), .C(men_men_n115_), .D(e), .Y(men_men_n515_));
  NO3        u0487(.A(men_men_n445_), .B(men_men_n93_), .C(men_men_n135_), .Y(men_men_n516_));
  NO4        u0488(.A(men_men_n516_), .B(men_men_n515_), .C(men_men_n513_), .D(men_men_n335_), .Y(men_men_n517_));
  NA2        u0489(.A(men_men_n517_), .B(men_men_n507_), .Y(men_men_n518_));
  NO3        u0490(.A(men_men_n518_), .B(men_men_n506_), .C(men_men_n499_), .Y(men_men_n519_));
  NA2        u0491(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n520_));
  NO2        u0492(.A(men_men_n194_), .B(men_men_n56_), .Y(men_men_n521_));
  NAi31      u0493(.An(j), .B(l), .C(i), .Y(men_men_n522_));
  OAI210     u0494(.A0(men_men_n522_), .A1(men_men_n136_), .B0(men_men_n105_), .Y(men_men_n523_));
  NA4        u0495(.A(men_men_n523_), .B(men_men_n521_), .C(d), .D(b), .Y(men_men_n524_));
  NO3        u0496(.A(men_men_n414_), .B(men_men_n360_), .C(men_men_n207_), .Y(men_men_n525_));
  NO2        u0497(.A(men_men_n414_), .B(men_men_n390_), .Y(men_men_n526_));
  NO4        u0498(.A(men_men_n526_), .B(men_men_n525_), .C(men_men_n191_), .D(men_men_n317_), .Y(men_men_n527_));
  NA4        u0499(.A(men_men_n527_), .B(men_men_n524_), .C(men_men_n520_), .D(men_men_n248_), .Y(men_men_n528_));
  OAI210     u0500(.A0(men_men_n131_), .A1(men_men_n129_), .B0(n), .Y(men_men_n529_));
  NO2        u0501(.A(men_men_n529_), .B(men_men_n135_), .Y(men_men_n530_));
  AO210      u0502(.A0(men_men_n309_), .A1(men_men_n221_), .B0(men_men_n250_), .Y(men_men_n531_));
  OA210      u0503(.A0(men_men_n531_), .A1(men_men_n530_), .B0(men_men_n199_), .Y(men_men_n532_));
  XO2        u0504(.A(i), .B(h), .Y(men_men_n533_));
  NAi31      u0505(.An(men_men_n309_), .B(men_men_n482_), .C(men_men_n403_), .Y(men_men_n534_));
  NOi32      u0506(.An(men_men_n534_), .Bn(men_men_n494_), .C(men_men_n278_), .Y(men_men_n535_));
  NAi31      u0507(.An(c), .B(f), .C(d), .Y(men_men_n536_));
  AOI210     u0508(.A0(men_men_n289_), .A1(men_men_n202_), .B0(men_men_n536_), .Y(men_men_n537_));
  NOi21      u0509(.An(men_men_n83_), .B(men_men_n537_), .Y(men_men_n538_));
  NA3        u0510(.A(men_men_n399_), .B(men_men_n99_), .C(men_men_n98_), .Y(men_men_n539_));
  NA2        u0511(.A(men_men_n234_), .B(men_men_n111_), .Y(men_men_n540_));
  AOI210     u0512(.A0(men_men_n540_), .A1(men_men_n187_), .B0(men_men_n536_), .Y(men_men_n541_));
  AOI210     u0513(.A0(men_men_n376_), .A1(men_men_n35_), .B0(men_men_n503_), .Y(men_men_n542_));
  NOi31      u0514(.An(men_men_n539_), .B(men_men_n542_), .C(men_men_n541_), .Y(men_men_n543_));
  AO220      u0515(.A0(men_men_n297_), .A1(men_men_n270_), .B0(men_men_n173_), .B1(men_men_n66_), .Y(men_men_n544_));
  NA3        u0516(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n545_));
  NO2        u0517(.A(men_men_n545_), .B(men_men_n457_), .Y(men_men_n546_));
  NO2        u0518(.A(men_men_n546_), .B(men_men_n305_), .Y(men_men_n547_));
  NAi41      u0519(.An(men_men_n544_), .B(men_men_n547_), .C(men_men_n543_), .D(men_men_n538_), .Y(men_men_n548_));
  NO4        u0520(.A(men_men_n548_), .B(men_men_n535_), .C(men_men_n532_), .D(men_men_n528_), .Y(men_men_n549_));
  NA4        u0521(.A(men_men_n549_), .B(men_men_n519_), .C(men_men_n486_), .D(men_men_n452_), .Y(men11));
  NO2        u0522(.A(men_men_n72_), .B(f), .Y(men_men_n551_));
  NA2        u0523(.A(j), .B(g), .Y(men_men_n552_));
  NAi31      u0524(.An(i), .B(m), .C(l), .Y(men_men_n553_));
  NA3        u0525(.A(m), .B(k), .C(j), .Y(men_men_n554_));
  OAI220     u0526(.A0(men_men_n554_), .A1(men_men_n135_), .B0(men_men_n553_), .B1(men_men_n552_), .Y(men_men_n555_));
  NA2        u0527(.A(men_men_n555_), .B(men_men_n551_), .Y(men_men_n556_));
  NOi32      u0528(.An(e), .Bn(b), .C(f), .Y(men_men_n557_));
  NA2        u0529(.A(men_men_n266_), .B(men_men_n116_), .Y(men_men_n558_));
  NA2        u0530(.A(men_men_n46_), .B(j), .Y(men_men_n559_));
  OAI220     u0531(.A0(men_men_n559_), .A1(men_men_n311_), .B0(men_men_n558_), .B1(men_men_n221_), .Y(men_men_n560_));
  NAi31      u0532(.An(d), .B(e), .C(a), .Y(men_men_n561_));
  NO2        u0533(.A(men_men_n561_), .B(n), .Y(men_men_n562_));
  AOI220     u0534(.A0(men_men_n562_), .A1(men_men_n103_), .B0(men_men_n560_), .B1(men_men_n557_), .Y(men_men_n563_));
  NAi41      u0535(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n564_));
  AN2        u0536(.A(men_men_n564_), .B(men_men_n389_), .Y(men_men_n565_));
  NA2        u0537(.A(j), .B(i), .Y(men_men_n566_));
  NAi31      u0538(.An(n), .B(m), .C(k), .Y(men_men_n567_));
  NO3        u0539(.A(men_men_n567_), .B(men_men_n566_), .C(men_men_n115_), .Y(men_men_n568_));
  NO4        u0540(.A(n), .B(d), .C(men_men_n119_), .D(a), .Y(men_men_n569_));
  OR2        u0541(.A(n), .B(c), .Y(men_men_n570_));
  NO2        u0542(.A(men_men_n570_), .B(men_men_n155_), .Y(men_men_n571_));
  NO2        u0543(.A(men_men_n571_), .B(men_men_n569_), .Y(men_men_n572_));
  NOi32      u0544(.An(g), .Bn(f), .C(i), .Y(men_men_n573_));
  AOI220     u0545(.A0(men_men_n573_), .A1(men_men_n101_), .B0(men_men_n555_), .B1(f), .Y(men_men_n574_));
  NO2        u0546(.A(men_men_n283_), .B(men_men_n49_), .Y(men_men_n575_));
  NO2        u0547(.A(men_men_n574_), .B(men_men_n572_), .Y(men_men_n576_));
  INV        u0548(.A(men_men_n576_), .Y(men_men_n577_));
  NA2        u0549(.A(men_men_n145_), .B(men_men_n34_), .Y(men_men_n578_));
  OAI220     u0550(.A0(men_men_n578_), .A1(m), .B0(men_men_n559_), .B1(men_men_n239_), .Y(men_men_n579_));
  NOi41      u0551(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n580_));
  NAi32      u0552(.An(e), .Bn(b), .C(c), .Y(men_men_n581_));
  AN2        u0553(.A(men_men_n353_), .B(men_men_n331_), .Y(men_men_n582_));
  NA2        u0554(.A(men_men_n582_), .B(men_men_n581_), .Y(men_men_n583_));
  OA210      u0555(.A0(men_men_n583_), .A1(men_men_n580_), .B0(men_men_n579_), .Y(men_men_n584_));
  OAI220     u0556(.A0(men_men_n416_), .A1(men_men_n415_), .B0(men_men_n553_), .B1(men_men_n552_), .Y(men_men_n585_));
  NAi31      u0557(.An(d), .B(c), .C(a), .Y(men_men_n586_));
  NO2        u0558(.A(men_men_n586_), .B(n), .Y(men_men_n587_));
  NA3        u0559(.A(men_men_n587_), .B(men_men_n585_), .C(e), .Y(men_men_n588_));
  NO3        u0560(.A(men_men_n61_), .B(men_men_n49_), .C(men_men_n221_), .Y(men_men_n589_));
  NO2        u0561(.A(men_men_n237_), .B(men_men_n113_), .Y(men_men_n590_));
  OAI210     u0562(.A0(men_men_n589_), .A1(men_men_n417_), .B0(men_men_n590_), .Y(men_men_n591_));
  NA2        u0563(.A(men_men_n591_), .B(men_men_n588_), .Y(men_men_n592_));
  NO2        u0564(.A(men_men_n285_), .B(n), .Y(men_men_n593_));
  NO2        u0565(.A(men_men_n447_), .B(men_men_n593_), .Y(men_men_n594_));
  NA2        u0566(.A(men_men_n585_), .B(f), .Y(men_men_n595_));
  NAi32      u0567(.An(d), .Bn(a), .C(b), .Y(men_men_n596_));
  NO2        u0568(.A(men_men_n596_), .B(men_men_n49_), .Y(men_men_n597_));
  NA2        u0569(.A(h), .B(f), .Y(men_men_n598_));
  NO2        u0570(.A(men_men_n598_), .B(men_men_n96_), .Y(men_men_n599_));
  NO3        u0571(.A(men_men_n183_), .B(men_men_n181_), .C(g), .Y(men_men_n600_));
  AOI220     u0572(.A0(men_men_n600_), .A1(men_men_n58_), .B0(men_men_n599_), .B1(men_men_n597_), .Y(men_men_n601_));
  OAI210     u0573(.A0(men_men_n595_), .A1(men_men_n594_), .B0(men_men_n601_), .Y(men_men_n602_));
  AN3        u0574(.A(j), .B(h), .C(g), .Y(men_men_n603_));
  NO2        u0575(.A(men_men_n152_), .B(c), .Y(men_men_n604_));
  NA3        u0576(.A(men_men_n604_), .B(men_men_n603_), .C(men_men_n481_), .Y(men_men_n605_));
  NA3        u0577(.A(f), .B(d), .C(b), .Y(men_men_n606_));
  NO4        u0578(.A(men_men_n606_), .B(men_men_n183_), .C(men_men_n181_), .D(g), .Y(men_men_n607_));
  NAi21      u0579(.An(men_men_n607_), .B(men_men_n605_), .Y(men_men_n608_));
  NO4        u0580(.A(men_men_n608_), .B(men_men_n602_), .C(men_men_n592_), .D(men_men_n584_), .Y(men_men_n609_));
  AN4        u0581(.A(men_men_n609_), .B(men_men_n577_), .C(men_men_n563_), .D(men_men_n556_), .Y(men_men_n610_));
  INV        u0582(.A(k), .Y(men_men_n611_));
  NA3        u0583(.A(l), .B(men_men_n611_), .C(i), .Y(men_men_n612_));
  INV        u0584(.A(men_men_n612_), .Y(men_men_n613_));
  NA4        u0585(.A(men_men_n413_), .B(men_men_n436_), .C(men_men_n188_), .D(men_men_n116_), .Y(men_men_n614_));
  NAi32      u0586(.An(h), .Bn(f), .C(g), .Y(men_men_n615_));
  NAi41      u0587(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n616_));
  OAI210     u0588(.A0(men_men_n561_), .A1(n), .B0(men_men_n616_), .Y(men_men_n617_));
  NA2        u0589(.A(men_men_n617_), .B(m), .Y(men_men_n618_));
  NAi31      u0590(.An(h), .B(g), .C(f), .Y(men_men_n619_));
  OR3        u0591(.A(men_men_n619_), .B(men_men_n285_), .C(men_men_n49_), .Y(men_men_n620_));
  NA4        u0592(.A(men_men_n436_), .B(men_men_n124_), .C(men_men_n116_), .D(e), .Y(men_men_n621_));
  AN2        u0593(.A(men_men_n621_), .B(men_men_n620_), .Y(men_men_n622_));
  OA210      u0594(.A0(men_men_n618_), .A1(men_men_n615_), .B0(men_men_n622_), .Y(men_men_n623_));
  NO3        u0595(.A(men_men_n615_), .B(men_men_n72_), .C(men_men_n74_), .Y(men_men_n624_));
  NO4        u0596(.A(men_men_n619_), .B(men_men_n570_), .C(men_men_n155_), .D(men_men_n74_), .Y(men_men_n625_));
  OR2        u0597(.A(men_men_n625_), .B(men_men_n624_), .Y(men_men_n626_));
  NAi31      u0598(.An(men_men_n626_), .B(men_men_n623_), .C(men_men_n614_), .Y(men_men_n627_));
  NAi31      u0599(.An(f), .B(h), .C(g), .Y(men_men_n628_));
  NO4        u0600(.A(men_men_n322_), .B(men_men_n628_), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n629_));
  NOi32      u0601(.An(b), .Bn(a), .C(c), .Y(men_men_n630_));
  NOi41      u0602(.An(men_men_n630_), .B(men_men_n369_), .C(men_men_n68_), .D(men_men_n120_), .Y(men_men_n631_));
  OR2        u0603(.A(men_men_n631_), .B(men_men_n629_), .Y(men_men_n632_));
  NOi32      u0604(.An(d), .Bn(a), .C(e), .Y(men_men_n633_));
  NA2        u0605(.A(men_men_n633_), .B(men_men_n116_), .Y(men_men_n634_));
  NO2        u0606(.A(n), .B(c), .Y(men_men_n635_));
  NA3        u0607(.A(men_men_n635_), .B(men_men_n29_), .C(m), .Y(men_men_n636_));
  NOi32      u0608(.An(e), .Bn(a), .C(d), .Y(men_men_n637_));
  AOI210     u0609(.A0(men_men_n29_), .A1(d), .B0(men_men_n637_), .Y(men_men_n638_));
  INV        u0610(.A(men_men_n578_), .Y(men_men_n639_));
  AOI210     u0611(.A0(men_men_n639_), .A1(men_men_n116_), .B0(men_men_n632_), .Y(men_men_n640_));
  OAI210     u0612(.A0(men_men_n255_), .A1(men_men_n88_), .B0(men_men_n640_), .Y(men_men_n641_));
  AOI210     u0613(.A0(men_men_n627_), .A1(men_men_n613_), .B0(men_men_n641_), .Y(men_men_n642_));
  NA2        u0614(.A(men_men_n483_), .B(men_men_n237_), .Y(men_men_n643_));
  NA2        u0615(.A(men_men_n75_), .B(men_men_n116_), .Y(men_men_n644_));
  NO2        u0616(.A(men_men_n644_), .B(men_men_n45_), .Y(men_men_n645_));
  NA3        u0617(.A(men_men_n580_), .B(men_men_n355_), .C(men_men_n46_), .Y(men_men_n646_));
  NOi32      u0618(.An(e), .Bn(c), .C(f), .Y(men_men_n647_));
  NOi21      u0619(.An(f), .B(g), .Y(men_men_n648_));
  NO2        u0620(.A(men_men_n648_), .B(men_men_n218_), .Y(men_men_n649_));
  NA2        u0621(.A(men_men_n649_), .B(men_men_n411_), .Y(men_men_n650_));
  NA3        u0622(.A(men_men_n650_), .B(men_men_n646_), .C(men_men_n185_), .Y(men_men_n651_));
  AOI210     u0623(.A0(men_men_n565_), .A1(men_men_n414_), .B0(men_men_n310_), .Y(men_men_n652_));
  NA2        u0624(.A(men_men_n652_), .B(men_men_n271_), .Y(men_men_n653_));
  NOi21      u0625(.An(j), .B(l), .Y(men_men_n654_));
  NAi21      u0626(.An(k), .B(h), .Y(men_men_n655_));
  NO2        u0627(.A(men_men_n655_), .B(men_men_n269_), .Y(men_men_n656_));
  NA2        u0628(.A(men_men_n656_), .B(men_men_n654_), .Y(men_men_n657_));
  OR2        u0629(.A(men_men_n657_), .B(men_men_n618_), .Y(men_men_n658_));
  NOi31      u0630(.An(m), .B(n), .C(k), .Y(men_men_n659_));
  NA2        u0631(.A(men_men_n654_), .B(men_men_n659_), .Y(men_men_n660_));
  AOI210     u0632(.A0(men_men_n414_), .A1(men_men_n389_), .B0(men_men_n310_), .Y(men_men_n661_));
  NAi21      u0633(.An(men_men_n660_), .B(men_men_n661_), .Y(men_men_n662_));
  NO2        u0634(.A(men_men_n285_), .B(men_men_n49_), .Y(men_men_n663_));
  NO2        u0635(.A(men_men_n322_), .B(men_men_n628_), .Y(men_men_n664_));
  NO2        u0636(.A(men_men_n561_), .B(men_men_n49_), .Y(men_men_n665_));
  AOI220     u0637(.A0(men_men_n665_), .A1(men_men_n664_), .B0(men_men_n663_), .B1(men_men_n599_), .Y(men_men_n666_));
  NA4        u0638(.A(men_men_n666_), .B(men_men_n662_), .C(men_men_n658_), .D(men_men_n653_), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n111_), .B(men_men_n36_), .Y(men_men_n668_));
  NO2        u0640(.A(k), .B(men_men_n221_), .Y(men_men_n669_));
  NO2        u0641(.A(men_men_n557_), .B(men_men_n378_), .Y(men_men_n670_));
  NO2        u0642(.A(men_men_n670_), .B(n), .Y(men_men_n671_));
  NAi31      u0643(.An(men_men_n668_), .B(men_men_n671_), .C(men_men_n669_), .Y(men_men_n672_));
  NO2        u0644(.A(men_men_n559_), .B(men_men_n183_), .Y(men_men_n673_));
  NA3        u0645(.A(men_men_n581_), .B(men_men_n278_), .C(men_men_n150_), .Y(men_men_n674_));
  NA2        u0646(.A(men_men_n674_), .B(men_men_n673_), .Y(men_men_n675_));
  AN3        u0647(.A(f), .B(d), .C(b), .Y(men_men_n676_));
  OAI210     u0648(.A0(men_men_n676_), .A1(men_men_n134_), .B0(n), .Y(men_men_n677_));
  NA3        u0649(.A(men_men_n533_), .B(men_men_n166_), .C(men_men_n221_), .Y(men_men_n678_));
  AOI210     u0650(.A0(men_men_n677_), .A1(men_men_n238_), .B0(men_men_n678_), .Y(men_men_n679_));
  NAi31      u0651(.An(m), .B(n), .C(k), .Y(men_men_n680_));
  OAI210     u0652(.A0(men_men_n139_), .A1(men_men_n680_), .B0(men_men_n257_), .Y(men_men_n681_));
  OAI210     u0653(.A0(men_men_n681_), .A1(men_men_n679_), .B0(j), .Y(men_men_n682_));
  NA3        u0654(.A(men_men_n682_), .B(men_men_n675_), .C(men_men_n672_), .Y(men_men_n683_));
  NO3        u0655(.A(men_men_n683_), .B(men_men_n667_), .C(men_men_n651_), .Y(men_men_n684_));
  NA2        u0656(.A(men_men_n399_), .B(men_men_n169_), .Y(men_men_n685_));
  NAi31      u0657(.An(g), .B(h), .C(f), .Y(men_men_n686_));
  OR3        u0658(.A(men_men_n686_), .B(men_men_n285_), .C(n), .Y(men_men_n687_));
  OA210      u0659(.A0(men_men_n561_), .A1(n), .B0(men_men_n616_), .Y(men_men_n688_));
  NA3        u0660(.A(men_men_n434_), .B(men_men_n124_), .C(men_men_n85_), .Y(men_men_n689_));
  OAI210     u0661(.A0(men_men_n688_), .A1(men_men_n92_), .B0(men_men_n689_), .Y(men_men_n690_));
  NOi21      u0662(.An(men_men_n687_), .B(men_men_n690_), .Y(men_men_n691_));
  AOI210     u0663(.A0(men_men_n691_), .A1(men_men_n685_), .B0(men_men_n554_), .Y(men_men_n692_));
  NO3        u0664(.A(g), .B(men_men_n220_), .C(men_men_n56_), .Y(men_men_n693_));
  NAi21      u0665(.An(h), .B(j), .Y(men_men_n694_));
  OAI220     u0666(.A0(men_men_n694_), .A1(men_men_n105_), .B0(men_men_n540_), .B1(men_men_n88_), .Y(men_men_n695_));
  OAI210     u0667(.A0(men_men_n695_), .A1(men_men_n411_), .B0(men_men_n693_), .Y(men_men_n696_));
  OR2        u0668(.A(men_men_n72_), .B(men_men_n74_), .Y(men_men_n697_));
  NA2        u0669(.A(men_men_n630_), .B(men_men_n357_), .Y(men_men_n698_));
  OA220      u0670(.A0(men_men_n660_), .A1(men_men_n698_), .B0(men_men_n657_), .B1(men_men_n697_), .Y(men_men_n699_));
  NA3        u0671(.A(men_men_n551_), .B(men_men_n101_), .C(men_men_n100_), .Y(men_men_n700_));
  AN2        u0672(.A(h), .B(f), .Y(men_men_n701_));
  NA2        u0673(.A(men_men_n701_), .B(men_men_n37_), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n101_), .B(men_men_n46_), .Y(men_men_n703_));
  OAI220     u0675(.A0(men_men_n703_), .A1(men_men_n346_), .B0(men_men_n702_), .B1(men_men_n488_), .Y(men_men_n704_));
  AOI210     u0676(.A0(men_men_n596_), .A1(men_men_n446_), .B0(men_men_n49_), .Y(men_men_n705_));
  OAI220     u0677(.A0(men_men_n619_), .A1(men_men_n612_), .B0(men_men_n339_), .B1(men_men_n552_), .Y(men_men_n706_));
  AOI210     u0678(.A0(men_men_n706_), .A1(men_men_n705_), .B0(men_men_n704_), .Y(men_men_n707_));
  NA4        u0679(.A(men_men_n707_), .B(men_men_n700_), .C(men_men_n699_), .D(men_men_n696_), .Y(men_men_n708_));
  NO2        u0680(.A(men_men_n259_), .B(f), .Y(men_men_n709_));
  NO2        u0681(.A(men_men_n648_), .B(men_men_n60_), .Y(men_men_n710_));
  NO3        u0682(.A(men_men_n710_), .B(men_men_n709_), .C(men_men_n34_), .Y(men_men_n711_));
  NA2        u0683(.A(men_men_n342_), .B(men_men_n145_), .Y(men_men_n712_));
  NA2        u0684(.A(men_men_n136_), .B(men_men_n49_), .Y(men_men_n713_));
  AOI220     u0685(.A0(men_men_n713_), .A1(men_men_n557_), .B0(men_men_n378_), .B1(men_men_n116_), .Y(men_men_n714_));
  OA220      u0686(.A0(men_men_n714_), .A1(men_men_n578_), .B0(men_men_n376_), .B1(men_men_n114_), .Y(men_men_n715_));
  OAI210     u0687(.A0(men_men_n712_), .A1(men_men_n711_), .B0(men_men_n715_), .Y(men_men_n716_));
  NO3        u0688(.A(men_men_n421_), .B(men_men_n199_), .C(men_men_n198_), .Y(men_men_n717_));
  NA2        u0689(.A(men_men_n717_), .B(men_men_n237_), .Y(men_men_n718_));
  NA3        u0690(.A(men_men_n718_), .B(men_men_n261_), .C(j), .Y(men_men_n719_));
  NO3        u0691(.A(men_men_n483_), .B(men_men_n181_), .C(i), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n487_), .B(men_men_n85_), .Y(men_men_n721_));
  NO4        u0693(.A(men_men_n554_), .B(men_men_n721_), .C(men_men_n135_), .D(men_men_n220_), .Y(men_men_n722_));
  INV        u0694(.A(men_men_n722_), .Y(men_men_n723_));
  NA4        u0695(.A(men_men_n723_), .B(men_men_n719_), .C(men_men_n539_), .D(men_men_n419_), .Y(men_men_n724_));
  NO4        u0696(.A(men_men_n724_), .B(men_men_n716_), .C(men_men_n708_), .D(men_men_n692_), .Y(men_men_n725_));
  NA4        u0697(.A(men_men_n725_), .B(men_men_n684_), .C(men_men_n642_), .D(men_men_n610_), .Y(men08));
  NO2        u0698(.A(k), .B(h), .Y(men_men_n727_));
  AO210      u0699(.A0(men_men_n259_), .A1(men_men_n471_), .B0(men_men_n727_), .Y(men_men_n728_));
  NO2        u0700(.A(men_men_n728_), .B(men_men_n308_), .Y(men_men_n729_));
  NA2        u0701(.A(men_men_n647_), .B(men_men_n85_), .Y(men_men_n730_));
  INV        u0702(.A(men_men_n516_), .Y(men_men_n731_));
  NA2        u0703(.A(men_men_n85_), .B(men_men_n113_), .Y(men_men_n732_));
  NO2        u0704(.A(men_men_n732_), .B(men_men_n57_), .Y(men_men_n733_));
  NO4        u0705(.A(men_men_n396_), .B(men_men_n115_), .C(j), .D(men_men_n221_), .Y(men_men_n734_));
  OAI210     u0706(.A0(men_men_n606_), .A1(men_men_n85_), .B0(men_men_n238_), .Y(men_men_n735_));
  AOI220     u0707(.A0(men_men_n735_), .A1(men_men_n363_), .B0(men_men_n734_), .B1(men_men_n733_), .Y(men_men_n736_));
  AOI210     u0708(.A0(men_men_n606_), .A1(men_men_n162_), .B0(men_men_n85_), .Y(men_men_n737_));
  NA4        u0709(.A(men_men_n223_), .B(men_men_n145_), .C(men_men_n45_), .D(h), .Y(men_men_n738_));
  AN2        u0710(.A(l), .B(k), .Y(men_men_n739_));
  NA4        u0711(.A(men_men_n739_), .B(men_men_n111_), .C(men_men_n74_), .D(men_men_n221_), .Y(men_men_n740_));
  OAI210     u0712(.A0(men_men_n738_), .A1(g), .B0(men_men_n740_), .Y(men_men_n741_));
  NA2        u0713(.A(men_men_n741_), .B(men_men_n737_), .Y(men_men_n742_));
  NA4        u0714(.A(men_men_n742_), .B(men_men_n736_), .C(men_men_n731_), .D(men_men_n365_), .Y(men_men_n743_));
  AN2        u0715(.A(men_men_n562_), .B(men_men_n97_), .Y(men_men_n744_));
  NO4        u0716(.A(men_men_n181_), .B(men_men_n410_), .C(men_men_n115_), .D(g), .Y(men_men_n745_));
  AOI210     u0717(.A0(men_men_n745_), .A1(men_men_n735_), .B0(men_men_n546_), .Y(men_men_n746_));
  NO2        u0718(.A(men_men_n38_), .B(men_men_n220_), .Y(men_men_n747_));
  AOI220     u0719(.A0(men_men_n649_), .A1(men_men_n362_), .B0(men_men_n747_), .B1(men_men_n593_), .Y(men_men_n748_));
  NAi31      u0720(.An(men_men_n744_), .B(men_men_n748_), .C(men_men_n746_), .Y(men_men_n749_));
  NO2        u0721(.A(men_men_n565_), .B(men_men_n35_), .Y(men_men_n750_));
  OAI210     u0722(.A0(men_men_n581_), .A1(men_men_n47_), .B0(men_men_n139_), .Y(men_men_n751_));
  NO2        u0723(.A(men_men_n509_), .B(men_men_n136_), .Y(men_men_n752_));
  AOI210     u0724(.A0(men_men_n752_), .A1(men_men_n751_), .B0(men_men_n750_), .Y(men_men_n753_));
  NO3        u0725(.A(men_men_n329_), .B(men_men_n135_), .C(men_men_n41_), .Y(men_men_n754_));
  NAi21      u0726(.An(men_men_n754_), .B(men_men_n740_), .Y(men_men_n755_));
  NA2        u0727(.A(men_men_n728_), .B(men_men_n140_), .Y(men_men_n756_));
  AOI220     u0728(.A0(men_men_n756_), .A1(men_men_n420_), .B0(men_men_n755_), .B1(men_men_n77_), .Y(men_men_n757_));
  OAI210     u0729(.A0(men_men_n753_), .A1(men_men_n88_), .B0(men_men_n757_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n378_), .B(men_men_n43_), .Y(men_men_n759_));
  NA3        u0731(.A(men_men_n718_), .B(men_men_n348_), .C(men_men_n402_), .Y(men_men_n760_));
  NA2        u0732(.A(men_men_n739_), .B(men_men_n228_), .Y(men_men_n761_));
  NO2        u0733(.A(men_men_n761_), .B(men_men_n341_), .Y(men_men_n762_));
  AOI210     u0734(.A0(men_men_n762_), .A1(men_men_n709_), .B0(men_men_n515_), .Y(men_men_n763_));
  NA3        u0735(.A(m), .B(l), .C(k), .Y(men_men_n764_));
  AOI210     u0736(.A0(men_men_n689_), .A1(men_men_n687_), .B0(men_men_n764_), .Y(men_men_n765_));
  NO2        u0737(.A(men_men_n564_), .B(men_men_n279_), .Y(men_men_n766_));
  NOi21      u0738(.An(men_men_n766_), .B(men_men_n558_), .Y(men_men_n767_));
  NA4        u0739(.A(men_men_n116_), .B(l), .C(k), .D(men_men_n88_), .Y(men_men_n768_));
  NA3        u0740(.A(men_men_n124_), .B(men_men_n429_), .C(i), .Y(men_men_n769_));
  NO2        u0741(.A(men_men_n769_), .B(men_men_n768_), .Y(men_men_n770_));
  NO3        u0742(.A(men_men_n770_), .B(men_men_n767_), .C(men_men_n765_), .Y(men_men_n771_));
  NA4        u0743(.A(men_men_n771_), .B(men_men_n763_), .C(men_men_n760_), .D(men_men_n759_), .Y(men_men_n772_));
  NO4        u0744(.A(men_men_n772_), .B(men_men_n758_), .C(men_men_n749_), .D(men_men_n743_), .Y(men_men_n773_));
  NA2        u0745(.A(men_men_n649_), .B(men_men_n411_), .Y(men_men_n774_));
  NOi31      u0746(.An(g), .B(h), .C(f), .Y(men_men_n775_));
  NA2        u0747(.A(men_men_n665_), .B(men_men_n775_), .Y(men_men_n776_));
  AO210      u0748(.A0(men_men_n776_), .A1(men_men_n620_), .B0(men_men_n566_), .Y(men_men_n777_));
  NO3        u0749(.A(men_men_n414_), .B(men_men_n552_), .C(h), .Y(men_men_n778_));
  AOI210     u0750(.A0(men_men_n778_), .A1(men_men_n116_), .B0(men_men_n526_), .Y(men_men_n779_));
  NA4        u0751(.A(men_men_n779_), .B(men_men_n777_), .C(men_men_n774_), .D(men_men_n258_), .Y(men_men_n780_));
  NA2        u0752(.A(men_men_n739_), .B(men_men_n74_), .Y(men_men_n781_));
  NO4        u0753(.A(men_men_n717_), .B(men_men_n181_), .C(n), .D(i), .Y(men_men_n782_));
  NOi21      u0754(.An(h), .B(j), .Y(men_men_n783_));
  NA2        u0755(.A(men_men_n783_), .B(f), .Y(men_men_n784_));
  NO2        u0756(.A(men_men_n784_), .B(men_men_n252_), .Y(men_men_n785_));
  NO3        u0757(.A(men_men_n785_), .B(men_men_n782_), .C(men_men_n720_), .Y(men_men_n786_));
  OAI220     u0758(.A0(men_men_n786_), .A1(men_men_n781_), .B0(men_men_n622_), .B1(men_men_n61_), .Y(men_men_n787_));
  AOI210     u0759(.A0(men_men_n780_), .A1(l), .B0(men_men_n787_), .Y(men_men_n788_));
  NO2        u0760(.A(j), .B(i), .Y(men_men_n789_));
  NA3        u0761(.A(men_men_n789_), .B(men_men_n81_), .C(l), .Y(men_men_n790_));
  NA2        u0762(.A(men_men_n789_), .B(men_men_n33_), .Y(men_men_n791_));
  NA2        u0763(.A(men_men_n439_), .B(men_men_n124_), .Y(men_men_n792_));
  OA220      u0764(.A0(men_men_n792_), .A1(men_men_n791_), .B0(men_men_n790_), .B1(men_men_n618_), .Y(men_men_n793_));
  NO3        u0765(.A(men_men_n157_), .B(men_men_n49_), .C(men_men_n113_), .Y(men_men_n794_));
  NO3        u0766(.A(men_men_n570_), .B(men_men_n155_), .C(men_men_n74_), .Y(men_men_n795_));
  NO3        u0767(.A(men_men_n509_), .B(men_men_n458_), .C(j), .Y(men_men_n796_));
  OAI210     u0768(.A0(men_men_n795_), .A1(men_men_n794_), .B0(men_men_n796_), .Y(men_men_n797_));
  OAI210     u0769(.A0(men_men_n776_), .A1(men_men_n61_), .B0(men_men_n797_), .Y(men_men_n798_));
  NA2        u0770(.A(k), .B(j), .Y(men_men_n799_));
  NO3        u0771(.A(men_men_n308_), .B(men_men_n799_), .C(men_men_n40_), .Y(men_men_n800_));
  AOI210     u0772(.A0(men_men_n557_), .A1(n), .B0(men_men_n580_), .Y(men_men_n801_));
  NA2        u0773(.A(men_men_n801_), .B(men_men_n582_), .Y(men_men_n802_));
  AN3        u0774(.A(men_men_n802_), .B(men_men_n800_), .C(men_men_n100_), .Y(men_men_n803_));
  NO3        u0775(.A(men_men_n181_), .B(men_men_n410_), .C(men_men_n115_), .Y(men_men_n804_));
  AOI220     u0776(.A0(men_men_n804_), .A1(men_men_n253_), .B0(men_men_n643_), .B1(men_men_n319_), .Y(men_men_n805_));
  NAi31      u0777(.An(men_men_n638_), .B(men_men_n94_), .C(men_men_n85_), .Y(men_men_n806_));
  NA2        u0778(.A(men_men_n806_), .B(men_men_n805_), .Y(men_men_n807_));
  NO2        u0779(.A(men_men_n308_), .B(men_men_n140_), .Y(men_men_n808_));
  AOI220     u0780(.A0(men_men_n808_), .A1(men_men_n649_), .B0(men_men_n754_), .B1(men_men_n737_), .Y(men_men_n809_));
  NO2        u0781(.A(men_men_n764_), .B(men_men_n92_), .Y(men_men_n810_));
  NA2        u0782(.A(men_men_n810_), .B(men_men_n617_), .Y(men_men_n811_));
  NO2        u0783(.A(men_men_n619_), .B(men_men_n120_), .Y(men_men_n812_));
  OAI210     u0784(.A0(men_men_n812_), .A1(men_men_n796_), .B0(men_men_n705_), .Y(men_men_n813_));
  NA3        u0785(.A(men_men_n813_), .B(men_men_n811_), .C(men_men_n809_), .Y(men_men_n814_));
  OR4        u0786(.A(men_men_n814_), .B(men_men_n807_), .C(men_men_n803_), .D(men_men_n798_), .Y(men_men_n815_));
  NA3        u0787(.A(men_men_n801_), .B(men_men_n582_), .C(men_men_n581_), .Y(men_men_n816_));
  NA4        u0788(.A(men_men_n816_), .B(men_men_n223_), .C(men_men_n471_), .D(men_men_n34_), .Y(men_men_n817_));
  NO4        u0789(.A(men_men_n509_), .B(men_men_n453_), .C(j), .D(f), .Y(men_men_n818_));
  OAI220     u0790(.A0(men_men_n738_), .A1(men_men_n730_), .B0(men_men_n346_), .B1(men_men_n38_), .Y(men_men_n819_));
  AOI210     u0791(.A0(men_men_n818_), .A1(men_men_n264_), .B0(men_men_n819_), .Y(men_men_n820_));
  NA3        u0792(.A(men_men_n573_), .B(men_men_n301_), .C(h), .Y(men_men_n821_));
  NOi21      u0793(.An(men_men_n705_), .B(men_men_n821_), .Y(men_men_n822_));
  NO2        u0794(.A(men_men_n93_), .B(men_men_n47_), .Y(men_men_n823_));
  OAI220     u0795(.A0(men_men_n821_), .A1(men_men_n636_), .B0(men_men_n790_), .B1(men_men_n697_), .Y(men_men_n824_));
  AOI210     u0796(.A0(men_men_n823_), .A1(men_men_n671_), .B0(men_men_n824_), .Y(men_men_n825_));
  NAi41      u0797(.An(men_men_n822_), .B(men_men_n825_), .C(men_men_n820_), .D(men_men_n817_), .Y(men_men_n826_));
  OR2        u0798(.A(men_men_n810_), .B(men_men_n97_), .Y(men_men_n827_));
  AOI220     u0799(.A0(men_men_n827_), .A1(men_men_n243_), .B0(men_men_n796_), .B1(men_men_n663_), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n688_), .B(men_men_n74_), .Y(men_men_n829_));
  AOI210     u0801(.A0(men_men_n818_), .A1(men_men_n829_), .B0(men_men_n350_), .Y(men_men_n830_));
  OAI210     u0802(.A0(men_men_n764_), .A1(men_men_n686_), .B0(men_men_n545_), .Y(men_men_n831_));
  NA3        u0803(.A(men_men_n256_), .B(men_men_n59_), .C(b), .Y(men_men_n832_));
  AOI220     u0804(.A0(men_men_n635_), .A1(men_men_n29_), .B0(men_men_n487_), .B1(men_men_n85_), .Y(men_men_n833_));
  NA2        u0805(.A(men_men_n833_), .B(men_men_n832_), .Y(men_men_n834_));
  NO2        u0806(.A(men_men_n821_), .B(men_men_n514_), .Y(men_men_n835_));
  AOI210     u0807(.A0(men_men_n834_), .A1(men_men_n831_), .B0(men_men_n835_), .Y(men_men_n836_));
  NA3        u0808(.A(men_men_n836_), .B(men_men_n830_), .C(men_men_n828_), .Y(men_men_n837_));
  NOi41      u0809(.An(men_men_n793_), .B(men_men_n837_), .C(men_men_n826_), .D(men_men_n815_), .Y(men_men_n838_));
  OR3        u0810(.A(men_men_n738_), .B(men_men_n238_), .C(g), .Y(men_men_n839_));
  NO3        u0811(.A(men_men_n356_), .B(men_men_n310_), .C(men_men_n115_), .Y(men_men_n840_));
  NA2        u0812(.A(men_men_n840_), .B(men_men_n802_), .Y(men_men_n841_));
  NA2        u0813(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n842_));
  NO3        u0814(.A(men_men_n842_), .B(men_men_n791_), .C(men_men_n285_), .Y(men_men_n843_));
  NO3        u0815(.A(men_men_n552_), .B(men_men_n95_), .C(h), .Y(men_men_n844_));
  AOI210     u0816(.A0(men_men_n844_), .A1(men_men_n733_), .B0(men_men_n843_), .Y(men_men_n845_));
  NA4        u0817(.A(men_men_n845_), .B(men_men_n841_), .C(men_men_n839_), .D(men_men_n422_), .Y(men_men_n846_));
  OR2        u0818(.A(men_men_n686_), .B(men_men_n93_), .Y(men_men_n847_));
  NOi31      u0819(.An(b), .B(d), .C(a), .Y(men_men_n848_));
  NO2        u0820(.A(men_men_n848_), .B(men_men_n633_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n849_), .B(n), .Y(men_men_n850_));
  NOi21      u0822(.An(men_men_n833_), .B(men_men_n850_), .Y(men_men_n851_));
  OAI220     u0823(.A0(men_men_n851_), .A1(men_men_n847_), .B0(men_men_n821_), .B1(men_men_n634_), .Y(men_men_n852_));
  NO2        u0824(.A(men_men_n581_), .B(men_men_n85_), .Y(men_men_n853_));
  NO3        u0825(.A(men_men_n648_), .B(men_men_n341_), .C(men_men_n120_), .Y(men_men_n854_));
  NOi21      u0826(.An(men_men_n854_), .B(men_men_n167_), .Y(men_men_n855_));
  AOI210     u0827(.A0(men_men_n840_), .A1(men_men_n853_), .B0(men_men_n855_), .Y(men_men_n856_));
  OAI210     u0828(.A0(men_men_n738_), .A1(men_men_n412_), .B0(men_men_n856_), .Y(men_men_n857_));
  NO2        u0829(.A(men_men_n717_), .B(n), .Y(men_men_n858_));
  AOI220     u0830(.A0(men_men_n808_), .A1(men_men_n693_), .B0(men_men_n858_), .B1(men_men_n729_), .Y(men_men_n859_));
  NO2        u0831(.A(men_men_n336_), .B(men_men_n242_), .Y(men_men_n860_));
  OAI210     u0832(.A0(men_men_n97_), .A1(men_men_n94_), .B0(men_men_n860_), .Y(men_men_n861_));
  NA2        u0833(.A(men_men_n124_), .B(men_men_n85_), .Y(men_men_n862_));
  AOI210     u0834(.A0(men_men_n443_), .A1(men_men_n435_), .B0(men_men_n862_), .Y(men_men_n863_));
  NAi21      u0835(.An(men_men_n863_), .B(men_men_n861_), .Y(men_men_n864_));
  NA2        u0836(.A(men_men_n762_), .B(men_men_n34_), .Y(men_men_n865_));
  NAi21      u0837(.An(men_men_n768_), .B(men_men_n454_), .Y(men_men_n866_));
  NO2        u0838(.A(men_men_n279_), .B(i), .Y(men_men_n867_));
  NA2        u0839(.A(men_men_n745_), .B(men_men_n364_), .Y(men_men_n868_));
  OAI210     u0840(.A0(men_men_n625_), .A1(men_men_n624_), .B0(men_men_n379_), .Y(men_men_n869_));
  AN3        u0841(.A(men_men_n869_), .B(men_men_n868_), .C(men_men_n866_), .Y(men_men_n870_));
  NAi41      u0842(.An(men_men_n864_), .B(men_men_n870_), .C(men_men_n865_), .D(men_men_n859_), .Y(men_men_n871_));
  NO4        u0843(.A(men_men_n871_), .B(men_men_n857_), .C(men_men_n852_), .D(men_men_n846_), .Y(men_men_n872_));
  NA4        u0844(.A(men_men_n872_), .B(men_men_n838_), .C(men_men_n788_), .D(men_men_n773_), .Y(men09));
  INV        u0845(.A(men_men_n125_), .Y(men_men_n874_));
  NA2        u0846(.A(f), .B(e), .Y(men_men_n875_));
  NO2        u0847(.A(men_men_n232_), .B(men_men_n115_), .Y(men_men_n876_));
  NA2        u0848(.A(men_men_n876_), .B(g), .Y(men_men_n877_));
  NA4        u0849(.A(men_men_n322_), .B(men_men_n496_), .C(men_men_n267_), .D(men_men_n122_), .Y(men_men_n878_));
  AOI210     u0850(.A0(men_men_n878_), .A1(g), .B0(men_men_n493_), .Y(men_men_n879_));
  AOI210     u0851(.A0(men_men_n879_), .A1(men_men_n877_), .B0(men_men_n875_), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n464_), .B(e), .Y(men_men_n881_));
  NO2        u0853(.A(men_men_n881_), .B(men_men_n536_), .Y(men_men_n882_));
  AOI210     u0854(.A0(men_men_n880_), .A1(men_men_n874_), .B0(men_men_n882_), .Y(men_men_n883_));
  NO2        u0855(.A(men_men_n210_), .B(men_men_n220_), .Y(men_men_n884_));
  NA3        u0856(.A(m), .B(l), .C(i), .Y(men_men_n885_));
  OAI220     u0857(.A0(men_men_n619_), .A1(men_men_n885_), .B0(men_men_n369_), .B1(men_men_n553_), .Y(men_men_n886_));
  NA4        u0858(.A(men_men_n89_), .B(men_men_n88_), .C(g), .D(f), .Y(men_men_n887_));
  NAi31      u0859(.An(men_men_n886_), .B(men_men_n887_), .C(men_men_n459_), .Y(men_men_n888_));
  OA210      u0860(.A0(men_men_n888_), .A1(men_men_n884_), .B0(men_men_n593_), .Y(men_men_n889_));
  NA3        u0861(.A(men_men_n847_), .B(men_men_n595_), .C(men_men_n545_), .Y(men_men_n890_));
  OA210      u0862(.A0(men_men_n890_), .A1(men_men_n889_), .B0(men_men_n850_), .Y(men_men_n891_));
  INV        u0863(.A(men_men_n353_), .Y(men_men_n892_));
  NO2        u0864(.A(men_men_n131_), .B(men_men_n129_), .Y(men_men_n893_));
  NOi31      u0865(.An(k), .B(m), .C(l), .Y(men_men_n894_));
  NO2        u0866(.A(men_men_n355_), .B(men_men_n894_), .Y(men_men_n895_));
  AOI210     u0867(.A0(men_men_n895_), .A1(men_men_n893_), .B0(men_men_n628_), .Y(men_men_n896_));
  NA2        u0868(.A(men_men_n832_), .B(men_men_n346_), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n357_), .B(men_men_n359_), .Y(men_men_n898_));
  OAI210     u0870(.A0(men_men_n210_), .A1(men_men_n220_), .B0(men_men_n898_), .Y(men_men_n899_));
  AOI220     u0871(.A0(men_men_n899_), .A1(men_men_n897_), .B0(men_men_n896_), .B1(men_men_n892_), .Y(men_men_n900_));
  NA3        u0872(.A(men_men_n1602_), .B(men_men_n196_), .C(men_men_n31_), .Y(men_men_n901_));
  NA4        u0873(.A(men_men_n901_), .B(men_men_n900_), .C(men_men_n650_), .D(men_men_n83_), .Y(men_men_n902_));
  NO2        u0874(.A(men_men_n615_), .B(men_men_n522_), .Y(men_men_n903_));
  NA2        u0875(.A(men_men_n903_), .B(men_men_n196_), .Y(men_men_n904_));
  NOi21      u0876(.An(f), .B(d), .Y(men_men_n905_));
  NA2        u0877(.A(men_men_n905_), .B(m), .Y(men_men_n906_));
  NO2        u0878(.A(men_men_n906_), .B(men_men_n52_), .Y(men_men_n907_));
  NOi32      u0879(.An(g), .Bn(f), .C(d), .Y(men_men_n908_));
  NA4        u0880(.A(men_men_n908_), .B(men_men_n635_), .C(men_men_n29_), .D(m), .Y(men_men_n909_));
  NOi21      u0881(.An(men_men_n323_), .B(men_men_n909_), .Y(men_men_n910_));
  AOI210     u0882(.A0(men_men_n907_), .A1(men_men_n571_), .B0(men_men_n910_), .Y(men_men_n911_));
  NA3        u0883(.A(men_men_n322_), .B(men_men_n267_), .C(men_men_n122_), .Y(men_men_n912_));
  AN2        u0884(.A(f), .B(d), .Y(men_men_n913_));
  NA3        u0885(.A(men_men_n501_), .B(men_men_n913_), .C(men_men_n85_), .Y(men_men_n914_));
  NO3        u0886(.A(men_men_n914_), .B(men_men_n74_), .C(men_men_n221_), .Y(men_men_n915_));
  NO2        u0887(.A(men_men_n294_), .B(men_men_n56_), .Y(men_men_n916_));
  OAI210     u0888(.A0(men_men_n916_), .A1(men_men_n912_), .B0(men_men_n915_), .Y(men_men_n917_));
  NAi41      u0889(.An(men_men_n513_), .B(men_men_n917_), .C(men_men_n911_), .D(men_men_n904_), .Y(men_men_n918_));
  NO4        u0890(.A(men_men_n648_), .B(men_men_n136_), .C(men_men_n341_), .D(men_men_n158_), .Y(men_men_n919_));
  NO2        u0891(.A(men_men_n680_), .B(men_men_n341_), .Y(men_men_n920_));
  AN2        u0892(.A(men_men_n920_), .B(men_men_n709_), .Y(men_men_n921_));
  NO3        u0893(.A(men_men_n921_), .B(men_men_n919_), .C(men_men_n240_), .Y(men_men_n922_));
  NA2        u0894(.A(men_men_n633_), .B(men_men_n85_), .Y(men_men_n923_));
  OAI220     u0895(.A0(men_men_n898_), .A1(men_men_n923_), .B0(men_men_n832_), .B1(men_men_n459_), .Y(men_men_n924_));
  NA3        u0896(.A(men_men_n166_), .B(men_men_n111_), .C(men_men_n110_), .Y(men_men_n925_));
  OAI220     u0897(.A0(men_men_n914_), .A1(men_men_n448_), .B0(men_men_n353_), .B1(men_men_n925_), .Y(men_men_n926_));
  NOi41      u0898(.An(men_men_n230_), .B(men_men_n926_), .C(men_men_n924_), .D(men_men_n317_), .Y(men_men_n927_));
  NA2        u0899(.A(c), .B(men_men_n119_), .Y(men_men_n928_));
  NO2        u0900(.A(men_men_n928_), .B(men_men_n426_), .Y(men_men_n929_));
  NA3        u0901(.A(men_men_n929_), .B(men_men_n534_), .C(f), .Y(men_men_n930_));
  OR2        u0902(.A(men_men_n686_), .B(men_men_n567_), .Y(men_men_n931_));
  OAI210     u0903(.A0(men_men_n598_), .A1(men_men_n644_), .B0(men_men_n931_), .Y(men_men_n932_));
  NA2        u0904(.A(men_men_n849_), .B(men_men_n114_), .Y(men_men_n933_));
  NA2        u0905(.A(men_men_n933_), .B(men_men_n932_), .Y(men_men_n934_));
  NA4        u0906(.A(men_men_n934_), .B(men_men_n930_), .C(men_men_n927_), .D(men_men_n922_), .Y(men_men_n935_));
  NO4        u0907(.A(men_men_n935_), .B(men_men_n918_), .C(men_men_n902_), .D(men_men_n891_), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n115_), .B(j), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n937_), .B(men_men_n149_), .Y(men_men_n938_));
  OAI210     u0910(.A0(men_men_n938_), .A1(men_men_n876_), .B0(g), .Y(men_men_n939_));
  AOI210     u0911(.A0(men_men_n939_), .A1(men_men_n302_), .B0(men_men_n914_), .Y(men_men_n940_));
  AOI210     u0912(.A0(men_men_n832_), .A1(men_men_n346_), .B0(men_men_n887_), .Y(men_men_n941_));
  NO2        u0913(.A(men_men_n140_), .B(men_men_n136_), .Y(men_men_n942_));
  NO2        u0914(.A(men_men_n237_), .B(men_men_n231_), .Y(men_men_n943_));
  AOI220     u0915(.A0(men_men_n943_), .A1(men_men_n234_), .B0(men_men_n315_), .B1(men_men_n942_), .Y(men_men_n944_));
  NO2        u0916(.A(men_men_n448_), .B(men_men_n875_), .Y(men_men_n945_));
  NA2        u0917(.A(men_men_n945_), .B(men_men_n587_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n946_), .B(men_men_n944_), .Y(men_men_n947_));
  NA2        u0919(.A(e), .B(d), .Y(men_men_n948_));
  AOI210     u0920(.A0(men_men_n540_), .A1(men_men_n187_), .B0(men_men_n237_), .Y(men_men_n949_));
  AOI210     u0921(.A0(men_men_n649_), .A1(men_men_n362_), .B0(men_men_n949_), .Y(men_men_n950_));
  NA2        u0922(.A(men_men_n294_), .B(men_men_n172_), .Y(men_men_n951_));
  NA3        u0923(.A(men_men_n915_), .B(men_men_n951_), .C(men_men_n56_), .Y(men_men_n952_));
  NA3        u0924(.A(men_men_n175_), .B(men_men_n86_), .C(men_men_n34_), .Y(men_men_n953_));
  NA3        u0925(.A(men_men_n953_), .B(men_men_n952_), .C(men_men_n950_), .Y(men_men_n954_));
  NO4        u0926(.A(men_men_n954_), .B(men_men_n947_), .C(men_men_n941_), .D(men_men_n940_), .Y(men_men_n955_));
  NA2        u0927(.A(men_men_n892_), .B(men_men_n31_), .Y(men_men_n956_));
  AO210      u0928(.A0(men_men_n956_), .A1(men_men_n730_), .B0(men_men_n224_), .Y(men_men_n957_));
  OAI220     u0929(.A0(men_men_n648_), .A1(men_men_n60_), .B0(men_men_n310_), .B1(j), .Y(men_men_n958_));
  NA2        u0930(.A(men_men_n958_), .B(men_men_n920_), .Y(men_men_n959_));
  OAI210     u0931(.A0(men_men_n881_), .A1(men_men_n179_), .B0(men_men_n959_), .Y(men_men_n960_));
  OAI210     u0932(.A0(men_men_n876_), .A1(men_men_n951_), .B0(men_men_n908_), .Y(men_men_n961_));
  NO2        u0933(.A(men_men_n961_), .B(men_men_n636_), .Y(men_men_n962_));
  AOI210     u0934(.A0(men_men_n121_), .A1(men_men_n120_), .B0(men_men_n266_), .Y(men_men_n963_));
  NO2        u0935(.A(men_men_n963_), .B(men_men_n909_), .Y(men_men_n964_));
  AO210      u0936(.A0(men_men_n897_), .A1(men_men_n886_), .B0(men_men_n964_), .Y(men_men_n965_));
  NOi31      u0937(.An(men_men_n571_), .B(men_men_n906_), .C(men_men_n302_), .Y(men_men_n966_));
  NO4        u0938(.A(men_men_n966_), .B(men_men_n965_), .C(men_men_n962_), .D(men_men_n960_), .Y(men_men_n967_));
  NA2        u0939(.A(men_men_n479_), .B(e), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n458_), .B(men_men_n70_), .Y(men_men_n969_));
  OAI210     u0941(.A0(men_men_n890_), .A1(men_men_n969_), .B0(men_men_n733_), .Y(men_men_n970_));
  AN4        u0942(.A(men_men_n970_), .B(men_men_n968_), .C(men_men_n967_), .D(men_men_n957_), .Y(men_men_n971_));
  NA4        u0943(.A(men_men_n971_), .B(men_men_n955_), .C(men_men_n936_), .D(men_men_n883_), .Y(men12));
  NO2        u0944(.A(men_men_n474_), .B(c), .Y(men_men_n973_));
  NO4        u0945(.A(men_men_n463_), .B(men_men_n259_), .C(men_men_n611_), .D(men_men_n221_), .Y(men_men_n974_));
  NA2        u0946(.A(men_men_n974_), .B(men_men_n973_), .Y(men_men_n975_));
  NA2        u0947(.A(men_men_n571_), .B(men_men_n969_), .Y(men_men_n976_));
  NO3        u0948(.A(men_men_n474_), .B(men_men_n85_), .C(men_men_n119_), .Y(men_men_n977_));
  NO2        u0949(.A(men_men_n893_), .B(men_men_n369_), .Y(men_men_n978_));
  NO2        u0950(.A(men_men_n686_), .B(men_men_n396_), .Y(men_men_n979_));
  AOI220     u0951(.A0(men_men_n979_), .A1(men_men_n569_), .B0(men_men_n978_), .B1(men_men_n977_), .Y(men_men_n980_));
  NA4        u0952(.A(men_men_n980_), .B(men_men_n976_), .C(men_men_n975_), .D(men_men_n462_), .Y(men_men_n981_));
  AOI210     u0953(.A0(men_men_n239_), .A1(men_men_n352_), .B0(men_men_n207_), .Y(men_men_n982_));
  OR2        u0954(.A(men_men_n982_), .B(men_men_n974_), .Y(men_men_n983_));
  AOI210     u0955(.A0(men_men_n349_), .A1(men_men_n408_), .B0(men_men_n221_), .Y(men_men_n984_));
  OAI210     u0956(.A0(men_men_n984_), .A1(men_men_n983_), .B0(men_men_n421_), .Y(men_men_n985_));
  NO2        u0957(.A(men_men_n668_), .B(men_men_n269_), .Y(men_men_n986_));
  NO2        u0958(.A(men_men_n619_), .B(men_men_n885_), .Y(men_men_n987_));
  AOI220     u0959(.A0(men_men_n987_), .A1(men_men_n593_), .B0(men_men_n860_), .B1(men_men_n986_), .Y(men_men_n988_));
  NO2        u0960(.A(men_men_n157_), .B(men_men_n242_), .Y(men_men_n989_));
  NA3        u0961(.A(men_men_n989_), .B(men_men_n245_), .C(i), .Y(men_men_n990_));
  NA3        u0962(.A(men_men_n990_), .B(men_men_n988_), .C(men_men_n985_), .Y(men_men_n991_));
  OR2        u0963(.A(men_men_n337_), .B(men_men_n977_), .Y(men_men_n992_));
  NA2        u0964(.A(men_men_n992_), .B(men_men_n370_), .Y(men_men_n993_));
  NO3        u0965(.A(men_men_n136_), .B(men_men_n158_), .C(men_men_n221_), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n994_), .B(men_men_n557_), .Y(men_men_n995_));
  NA4        u0967(.A(men_men_n464_), .B(men_men_n456_), .C(men_men_n188_), .D(g), .Y(men_men_n996_));
  NA3        u0968(.A(men_men_n996_), .B(men_men_n995_), .C(men_men_n993_), .Y(men_men_n997_));
  NO3        u0969(.A(men_men_n691_), .B(men_men_n93_), .C(men_men_n45_), .Y(men_men_n998_));
  NO4        u0970(.A(men_men_n998_), .B(men_men_n997_), .C(men_men_n991_), .D(men_men_n981_), .Y(men_men_n999_));
  NO2        u0971(.A(men_men_n386_), .B(men_men_n385_), .Y(men_men_n1000_));
  NA2        u0972(.A(men_men_n616_), .B(men_men_n72_), .Y(men_men_n1001_));
  NA2        u0973(.A(men_men_n581_), .B(men_men_n150_), .Y(men_men_n1002_));
  NOi21      u0974(.An(men_men_n34_), .B(men_men_n680_), .Y(men_men_n1003_));
  AOI220     u0975(.A0(men_men_n1003_), .A1(men_men_n1002_), .B0(men_men_n1001_), .B1(men_men_n1000_), .Y(men_men_n1004_));
  OAI210     u0976(.A0(men_men_n257_), .A1(men_men_n45_), .B0(men_men_n1004_), .Y(men_men_n1005_));
  NA2        u0977(.A(men_men_n454_), .B(men_men_n271_), .Y(men_men_n1006_));
  NO3        u0978(.A(men_men_n862_), .B(men_men_n90_), .C(men_men_n426_), .Y(men_men_n1007_));
  NAi31      u0979(.An(men_men_n1007_), .B(men_men_n1006_), .C(men_men_n333_), .Y(men_men_n1008_));
  NO2        u0980(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n1009_));
  NO2        u0981(.A(men_men_n529_), .B(men_men_n310_), .Y(men_men_n1010_));
  NO2        u0982(.A(men_men_n1010_), .B(men_men_n382_), .Y(men_men_n1011_));
  NO2        u0983(.A(men_men_n1011_), .B(men_men_n150_), .Y(men_men_n1012_));
  NA2        u0984(.A(men_men_n659_), .B(men_men_n379_), .Y(men_men_n1013_));
  OAI210     u0985(.A0(men_men_n769_), .A1(men_men_n1013_), .B0(men_men_n383_), .Y(men_men_n1014_));
  NO4        u0986(.A(men_men_n1014_), .B(men_men_n1012_), .C(men_men_n1008_), .D(men_men_n1005_), .Y(men_men_n1015_));
  NA2        u0987(.A(men_men_n362_), .B(g), .Y(men_men_n1016_));
  NA2        u0988(.A(men_men_n169_), .B(i), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n46_), .B(i), .Y(men_men_n1018_));
  OAI220     u0990(.A0(men_men_n1018_), .A1(men_men_n206_), .B0(men_men_n1017_), .B1(men_men_n93_), .Y(men_men_n1019_));
  AOI210     u0991(.A0(men_men_n437_), .A1(men_men_n37_), .B0(men_men_n1019_), .Y(men_men_n1020_));
  NO2        u0992(.A(men_men_n150_), .B(men_men_n85_), .Y(men_men_n1021_));
  OR2        u0993(.A(men_men_n1021_), .B(men_men_n580_), .Y(men_men_n1022_));
  NA2        u0994(.A(men_men_n581_), .B(men_men_n400_), .Y(men_men_n1023_));
  AOI210     u0995(.A0(men_men_n1023_), .A1(n), .B0(men_men_n1022_), .Y(men_men_n1024_));
  OAI220     u0996(.A0(men_men_n1024_), .A1(men_men_n1016_), .B0(men_men_n1020_), .B1(men_men_n346_), .Y(men_men_n1025_));
  NO2        u0997(.A(men_men_n686_), .B(men_men_n522_), .Y(men_men_n1026_));
  NA3        u0998(.A(men_men_n357_), .B(men_men_n654_), .C(i), .Y(men_men_n1027_));
  OAI210     u0999(.A0(men_men_n458_), .A1(men_men_n322_), .B0(men_men_n1027_), .Y(men_men_n1028_));
  OAI220     u1000(.A0(men_men_n1028_), .A1(men_men_n1026_), .B0(men_men_n705_), .B1(men_men_n795_), .Y(men_men_n1029_));
  NA2        u1001(.A(men_men_n637_), .B(men_men_n116_), .Y(men_men_n1030_));
  OR3        u1002(.A(men_men_n322_), .B(men_men_n453_), .C(f), .Y(men_men_n1031_));
  NA3        u1003(.A(men_men_n654_), .B(men_men_n81_), .C(i), .Y(men_men_n1032_));
  OA220      u1004(.A0(men_men_n1032_), .A1(men_men_n1030_), .B0(men_men_n1031_), .B1(men_men_n618_), .Y(men_men_n1033_));
  NA3        u1005(.A(men_men_n338_), .B(men_men_n121_), .C(g), .Y(men_men_n1034_));
  AOI210     u1006(.A0(men_men_n702_), .A1(men_men_n1034_), .B0(m), .Y(men_men_n1035_));
  NA2        u1007(.A(men_men_n978_), .B(men_men_n337_), .Y(men_men_n1036_));
  NA2        u1008(.A(men_men_n721_), .B(men_men_n923_), .Y(men_men_n1037_));
  NA2        u1009(.A(men_men_n887_), .B(men_men_n459_), .Y(men_men_n1038_));
  NA2        u1010(.A(i), .B(men_men_n78_), .Y(men_men_n1039_));
  NA3        u1011(.A(men_men_n1039_), .B(men_men_n1032_), .C(men_men_n1031_), .Y(men_men_n1040_));
  AOI220     u1012(.A0(men_men_n1040_), .A1(men_men_n264_), .B0(men_men_n1038_), .B1(men_men_n1037_), .Y(men_men_n1041_));
  NA4        u1013(.A(men_men_n1041_), .B(men_men_n1036_), .C(men_men_n1033_), .D(men_men_n1029_), .Y(men_men_n1042_));
  NO2        u1014(.A(men_men_n396_), .B(men_men_n92_), .Y(men_men_n1043_));
  OAI210     u1015(.A0(men_men_n1043_), .A1(men_men_n986_), .B0(men_men_n243_), .Y(men_men_n1044_));
  NA2        u1016(.A(men_men_n690_), .B(men_men_n89_), .Y(men_men_n1045_));
  NO2        u1017(.A(men_men_n482_), .B(men_men_n221_), .Y(men_men_n1046_));
  AOI220     u1018(.A0(men_men_n1046_), .A1(men_men_n401_), .B0(men_men_n992_), .B1(men_men_n225_), .Y(men_men_n1047_));
  AOI220     u1019(.A0(men_men_n979_), .A1(men_men_n989_), .B0(men_men_n617_), .B1(men_men_n91_), .Y(men_men_n1048_));
  NA4        u1020(.A(men_men_n1048_), .B(men_men_n1047_), .C(men_men_n1045_), .D(men_men_n1044_), .Y(men_men_n1049_));
  OAI210     u1021(.A0(men_men_n1038_), .A1(men_men_n987_), .B0(men_men_n569_), .Y(men_men_n1050_));
  AOI210     u1022(.A0(men_men_n438_), .A1(men_men_n430_), .B0(men_men_n862_), .Y(men_men_n1051_));
  OAI210     u1023(.A0(men_men_n386_), .A1(men_men_n385_), .B0(men_men_n112_), .Y(men_men_n1052_));
  AOI210     u1024(.A0(men_men_n1052_), .A1(men_men_n562_), .B0(men_men_n1051_), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n1035_), .B(men_men_n977_), .Y(men_men_n1054_));
  NO3        u1026(.A(men_men_n937_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1055_));
  AOI220     u1027(.A0(men_men_n1055_), .A1(men_men_n652_), .B0(men_men_n673_), .B1(men_men_n557_), .Y(men_men_n1056_));
  NA4        u1028(.A(men_men_n1056_), .B(men_men_n1054_), .C(men_men_n1053_), .D(men_men_n1050_), .Y(men_men_n1057_));
  NO4        u1029(.A(men_men_n1057_), .B(men_men_n1049_), .C(men_men_n1042_), .D(men_men_n1025_), .Y(men_men_n1058_));
  NAi31      u1030(.An(men_men_n146_), .B(men_men_n439_), .C(n), .Y(men_men_n1059_));
  NO3        u1031(.A(men_men_n129_), .B(men_men_n355_), .C(men_men_n894_), .Y(men_men_n1060_));
  NO2        u1032(.A(men_men_n1060_), .B(men_men_n1059_), .Y(men_men_n1061_));
  NO3        u1033(.A(men_men_n279_), .B(men_men_n146_), .C(men_men_n426_), .Y(men_men_n1062_));
  AOI210     u1034(.A0(men_men_n1062_), .A1(men_men_n523_), .B0(men_men_n1061_), .Y(men_men_n1063_));
  NA2        u1035(.A(men_men_n516_), .B(i), .Y(men_men_n1064_));
  NA2        u1036(.A(men_men_n1064_), .B(men_men_n1063_), .Y(men_men_n1065_));
  NA2        u1037(.A(men_men_n237_), .B(men_men_n180_), .Y(men_men_n1066_));
  NO2        u1038(.A(men_men_n319_), .B(men_men_n464_), .Y(men_men_n1067_));
  NOi31      u1039(.An(men_men_n1066_), .B(men_men_n1067_), .C(men_men_n221_), .Y(men_men_n1068_));
  NAi21      u1040(.An(men_men_n581_), .B(men_men_n1046_), .Y(men_men_n1069_));
  NA2        u1041(.A(men_men_n457_), .B(men_men_n923_), .Y(men_men_n1070_));
  NO3        u1042(.A(men_men_n458_), .B(men_men_n322_), .C(men_men_n74_), .Y(men_men_n1071_));
  NA2        u1043(.A(men_men_n1071_), .B(men_men_n1070_), .Y(men_men_n1072_));
  NA2        u1044(.A(men_men_n1072_), .B(men_men_n1069_), .Y(men_men_n1073_));
  OAI220     u1045(.A0(men_men_n1059_), .A1(men_men_n239_), .B0(men_men_n1027_), .B1(men_men_n634_), .Y(men_men_n1074_));
  NO2        u1046(.A(men_men_n687_), .B(men_men_n396_), .Y(men_men_n1075_));
  NA2        u1047(.A(men_men_n982_), .B(men_men_n973_), .Y(men_men_n1076_));
  NO3        u1048(.A(men_men_n570_), .B(men_men_n155_), .C(men_men_n220_), .Y(men_men_n1077_));
  OAI210     u1049(.A0(men_men_n1077_), .A1(men_men_n551_), .B0(men_men_n397_), .Y(men_men_n1078_));
  OAI220     u1050(.A0(men_men_n979_), .A1(men_men_n987_), .B0(men_men_n571_), .B1(men_men_n447_), .Y(men_men_n1079_));
  NA4        u1051(.A(men_men_n1079_), .B(men_men_n1078_), .C(men_men_n1076_), .D(men_men_n646_), .Y(men_men_n1080_));
  OAI210     u1052(.A0(men_men_n982_), .A1(men_men_n974_), .B0(men_men_n1066_), .Y(men_men_n1081_));
  NA3        u1053(.A(men_men_n1023_), .B(men_men_n511_), .C(men_men_n46_), .Y(men_men_n1082_));
  AOI210     u1054(.A0(men_men_n399_), .A1(men_men_n397_), .B0(men_men_n345_), .Y(men_men_n1083_));
  NA4        u1055(.A(men_men_n1083_), .B(men_men_n1082_), .C(men_men_n1081_), .D(men_men_n280_), .Y(men_men_n1084_));
  OR4        u1056(.A(men_men_n1084_), .B(men_men_n1080_), .C(men_men_n1075_), .D(men_men_n1074_), .Y(men_men_n1085_));
  NO4        u1057(.A(men_men_n1085_), .B(men_men_n1073_), .C(men_men_n1068_), .D(men_men_n1065_), .Y(men_men_n1086_));
  NA4        u1058(.A(men_men_n1086_), .B(men_men_n1058_), .C(men_men_n1015_), .D(men_men_n999_), .Y(men13));
  NA2        u1059(.A(men_men_n46_), .B(men_men_n88_), .Y(men_men_n1088_));
  AN2        u1060(.A(c), .B(b), .Y(men_men_n1089_));
  NA3        u1061(.A(men_men_n256_), .B(men_men_n1089_), .C(m), .Y(men_men_n1090_));
  NO4        u1062(.A(e), .B(men_men_n1090_), .C(men_men_n1088_), .D(men_men_n612_), .Y(men_men_n1091_));
  NA2        u1063(.A(men_men_n271_), .B(men_men_n1089_), .Y(men_men_n1092_));
  NO4        u1064(.A(men_men_n1092_), .B(e), .C(men_men_n1017_), .D(a), .Y(men_men_n1093_));
  NAi32      u1065(.An(d), .Bn(c), .C(e), .Y(men_men_n1094_));
  NA2        u1066(.A(men_men_n145_), .B(men_men_n45_), .Y(men_men_n1095_));
  NO4        u1067(.A(men_men_n1095_), .B(men_men_n1094_), .C(men_men_n619_), .D(men_men_n318_), .Y(men_men_n1096_));
  NA2        u1068(.A(men_men_n694_), .B(men_men_n231_), .Y(men_men_n1097_));
  NA2        u1069(.A(men_men_n429_), .B(men_men_n220_), .Y(men_men_n1098_));
  AN2        u1070(.A(d), .B(c), .Y(men_men_n1099_));
  NA2        u1071(.A(men_men_n1099_), .B(men_men_n119_), .Y(men_men_n1100_));
  NO4        u1072(.A(men_men_n1100_), .B(men_men_n1098_), .C(men_men_n183_), .D(men_men_n176_), .Y(men_men_n1101_));
  NA2        u1073(.A(d), .B(c), .Y(men_men_n1102_));
  NO4        u1074(.A(men_men_n1095_), .B(men_men_n615_), .C(men_men_n1102_), .D(men_men_n318_), .Y(men_men_n1103_));
  AO210      u1075(.A0(men_men_n1101_), .A1(men_men_n1097_), .B0(men_men_n1103_), .Y(men_men_n1104_));
  OR4        u1076(.A(men_men_n1104_), .B(men_men_n1096_), .C(men_men_n1093_), .D(men_men_n1091_), .Y(men_men_n1105_));
  NAi32      u1077(.An(f), .Bn(e), .C(c), .Y(men_men_n1106_));
  OR3        u1078(.A(men_men_n231_), .B(men_men_n183_), .C(men_men_n176_), .Y(men_men_n1107_));
  NO2        u1079(.A(men_men_n1107_), .B(men_men_n1106_), .Y(men_men_n1108_));
  NO2        u1080(.A(men_men_n1102_), .B(men_men_n318_), .Y(men_men_n1109_));
  NO2        u1081(.A(j), .B(men_men_n45_), .Y(men_men_n1110_));
  NA2        u1082(.A(men_men_n656_), .B(men_men_n1110_), .Y(men_men_n1111_));
  NOi21      u1083(.An(men_men_n1109_), .B(men_men_n1111_), .Y(men_men_n1112_));
  NO2        u1084(.A(men_men_n799_), .B(men_men_n115_), .Y(men_men_n1113_));
  NOi41      u1085(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1114_));
  NA2        u1086(.A(men_men_n1114_), .B(men_men_n1113_), .Y(men_men_n1115_));
  NO2        u1087(.A(men_men_n1115_), .B(men_men_n1106_), .Y(men_men_n1116_));
  OR3        u1088(.A(e), .B(d), .C(c), .Y(men_men_n1117_));
  NA3        u1089(.A(k), .B(j), .C(i), .Y(men_men_n1118_));
  NO3        u1090(.A(men_men_n1118_), .B(men_men_n318_), .C(men_men_n92_), .Y(men_men_n1119_));
  OR4        u1091(.A(men_men_n1119_), .B(men_men_n1116_), .C(men_men_n1112_), .D(men_men_n1108_), .Y(men_men_n1120_));
  NA3        u1092(.A(men_men_n490_), .B(men_men_n348_), .C(men_men_n56_), .Y(men_men_n1121_));
  NO2        u1093(.A(men_men_n1121_), .B(men_men_n1111_), .Y(men_men_n1122_));
  NO4        u1094(.A(men_men_n1121_), .B(men_men_n615_), .C(men_men_n471_), .D(men_men_n45_), .Y(men_men_n1123_));
  NO2        u1095(.A(f), .B(c), .Y(men_men_n1124_));
  NOi21      u1096(.An(men_men_n1124_), .B(men_men_n463_), .Y(men_men_n1125_));
  NA2        u1097(.A(men_men_n1125_), .B(men_men_n59_), .Y(men_men_n1126_));
  OR2        u1098(.A(k), .B(i), .Y(men_men_n1127_));
  NO3        u1099(.A(men_men_n1127_), .B(men_men_n249_), .C(l), .Y(men_men_n1128_));
  NOi31      u1100(.An(men_men_n1128_), .B(men_men_n1126_), .C(j), .Y(men_men_n1129_));
  OR3        u1101(.A(men_men_n1129_), .B(men_men_n1123_), .C(men_men_n1122_), .Y(men_men_n1130_));
  OR3        u1102(.A(men_men_n1130_), .B(men_men_n1120_), .C(men_men_n1105_), .Y(men02));
  OR2        u1103(.A(l), .B(k), .Y(men_men_n1132_));
  OR3        u1104(.A(n), .B(m), .C(i), .Y(men_men_n1133_));
  NO4        u1105(.A(men_men_n1133_), .B(h), .C(men_men_n1132_), .D(men_men_n1117_), .Y(men_men_n1134_));
  NOi31      u1106(.An(e), .B(d), .C(c), .Y(men_men_n1135_));
  AOI210     u1107(.A0(men_men_n1119_), .A1(men_men_n1135_), .B0(men_men_n1096_), .Y(men_men_n1136_));
  AN3        u1108(.A(g), .B(f), .C(c), .Y(men_men_n1137_));
  NA3        u1109(.A(men_men_n1137_), .B(men_men_n490_), .C(h), .Y(men_men_n1138_));
  OR2        u1110(.A(men_men_n1118_), .B(men_men_n318_), .Y(men_men_n1139_));
  OR2        u1111(.A(men_men_n1139_), .B(men_men_n1138_), .Y(men_men_n1140_));
  NO3        u1112(.A(men_men_n1121_), .B(men_men_n1095_), .C(men_men_n615_), .Y(men_men_n1141_));
  NO2        u1113(.A(men_men_n1141_), .B(men_men_n1108_), .Y(men_men_n1142_));
  NA3        u1114(.A(l), .B(k), .C(j), .Y(men_men_n1143_));
  NA2        u1115(.A(i), .B(h), .Y(men_men_n1144_));
  NO3        u1116(.A(men_men_n1144_), .B(men_men_n1143_), .C(men_men_n136_), .Y(men_men_n1145_));
  NO3        u1117(.A(men_men_n147_), .B(men_men_n292_), .C(men_men_n221_), .Y(men_men_n1146_));
  AOI210     u1118(.A0(men_men_n1146_), .A1(men_men_n1145_), .B0(men_men_n1112_), .Y(men_men_n1147_));
  NA3        u1119(.A(c), .B(b), .C(a), .Y(men_men_n1148_));
  NO3        u1120(.A(men_men_n1148_), .B(men_men_n948_), .C(men_men_n220_), .Y(men_men_n1149_));
  NO4        u1121(.A(men_men_n1118_), .B(men_men_n310_), .C(men_men_n49_), .D(men_men_n115_), .Y(men_men_n1150_));
  AOI210     u1122(.A0(men_men_n1150_), .A1(men_men_n1149_), .B0(men_men_n1122_), .Y(men_men_n1151_));
  AN4        u1123(.A(men_men_n1151_), .B(men_men_n1147_), .C(men_men_n1142_), .D(men_men_n1140_), .Y(men_men_n1152_));
  NO2        u1124(.A(men_men_n1100_), .B(men_men_n1098_), .Y(men_men_n1153_));
  NA2        u1125(.A(men_men_n1115_), .B(men_men_n1107_), .Y(men_men_n1154_));
  AOI210     u1126(.A0(men_men_n1154_), .A1(men_men_n1153_), .B0(men_men_n1091_), .Y(men_men_n1155_));
  NAi41      u1127(.An(men_men_n1134_), .B(men_men_n1155_), .C(men_men_n1152_), .D(men_men_n1136_), .Y(men03));
  NO2        u1128(.A(men_men_n553_), .B(men_men_n628_), .Y(men_men_n1157_));
  NA4        u1129(.A(men_men_n89_), .B(men_men_n88_), .C(g), .D(men_men_n220_), .Y(men_men_n1158_));
  NA4        u1130(.A(men_men_n603_), .B(m), .C(men_men_n115_), .D(men_men_n220_), .Y(men_men_n1159_));
  NA3        u1131(.A(men_men_n1159_), .B(men_men_n387_), .C(men_men_n1158_), .Y(men_men_n1160_));
  NO3        u1132(.A(men_men_n1160_), .B(men_men_n1157_), .C(men_men_n1052_), .Y(men_men_n1161_));
  NOi41      u1133(.An(men_men_n847_), .B(men_men_n899_), .C(men_men_n888_), .D(men_men_n747_), .Y(men_men_n1162_));
  OAI220     u1134(.A0(men_men_n1162_), .A1(men_men_n721_), .B0(men_men_n1161_), .B1(men_men_n616_), .Y(men_men_n1163_));
  NOi31      u1135(.An(i), .B(k), .C(j), .Y(men_men_n1164_));
  NA4        u1136(.A(men_men_n1164_), .B(men_men_n1135_), .C(men_men_n357_), .D(men_men_n348_), .Y(men_men_n1165_));
  OAI210     u1137(.A0(men_men_n862_), .A1(men_men_n440_), .B0(men_men_n1165_), .Y(men_men_n1166_));
  NOi31      u1138(.An(m), .B(n), .C(f), .Y(men_men_n1167_));
  NA2        u1139(.A(men_men_n1167_), .B(men_men_n51_), .Y(men_men_n1168_));
  AN2        u1140(.A(e), .B(c), .Y(men_men_n1169_));
  NA2        u1141(.A(men_men_n1169_), .B(a), .Y(men_men_n1170_));
  OAI220     u1142(.A0(men_men_n1170_), .A1(men_men_n1168_), .B0(men_men_n931_), .B1(men_men_n446_), .Y(men_men_n1171_));
  NA2        u1143(.A(men_men_n533_), .B(l), .Y(men_men_n1172_));
  NOi31      u1144(.An(men_men_n908_), .B(men_men_n1090_), .C(men_men_n1172_), .Y(men_men_n1173_));
  NO4        u1145(.A(men_men_n1173_), .B(men_men_n1171_), .C(men_men_n1166_), .D(men_men_n1051_), .Y(men_men_n1174_));
  NO2        u1146(.A(men_men_n292_), .B(a), .Y(men_men_n1175_));
  INV        u1147(.A(men_men_n1096_), .Y(men_men_n1176_));
  NO2        u1148(.A(men_men_n1144_), .B(men_men_n509_), .Y(men_men_n1177_));
  NO2        u1149(.A(men_men_n88_), .B(g), .Y(men_men_n1178_));
  AOI210     u1150(.A0(men_men_n1178_), .A1(men_men_n1177_), .B0(men_men_n1128_), .Y(men_men_n1179_));
  OR2        u1151(.A(men_men_n1179_), .B(men_men_n1126_), .Y(men_men_n1180_));
  NA3        u1152(.A(men_men_n1180_), .B(men_men_n1176_), .C(men_men_n1174_), .Y(men_men_n1181_));
  NO4        u1153(.A(men_men_n1181_), .B(men_men_n1163_), .C(men_men_n864_), .D(men_men_n592_), .Y(men_men_n1182_));
  NA2        u1154(.A(c), .B(b), .Y(men_men_n1183_));
  NO2        u1155(.A(men_men_n732_), .B(men_men_n1183_), .Y(men_men_n1184_));
  OAI210     u1156(.A0(men_men_n906_), .A1(men_men_n879_), .B0(men_men_n433_), .Y(men_men_n1185_));
  OAI210     u1157(.A0(men_men_n1185_), .A1(men_men_n907_), .B0(men_men_n1184_), .Y(men_men_n1186_));
  NAi21      u1158(.An(men_men_n441_), .B(men_men_n1184_), .Y(men_men_n1187_));
  NA3        u1159(.A(men_men_n447_), .B(men_men_n585_), .C(f), .Y(men_men_n1188_));
  OAI210     u1160(.A0(men_men_n575_), .A1(men_men_n39_), .B0(men_men_n1175_), .Y(men_men_n1189_));
  NA3        u1161(.A(men_men_n1189_), .B(men_men_n1188_), .C(men_men_n1187_), .Y(men_men_n1190_));
  NA2        u1162(.A(men_men_n267_), .B(men_men_n122_), .Y(men_men_n1191_));
  OAI210     u1163(.A0(men_men_n1191_), .A1(men_men_n296_), .B0(g), .Y(men_men_n1192_));
  NO2        u1164(.A(f), .B(men_men_n1148_), .Y(men_men_n1193_));
  INV        u1165(.A(men_men_n1193_), .Y(men_men_n1194_));
  AOI210     u1166(.A0(men_men_n1192_), .A1(men_men_n302_), .B0(men_men_n1194_), .Y(men_men_n1195_));
  AOI210     u1167(.A0(men_men_n1195_), .A1(men_men_n116_), .B0(men_men_n1190_), .Y(men_men_n1196_));
  NA2        u1168(.A(men_men_n493_), .B(men_men_n492_), .Y(men_men_n1197_));
  NO2        u1169(.A(men_men_n189_), .B(men_men_n242_), .Y(men_men_n1198_));
  NA2        u1170(.A(men_men_n1198_), .B(m), .Y(men_men_n1199_));
  NA3        u1171(.A(men_men_n963_), .B(men_men_n1172_), .C(men_men_n496_), .Y(men_men_n1200_));
  OAI210     u1172(.A0(men_men_n1200_), .A1(men_men_n323_), .B0(men_men_n494_), .Y(men_men_n1201_));
  AOI210     u1173(.A0(men_men_n1201_), .A1(men_men_n1197_), .B0(men_men_n1199_), .Y(men_men_n1202_));
  NA2        u1174(.A(men_men_n587_), .B(men_men_n428_), .Y(men_men_n1203_));
  NA2        u1175(.A(men_men_n165_), .B(men_men_n33_), .Y(men_men_n1204_));
  AOI210     u1176(.A0(men_men_n1013_), .A1(men_men_n1204_), .B0(men_men_n221_), .Y(men_men_n1205_));
  OAI210     u1177(.A0(men_men_n1205_), .A1(men_men_n467_), .B0(men_men_n1193_), .Y(men_men_n1206_));
  NO2        u1178(.A(men_men_n390_), .B(men_men_n389_), .Y(men_men_n1207_));
  AOI210     u1179(.A0(men_men_n1198_), .A1(men_men_n449_), .B0(men_men_n1007_), .Y(men_men_n1208_));
  NAi41      u1180(.An(men_men_n1207_), .B(men_men_n1208_), .C(men_men_n1206_), .D(men_men_n1203_), .Y(men_men_n1209_));
  NO2        u1181(.A(men_men_n1209_), .B(men_men_n1202_), .Y(men_men_n1210_));
  NA4        u1182(.A(men_men_n1210_), .B(men_men_n1196_), .C(men_men_n1186_), .D(men_men_n1182_), .Y(men00));
  AOI210     u1183(.A0(men_men_n309_), .A1(men_men_n221_), .B0(men_men_n284_), .Y(men_men_n1212_));
  NO2        u1184(.A(men_men_n1212_), .B(men_men_n606_), .Y(men_men_n1213_));
  AOI210     u1185(.A0(men_men_n945_), .A1(men_men_n989_), .B0(men_men_n1166_), .Y(men_men_n1214_));
  NO3        u1186(.A(men_men_n1141_), .B(men_men_n1007_), .C(men_men_n744_), .Y(men_men_n1215_));
  NA3        u1187(.A(men_men_n1215_), .B(men_men_n1214_), .C(men_men_n1053_), .Y(men_men_n1216_));
  NA2        u1188(.A(men_men_n534_), .B(f), .Y(men_men_n1217_));
  NA3        u1189(.A(men_men_n1603_), .B(men_men_n263_), .C(n), .Y(men_men_n1218_));
  AOI210     u1190(.A0(men_men_n1218_), .A1(men_men_n1217_), .B0(men_men_n1100_), .Y(men_men_n1219_));
  NO4        u1191(.A(men_men_n1219_), .B(men_men_n1216_), .C(men_men_n1213_), .D(men_men_n1120_), .Y(men_men_n1220_));
  NA3        u1192(.A(men_men_n175_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1221_));
  NA3        u1193(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1222_));
  NOi31      u1194(.An(n), .B(m), .C(i), .Y(men_men_n1223_));
  NA3        u1195(.A(men_men_n1223_), .B(men_men_n676_), .C(men_men_n51_), .Y(men_men_n1224_));
  OAI210     u1196(.A0(men_men_n1222_), .A1(men_men_n1221_), .B0(men_men_n1224_), .Y(men_men_n1225_));
  INV        u1197(.A(men_men_n605_), .Y(men_men_n1226_));
  NO4        u1198(.A(men_men_n1226_), .B(men_men_n1225_), .C(men_men_n1207_), .D(men_men_n966_), .Y(men_men_n1227_));
  NO4        u1199(.A(men_men_n512_), .B(men_men_n372_), .C(men_men_n1183_), .D(men_men_n59_), .Y(men_men_n1228_));
  NA3        u1200(.A(men_men_n402_), .B(men_men_n228_), .C(g), .Y(men_men_n1229_));
  OA220      u1201(.A0(men_men_n1229_), .A1(men_men_n1222_), .B0(men_men_n403_), .B1(men_men_n139_), .Y(men_men_n1230_));
  NO2        u1202(.A(h), .B(g), .Y(men_men_n1231_));
  NA4        u1203(.A(men_men_n523_), .B(men_men_n490_), .C(men_men_n1231_), .D(men_men_n1089_), .Y(men_men_n1232_));
  OAI220     u1204(.A0(men_men_n553_), .A1(men_men_n628_), .B0(men_men_n93_), .B1(men_men_n92_), .Y(men_men_n1233_));
  AOI220     u1205(.A0(men_men_n1233_), .A1(men_men_n562_), .B0(men_men_n994_), .B1(men_men_n604_), .Y(men_men_n1234_));
  AOI220     u1206(.A0(men_men_n330_), .A1(men_men_n253_), .B0(men_men_n184_), .B1(men_men_n154_), .Y(men_men_n1235_));
  NA4        u1207(.A(men_men_n1235_), .B(men_men_n1234_), .C(men_men_n1232_), .D(men_men_n1230_), .Y(men_men_n1236_));
  NO3        u1208(.A(men_men_n1236_), .B(men_men_n1228_), .C(men_men_n273_), .Y(men_men_n1237_));
  INV        u1209(.A(men_men_n335_), .Y(men_men_n1238_));
  AOI210     u1210(.A0(men_men_n253_), .A1(men_men_n362_), .B0(men_men_n607_), .Y(men_men_n1239_));
  NA3        u1211(.A(men_men_n1239_), .B(men_men_n1238_), .C(men_men_n160_), .Y(men_men_n1240_));
  NO2        u1212(.A(men_men_n244_), .B(men_men_n188_), .Y(men_men_n1241_));
  NA2        u1213(.A(men_men_n1241_), .B(men_men_n447_), .Y(men_men_n1242_));
  NA3        u1214(.A(men_men_n186_), .B(men_men_n115_), .C(g), .Y(men_men_n1243_));
  NOi31      u1215(.An(men_men_n916_), .B(h), .C(men_men_n1243_), .Y(men_men_n1244_));
  NAi31      u1216(.An(men_men_n192_), .B(men_men_n903_), .C(men_men_n490_), .Y(men_men_n1245_));
  NAi31      u1217(.An(men_men_n1244_), .B(men_men_n1245_), .C(men_men_n1242_), .Y(men_men_n1246_));
  NO2        u1218(.A(men_men_n283_), .B(men_men_n74_), .Y(men_men_n1247_));
  NO3        u1219(.A(men_men_n446_), .B(men_men_n875_), .C(n), .Y(men_men_n1248_));
  AOI210     u1220(.A0(men_men_n1248_), .A1(men_men_n1247_), .B0(men_men_n1134_), .Y(men_men_n1249_));
  NAi31      u1221(.An(men_men_n1103_), .B(men_men_n1249_), .C(men_men_n73_), .Y(men_men_n1250_));
  NO4        u1222(.A(men_men_n1250_), .B(men_men_n1246_), .C(men_men_n1240_), .D(men_men_n544_), .Y(men_men_n1251_));
  AN3        u1223(.A(men_men_n1251_), .B(men_men_n1237_), .C(men_men_n1227_), .Y(men_men_n1252_));
  NA2        u1224(.A(men_men_n562_), .B(men_men_n103_), .Y(men_men_n1253_));
  NA3        u1225(.A(men_men_n1167_), .B(men_men_n637_), .C(men_men_n489_), .Y(men_men_n1254_));
  NA4        u1226(.A(men_men_n1254_), .B(men_men_n588_), .C(men_men_n1253_), .D(men_men_n247_), .Y(men_men_n1255_));
  NA2        u1227(.A(men_men_n1160_), .B(men_men_n562_), .Y(men_men_n1256_));
  NA4        u1228(.A(men_men_n676_), .B(men_men_n212_), .C(men_men_n228_), .D(men_men_n169_), .Y(men_men_n1257_));
  NA3        u1229(.A(men_men_n1257_), .B(men_men_n1256_), .C(men_men_n306_), .Y(men_men_n1258_));
  OAI210     u1230(.A0(men_men_n488_), .A1(men_men_n123_), .B0(men_men_n909_), .Y(men_men_n1259_));
  AOI220     u1231(.A0(men_men_n1259_), .A1(men_men_n1200_), .B0(men_men_n587_), .B1(men_men_n428_), .Y(men_men_n1260_));
  OR4        u1232(.A(men_men_n1100_), .B(men_men_n279_), .C(men_men_n229_), .D(e), .Y(men_men_n1261_));
  NO2        u1233(.A(men_men_n224_), .B(men_men_n221_), .Y(men_men_n1262_));
  NA2        u1234(.A(n), .B(e), .Y(men_men_n1263_));
  NO2        u1235(.A(men_men_n1263_), .B(men_men_n152_), .Y(men_men_n1264_));
  AOI220     u1236(.A0(men_men_n1264_), .A1(men_men_n281_), .B0(men_men_n892_), .B1(men_men_n1262_), .Y(men_men_n1265_));
  OAI210     u1237(.A0(men_men_n373_), .A1(men_men_n324_), .B0(men_men_n469_), .Y(men_men_n1266_));
  NA4        u1238(.A(men_men_n1266_), .B(men_men_n1265_), .C(men_men_n1261_), .D(men_men_n1260_), .Y(men_men_n1267_));
  AOI210     u1239(.A0(men_men_n1264_), .A1(men_men_n896_), .B0(men_men_n863_), .Y(men_men_n1268_));
  AOI220     u1240(.A0(men_men_n1003_), .A1(men_men_n604_), .B0(men_men_n676_), .B1(men_men_n250_), .Y(men_men_n1269_));
  NO2        u1241(.A(men_men_n67_), .B(h), .Y(men_men_n1270_));
  NO3        u1242(.A(men_men_n1100_), .B(men_men_n1098_), .C(men_men_n761_), .Y(men_men_n1271_));
  NO2        u1243(.A(men_men_n1132_), .B(men_men_n136_), .Y(men_men_n1272_));
  AN2        u1244(.A(men_men_n1272_), .B(men_men_n1146_), .Y(men_men_n1273_));
  OAI210     u1245(.A0(men_men_n1273_), .A1(men_men_n1271_), .B0(men_men_n1270_), .Y(men_men_n1274_));
  NA4        u1246(.A(men_men_n1274_), .B(men_men_n1269_), .C(men_men_n1268_), .D(men_men_n911_), .Y(men_men_n1275_));
  NO4        u1247(.A(men_men_n1275_), .B(men_men_n1267_), .C(men_men_n1258_), .D(men_men_n1255_), .Y(men_men_n1276_));
  NA2        u1248(.A(men_men_n880_), .B(men_men_n794_), .Y(men_men_n1277_));
  NA4        u1249(.A(men_men_n1277_), .B(men_men_n1276_), .C(men_men_n1252_), .D(men_men_n1220_), .Y(men01));
  AN2        u1250(.A(men_men_n1078_), .B(men_men_n1076_), .Y(men_men_n1279_));
  NO4        u1251(.A(men_men_n843_), .B(men_men_n835_), .C(men_men_n504_), .D(men_men_n290_), .Y(men_men_n1280_));
  NO2        u1252(.A(men_men_n621_), .B(men_men_n299_), .Y(men_men_n1281_));
  NA2        u1253(.A(men_men_n1281_), .B(i), .Y(men_men_n1282_));
  NA3        u1254(.A(men_men_n1282_), .B(men_men_n1280_), .C(men_men_n1279_), .Y(men_men_n1283_));
  NA2        u1255(.A(men_men_n617_), .B(men_men_n91_), .Y(men_men_n1284_));
  NA2        u1256(.A(men_men_n581_), .B(men_men_n278_), .Y(men_men_n1285_));
  NA2        u1257(.A(men_men_n1010_), .B(men_men_n1285_), .Y(men_men_n1286_));
  NA4        u1258(.A(men_men_n1286_), .B(men_men_n1284_), .C(men_men_n959_), .D(men_men_n347_), .Y(men_men_n1287_));
  NA2        u1259(.A(men_men_n739_), .B(men_men_n98_), .Y(men_men_n1288_));
  OAI220     u1260(.A0(men_men_n1288_), .A1(i), .B0(men_men_n369_), .B1(men_men_n294_), .Y(men_men_n1289_));
  OAI210     u1261(.A0(men_men_n821_), .A1(men_men_n634_), .B0(men_men_n1257_), .Y(men_men_n1290_));
  AOI210     u1262(.A0(men_men_n1289_), .A1(men_men_n663_), .B0(men_men_n1290_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n121_), .B(l), .Y(men_men_n1292_));
  OA220      u1264(.A0(men_men_n1292_), .A1(men_men_n614_), .B0(men_men_n688_), .B1(men_men_n387_), .Y(men_men_n1293_));
  NAi41      u1265(.An(men_men_n168_), .B(men_men_n1293_), .C(men_men_n1291_), .D(men_men_n944_), .Y(men_men_n1294_));
  NO3        u1266(.A(men_men_n822_), .B(men_men_n704_), .C(men_men_n537_), .Y(men_men_n1295_));
  NA4        u1267(.A(men_men_n739_), .B(men_men_n98_), .C(men_men_n45_), .D(men_men_n220_), .Y(men_men_n1296_));
  OA220      u1268(.A0(men_men_n1296_), .A1(men_men_n697_), .B0(men_men_n202_), .B1(men_men_n200_), .Y(men_men_n1297_));
  NA3        u1269(.A(men_men_n1297_), .B(men_men_n1295_), .C(men_men_n142_), .Y(men_men_n1298_));
  NO4        u1270(.A(men_men_n1298_), .B(men_men_n1294_), .C(men_men_n1287_), .D(men_men_n1283_), .Y(men_men_n1299_));
  NA2        u1271(.A(men_men_n1229_), .B(men_men_n213_), .Y(men_men_n1300_));
  OAI210     u1272(.A0(men_men_n1300_), .A1(men_men_n312_), .B0(men_men_n557_), .Y(men_men_n1301_));
  NA2        u1273(.A(men_men_n75_), .B(i), .Y(men_men_n1302_));
  AOI210     u1274(.A0(men_men_n620_), .A1(men_men_n614_), .B0(men_men_n1302_), .Y(men_men_n1303_));
  NOi21      u1275(.An(men_men_n589_), .B(men_men_n611_), .Y(men_men_n1304_));
  AOI210     u1276(.A0(men_men_n1304_), .A1(a), .B0(men_men_n1303_), .Y(men_men_n1305_));
  AOI210     u1277(.A0(men_men_n210_), .A1(men_men_n90_), .B0(men_men_n220_), .Y(men_men_n1306_));
  OAI210     u1278(.A0(men_men_n850_), .A1(men_men_n447_), .B0(men_men_n1306_), .Y(men_men_n1307_));
  AN3        u1279(.A(m), .B(l), .C(k), .Y(men_men_n1308_));
  OAI210     u1280(.A0(men_men_n375_), .A1(men_men_n34_), .B0(men_men_n1308_), .Y(men_men_n1309_));
  NA2        u1281(.A(men_men_n209_), .B(men_men_n34_), .Y(men_men_n1310_));
  AO210      u1282(.A0(men_men_n1310_), .A1(men_men_n1309_), .B0(men_men_n346_), .Y(men_men_n1311_));
  NA4        u1283(.A(men_men_n1311_), .B(men_men_n1307_), .C(men_men_n1305_), .D(men_men_n1301_), .Y(men_men_n1312_));
  AOI210     u1284(.A0(men_men_n626_), .A1(men_men_n121_), .B0(men_men_n632_), .Y(men_men_n1313_));
  OAI210     u1285(.A0(men_men_n1292_), .A1(men_men_n623_), .B0(men_men_n1313_), .Y(men_men_n1314_));
  NA2        u1286(.A(men_men_n289_), .B(men_men_n202_), .Y(men_men_n1315_));
  OAI210     u1287(.A0(men_men_n1315_), .A1(men_men_n404_), .B0(men_men_n693_), .Y(men_men_n1316_));
  NO3        u1288(.A(men_men_n862_), .B(men_men_n210_), .C(men_men_n426_), .Y(men_men_n1317_));
  NO2        u1289(.A(men_men_n1317_), .B(men_men_n1007_), .Y(men_men_n1318_));
  OAI210     u1290(.A0(men_men_n1289_), .A1(men_men_n340_), .B0(men_men_n705_), .Y(men_men_n1319_));
  NA4        u1291(.A(men_men_n1319_), .B(men_men_n1318_), .C(men_men_n1316_), .D(men_men_n825_), .Y(men_men_n1320_));
  NO3        u1292(.A(men_men_n1320_), .B(men_men_n1314_), .C(men_men_n1312_), .Y(men_men_n1321_));
  NA3        u1293(.A(men_men_n635_), .B(men_men_n29_), .C(f), .Y(men_men_n1322_));
  NO2        u1294(.A(men_men_n1322_), .B(men_men_n210_), .Y(men_men_n1323_));
  AOI210     u1295(.A0(men_men_n530_), .A1(men_men_n58_), .B0(men_men_n1323_), .Y(men_men_n1324_));
  OR3        u1296(.A(men_men_n1288_), .B(men_men_n636_), .C(i), .Y(men_men_n1325_));
  NA3        u1297(.A(men_men_n775_), .B(men_men_n75_), .C(i), .Y(men_men_n1326_));
  AOI210     u1298(.A0(men_men_n1326_), .A1(men_men_n1296_), .B0(men_men_n1030_), .Y(men_men_n1327_));
  NO2        u1299(.A(men_men_n213_), .B(men_men_n114_), .Y(men_men_n1328_));
  NO3        u1300(.A(men_men_n1328_), .B(men_men_n1327_), .C(men_men_n1225_), .Y(men_men_n1329_));
  NA4        u1301(.A(men_men_n1329_), .B(men_men_n1325_), .C(men_men_n1324_), .D(men_men_n793_), .Y(men_men_n1330_));
  NO2        u1302(.A(men_men_n1017_), .B(men_men_n238_), .Y(men_men_n1331_));
  NO2        u1303(.A(men_men_n1018_), .B(men_men_n582_), .Y(men_men_n1332_));
  OAI210     u1304(.A0(men_men_n1332_), .A1(men_men_n1331_), .B0(men_men_n355_), .Y(men_men_n1333_));
  NA2        u1305(.A(men_men_n599_), .B(men_men_n597_), .Y(men_men_n1334_));
  NO3        u1306(.A(men_men_n80_), .B(men_men_n310_), .C(men_men_n45_), .Y(men_men_n1335_));
  NA2        u1307(.A(men_men_n1335_), .B(men_men_n580_), .Y(men_men_n1336_));
  NA3        u1308(.A(men_men_n1336_), .B(men_men_n1334_), .C(men_men_n699_), .Y(men_men_n1337_));
  OR2        u1309(.A(men_men_n1229_), .B(men_men_n1222_), .Y(men_men_n1338_));
  NO2        u1310(.A(men_men_n387_), .B(men_men_n72_), .Y(men_men_n1339_));
  AOI210     u1311(.A0(men_men_n766_), .A1(men_men_n645_), .B0(men_men_n1339_), .Y(men_men_n1340_));
  NA2        u1312(.A(men_men_n1335_), .B(men_men_n853_), .Y(men_men_n1341_));
  NA4        u1313(.A(men_men_n1341_), .B(men_men_n1340_), .C(men_men_n1338_), .D(men_men_n405_), .Y(men_men_n1342_));
  NOi41      u1314(.An(men_men_n1333_), .B(men_men_n1342_), .C(men_men_n1337_), .D(men_men_n1330_), .Y(men_men_n1343_));
  NO2        u1315(.A(men_men_n135_), .B(men_men_n45_), .Y(men_men_n1344_));
  AO220      u1316(.A0(i), .A1(men_men_n649_), .B0(men_men_n1344_), .B1(men_men_n737_), .Y(men_men_n1345_));
  NA2        u1317(.A(men_men_n1345_), .B(men_men_n355_), .Y(men_men_n1346_));
  NA2        u1318(.A(men_men_n483_), .B(men_men_n139_), .Y(men_men_n1347_));
  NO3        u1319(.A(men_men_n1144_), .B(men_men_n183_), .C(men_men_n88_), .Y(men_men_n1348_));
  AOI220     u1320(.A0(men_men_n1348_), .A1(men_men_n1347_), .B0(men_men_n1335_), .B1(men_men_n1021_), .Y(men_men_n1349_));
  NA2        u1321(.A(men_men_n1349_), .B(men_men_n1346_), .Y(men_men_n1350_));
  NO2        u1322(.A(men_men_n1350_), .B(men_men_n667_), .Y(men_men_n1351_));
  NA4        u1323(.A(men_men_n1351_), .B(men_men_n1343_), .C(men_men_n1321_), .D(men_men_n1299_), .Y(men06));
  NO2        u1324(.A(men_men_n427_), .B(men_men_n586_), .Y(men_men_n1353_));
  NO2        u1325(.A(men_men_n768_), .B(i), .Y(men_men_n1354_));
  OAI210     u1326(.A0(men_men_n1354_), .A1(men_men_n274_), .B0(men_men_n1353_), .Y(men_men_n1355_));
  NO2        u1327(.A(men_men_n231_), .B(men_men_n105_), .Y(men_men_n1356_));
  OAI210     u1328(.A0(men_men_n1356_), .A1(men_men_n1348_), .B0(men_men_n401_), .Y(men_men_n1357_));
  NO3        u1329(.A(men_men_n630_), .B(men_men_n848_), .C(men_men_n633_), .Y(men_men_n1358_));
  OR2        u1330(.A(men_men_n1358_), .B(men_men_n931_), .Y(men_men_n1359_));
  NA4        u1331(.A(men_men_n1359_), .B(men_men_n1357_), .C(men_men_n1355_), .D(men_men_n1333_), .Y(men_men_n1360_));
  NO3        u1332(.A(men_men_n1360_), .B(men_men_n1337_), .C(men_men_n262_), .Y(men_men_n1361_));
  NO2        u1333(.A(men_men_n310_), .B(men_men_n45_), .Y(men_men_n1362_));
  AOI210     u1334(.A0(men_men_n1362_), .A1(men_men_n1022_), .B0(men_men_n1331_), .Y(men_men_n1363_));
  AOI210     u1335(.A0(men_men_n1362_), .A1(men_men_n583_), .B0(men_men_n1345_), .Y(men_men_n1364_));
  AOI210     u1336(.A0(men_men_n1364_), .A1(men_men_n1363_), .B0(men_men_n352_), .Y(men_men_n1365_));
  OAI210     u1337(.A0(men_men_n90_), .A1(men_men_n40_), .B0(men_men_n703_), .Y(men_men_n1366_));
  NA2        u1338(.A(men_men_n1366_), .B(men_men_n671_), .Y(men_men_n1367_));
  NO2        u1339(.A(men_men_n540_), .B(men_men_n180_), .Y(men_men_n1368_));
  NOi21      u1340(.An(men_men_n141_), .B(men_men_n45_), .Y(men_men_n1369_));
  AOI210     u1341(.A0(men_men_n638_), .A1(men_men_n57_), .B0(men_men_n1168_), .Y(men_men_n1370_));
  OAI210     u1342(.A0(men_men_n483_), .A1(men_men_n254_), .B0(men_men_n953_), .Y(men_men_n1371_));
  NO4        u1343(.A(men_men_n1371_), .B(men_men_n1370_), .C(men_men_n1369_), .D(men_men_n1368_), .Y(men_men_n1372_));
  OR2        u1344(.A(men_men_n631_), .B(men_men_n629_), .Y(men_men_n1373_));
  NO2        u1345(.A(men_men_n386_), .B(men_men_n140_), .Y(men_men_n1374_));
  AOI210     u1346(.A0(men_men_n1374_), .A1(men_men_n617_), .B0(men_men_n1373_), .Y(men_men_n1375_));
  NA3        u1347(.A(men_men_n1375_), .B(men_men_n1372_), .C(men_men_n1367_), .Y(men_men_n1376_));
  NO2        u1348(.A(men_men_n784_), .B(men_men_n385_), .Y(men_men_n1377_));
  NO3        u1349(.A(men_men_n705_), .B(men_men_n795_), .C(men_men_n663_), .Y(men_men_n1378_));
  NOi21      u1350(.An(men_men_n1377_), .B(men_men_n1378_), .Y(men_men_n1379_));
  AN2        u1351(.A(men_men_n1003_), .B(men_men_n674_), .Y(men_men_n1380_));
  NO4        u1352(.A(men_men_n1380_), .B(men_men_n1379_), .C(men_men_n1376_), .D(men_men_n1365_), .Y(men_men_n1381_));
  NO2        u1353(.A(men_men_n842_), .B(men_men_n285_), .Y(men_men_n1382_));
  OAI220     u1354(.A0(men_men_n768_), .A1(men_men_n47_), .B0(men_men_n231_), .B1(men_men_n644_), .Y(men_men_n1383_));
  OAI210     u1355(.A0(men_men_n285_), .A1(c), .B0(men_men_n670_), .Y(men_men_n1384_));
  AOI220     u1356(.A0(men_men_n1384_), .A1(men_men_n1383_), .B0(men_men_n1382_), .B1(men_men_n274_), .Y(men_men_n1385_));
  NO3        u1357(.A(men_men_n249_), .B(men_men_n105_), .C(men_men_n292_), .Y(men_men_n1386_));
  OAI220     u1358(.A0(men_men_n730_), .A1(men_men_n254_), .B0(men_men_n536_), .B1(men_men_n540_), .Y(men_men_n1387_));
  OAI210     u1359(.A0(l), .A1(i), .B0(k), .Y(men_men_n1388_));
  NO3        u1360(.A(men_men_n1388_), .B(men_men_n628_), .C(j), .Y(men_men_n1389_));
  NOi21      u1361(.An(men_men_n1389_), .B(men_men_n697_), .Y(men_men_n1390_));
  NO4        u1362(.A(men_men_n1390_), .B(men_men_n1387_), .C(men_men_n1386_), .D(men_men_n1171_), .Y(men_men_n1391_));
  NA4        u1363(.A(men_men_n833_), .B(men_men_n832_), .C(men_men_n457_), .D(men_men_n923_), .Y(men_men_n1392_));
  NAi31      u1364(.An(men_men_n784_), .B(men_men_n1392_), .C(men_men_n209_), .Y(men_men_n1393_));
  NA4        u1365(.A(men_men_n1393_), .B(men_men_n1391_), .C(men_men_n1385_), .D(men_men_n1269_), .Y(men_men_n1394_));
  NOi31      u1366(.An(men_men_n1358_), .B(men_men_n487_), .C(men_men_n413_), .Y(men_men_n1395_));
  OR3        u1367(.A(men_men_n1395_), .B(men_men_n821_), .C(men_men_n567_), .Y(men_men_n1396_));
  OR3        u1368(.A(men_men_n389_), .B(men_men_n231_), .C(men_men_n644_), .Y(men_men_n1397_));
  AOI210     u1369(.A0(men_men_n599_), .A1(men_men_n469_), .B0(men_men_n391_), .Y(men_men_n1398_));
  NA2        u1370(.A(men_men_n1389_), .B(men_men_n829_), .Y(men_men_n1399_));
  NA4        u1371(.A(men_men_n1399_), .B(men_men_n1398_), .C(men_men_n1397_), .D(men_men_n1396_), .Y(men_men_n1400_));
  AOI220     u1372(.A0(men_men_n1377_), .A1(men_men_n794_), .B0(men_men_n1374_), .B1(men_men_n243_), .Y(men_men_n1401_));
  AO220      u1373(.A0(men_men_n1356_), .A1(men_men_n693_), .B0(men_men_n974_), .B1(men_men_n973_), .Y(men_men_n1402_));
  NO3        u1374(.A(men_men_n1402_), .B(men_men_n921_), .C(men_men_n526_), .Y(men_men_n1403_));
  NA3        u1375(.A(men_men_n1403_), .B(men_men_n1401_), .C(men_men_n1341_), .Y(men_men_n1404_));
  NO3        u1376(.A(men_men_n1404_), .B(men_men_n1400_), .C(men_men_n1394_), .Y(men_men_n1405_));
  NA4        u1377(.A(men_men_n1405_), .B(men_men_n1381_), .C(men_men_n1361_), .D(men_men_n1351_), .Y(men07));
  NOi21      u1378(.An(j), .B(k), .Y(men_men_n1407_));
  NA4        u1379(.A(men_men_n186_), .B(men_men_n111_), .C(men_men_n1407_), .D(f), .Y(men_men_n1408_));
  NAi32      u1380(.An(m), .Bn(b), .C(n), .Y(men_men_n1409_));
  NAi21      u1381(.An(f), .B(c), .Y(men_men_n1410_));
  OR2        u1382(.A(e), .B(d), .Y(men_men_n1411_));
  NOi31      u1383(.An(n), .B(m), .C(b), .Y(men_men_n1412_));
  NO3        u1384(.A(men_men_n136_), .B(men_men_n471_), .C(h), .Y(men_men_n1413_));
  INV        u1385(.A(men_men_n1408_), .Y(men_men_n1414_));
  NOi41      u1386(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1415_));
  NA3        u1387(.A(men_men_n1415_), .B(men_men_n913_), .C(men_men_n429_), .Y(men_men_n1416_));
  NOi21      u1388(.An(h), .B(k), .Y(men_men_n1417_));
  NO2        u1389(.A(men_men_n1416_), .B(men_men_n56_), .Y(men_men_n1418_));
  NO3        u1390(.A(men_men_n1106_), .B(men_men_n152_), .C(men_men_n221_), .Y(men_men_n1419_));
  OAI210     u1391(.A0(men_men_n1146_), .A1(men_men_n1419_), .B0(men_men_n228_), .Y(men_men_n1420_));
  NO2        u1392(.A(men_men_n1420_), .B(men_men_n60_), .Y(men_men_n1421_));
  NO2        u1393(.A(k), .B(i), .Y(men_men_n1422_));
  NO2        u1394(.A(men_men_n1118_), .B(men_men_n318_), .Y(men_men_n1423_));
  NA2        u1395(.A(men_men_n568_), .B(men_men_n81_), .Y(men_men_n1424_));
  NA2        u1396(.A(men_men_n1270_), .B(men_men_n300_), .Y(men_men_n1425_));
  NA2        u1397(.A(men_men_n1425_), .B(men_men_n1424_), .Y(men_men_n1426_));
  NO4        u1398(.A(men_men_n1426_), .B(men_men_n1421_), .C(men_men_n1418_), .D(men_men_n1414_), .Y(men_men_n1427_));
  OR2        u1399(.A(h), .B(f), .Y(men_men_n1428_));
  NO3        u1400(.A(n), .B(m), .C(i), .Y(men_men_n1429_));
  OAI210     u1401(.A0(men_men_n1169_), .A1(men_men_n163_), .B0(men_men_n1429_), .Y(men_men_n1430_));
  NO2        u1402(.A(i), .B(g), .Y(men_men_n1431_));
  OR3        u1403(.A(men_men_n1431_), .B(men_men_n1409_), .C(men_men_n71_), .Y(men_men_n1432_));
  OAI220     u1404(.A0(men_men_n1432_), .A1(men_men_n508_), .B0(men_men_n1430_), .B1(men_men_n1428_), .Y(men_men_n1433_));
  NA3        u1405(.A(men_men_n727_), .B(men_men_n713_), .C(men_men_n115_), .Y(men_men_n1434_));
  NA3        u1406(.A(men_men_n1412_), .B(men_men_n1113_), .C(men_men_n701_), .Y(men_men_n1435_));
  AOI210     u1407(.A0(men_men_n1435_), .A1(men_men_n1434_), .B0(men_men_n45_), .Y(men_men_n1436_));
  NA2        u1408(.A(men_men_n1429_), .B(men_men_n669_), .Y(men_men_n1437_));
  NO2        u1409(.A(l), .B(k), .Y(men_men_n1438_));
  NOi41      u1410(.An(men_men_n573_), .B(men_men_n1438_), .C(men_men_n502_), .D(men_men_n463_), .Y(men_men_n1439_));
  NO3        u1411(.A(men_men_n463_), .B(d), .C(c), .Y(men_men_n1440_));
  NO3        u1412(.A(men_men_n1439_), .B(men_men_n1436_), .C(men_men_n1433_), .Y(men_men_n1441_));
  NO2        u1413(.A(men_men_n153_), .B(h), .Y(men_men_n1442_));
  NO2        u1414(.A(g), .B(c), .Y(men_men_n1443_));
  NA3        u1415(.A(men_men_n1443_), .B(men_men_n147_), .C(men_men_n193_), .Y(men_men_n1444_));
  NO2        u1416(.A(men_men_n1444_), .B(men_men_n1600_), .Y(men_men_n1445_));
  NA2        u1417(.A(men_men_n1445_), .B(men_men_n186_), .Y(men_men_n1446_));
  OAI210     u1418(.A0(men_men_n1417_), .A1(men_men_n220_), .B0(men_men_n1127_), .Y(men_men_n1447_));
  NO2        u1419(.A(men_men_n474_), .B(a), .Y(men_men_n1448_));
  NA3        u1420(.A(men_men_n1448_), .B(men_men_n1447_), .C(men_men_n116_), .Y(men_men_n1449_));
  NO2        u1421(.A(i), .B(h), .Y(men_men_n1450_));
  NA2        u1422(.A(men_men_n1450_), .B(men_men_n228_), .Y(men_men_n1451_));
  AOI210     u1423(.A0(men_men_n263_), .A1(men_men_n119_), .B0(men_men_n557_), .Y(men_men_n1452_));
  NO2        u1424(.A(men_men_n1452_), .B(men_men_n1451_), .Y(men_men_n1453_));
  NO2        u1425(.A(men_men_n791_), .B(men_men_n194_), .Y(men_men_n1454_));
  NOi31      u1426(.An(m), .B(n), .C(b), .Y(men_men_n1455_));
  NOi31      u1427(.An(f), .B(d), .C(c), .Y(men_men_n1456_));
  NA2        u1428(.A(men_men_n1456_), .B(men_men_n1455_), .Y(men_men_n1457_));
  INV        u1429(.A(men_men_n1457_), .Y(men_men_n1458_));
  NO3        u1430(.A(men_men_n1458_), .B(men_men_n1454_), .C(men_men_n1453_), .Y(men_men_n1459_));
  NA2        u1431(.A(men_men_n1137_), .B(men_men_n490_), .Y(men_men_n1460_));
  NO4        u1432(.A(men_men_n1460_), .B(men_men_n1113_), .C(men_men_n463_), .D(men_men_n45_), .Y(men_men_n1461_));
  OAI210     u1433(.A0(men_men_n189_), .A1(men_men_n552_), .B0(men_men_n1114_), .Y(men_men_n1462_));
  NO3        u1434(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1463_));
  INV        u1435(.A(men_men_n1462_), .Y(men_men_n1464_));
  NO2        u1436(.A(men_men_n1464_), .B(men_men_n1461_), .Y(men_men_n1465_));
  AN4        u1437(.A(men_men_n1465_), .B(men_men_n1459_), .C(men_men_n1449_), .D(men_men_n1446_), .Y(men_men_n1466_));
  NA2        u1438(.A(men_men_n1412_), .B(men_men_n398_), .Y(men_men_n1467_));
  NO2        u1439(.A(men_men_n1467_), .B(men_men_n1097_), .Y(men_men_n1468_));
  NO2        u1440(.A(men_men_n194_), .B(b), .Y(men_men_n1469_));
  AOI220     u1441(.A0(men_men_n1223_), .A1(men_men_n1469_), .B0(men_men_n1145_), .B1(men_men_n1460_), .Y(men_men_n1470_));
  NO2        u1442(.A(i), .B(men_men_n220_), .Y(men_men_n1471_));
  NA4        u1443(.A(men_men_n1198_), .B(men_men_n1471_), .C(men_men_n106_), .D(m), .Y(men_men_n1472_));
  NAi31      u1444(.An(men_men_n1468_), .B(men_men_n1472_), .C(men_men_n1470_), .Y(men_men_n1473_));
  NO4        u1445(.A(men_men_n136_), .B(g), .C(f), .D(e), .Y(men_men_n1474_));
  NA2        u1446(.A(men_men_n301_), .B(h), .Y(men_men_n1475_));
  NA2        u1447(.A(men_men_n201_), .B(men_men_n100_), .Y(men_men_n1476_));
  OR2        u1448(.A(e), .B(a), .Y(men_men_n1477_));
  NA2        u1449(.A(men_men_n30_), .B(h), .Y(men_men_n1478_));
  NO2        u1450(.A(men_men_n1478_), .B(men_men_n1133_), .Y(men_men_n1479_));
  NOi41      u1451(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1480_));
  NA2        u1452(.A(men_men_n1480_), .B(men_men_n116_), .Y(men_men_n1481_));
  NA2        u1453(.A(men_men_n1415_), .B(men_men_n1438_), .Y(men_men_n1482_));
  NA2        u1454(.A(men_men_n1482_), .B(men_men_n1481_), .Y(men_men_n1483_));
  OR3        u1455(.A(men_men_n567_), .B(men_men_n566_), .C(men_men_n115_), .Y(men_men_n1484_));
  NA2        u1456(.A(men_men_n1167_), .B(men_men_n426_), .Y(men_men_n1485_));
  OAI220     u1457(.A0(men_men_n1485_), .A1(men_men_n456_), .B0(men_men_n1484_), .B1(men_men_n310_), .Y(men_men_n1486_));
  AO210      u1458(.A0(men_men_n1486_), .A1(men_men_n119_), .B0(men_men_n1483_), .Y(men_men_n1487_));
  NO3        u1459(.A(men_men_n1487_), .B(men_men_n1479_), .C(men_men_n1473_), .Y(men_men_n1488_));
  NA4        u1460(.A(men_men_n1488_), .B(men_men_n1466_), .C(men_men_n1441_), .D(men_men_n1427_), .Y(men_men_n1489_));
  NO2        u1461(.A(men_men_n1183_), .B(men_men_n113_), .Y(men_men_n1490_));
  NA2        u1462(.A(men_men_n398_), .B(men_men_n56_), .Y(men_men_n1491_));
  AOI210     u1463(.A0(men_men_n1491_), .A1(men_men_n1106_), .B0(men_men_n1437_), .Y(men_men_n1492_));
  NA2        u1464(.A(men_men_n222_), .B(men_men_n186_), .Y(men_men_n1493_));
  AOI210     u1465(.A0(men_men_n1493_), .A1(men_men_n1243_), .B0(men_men_n1491_), .Y(men_men_n1494_));
  NO2        u1466(.A(men_men_n1138_), .B(men_men_n1133_), .Y(men_men_n1495_));
  NO3        u1467(.A(men_men_n1495_), .B(men_men_n1494_), .C(men_men_n1492_), .Y(men_men_n1496_));
  NA3        u1468(.A(men_men_n1463_), .B(men_men_n1411_), .C(men_men_n1167_), .Y(men_men_n1497_));
  NO3        u1469(.A(men_men_n1133_), .B(men_men_n611_), .C(g), .Y(men_men_n1498_));
  NOi21      u1470(.An(men_men_n1493_), .B(men_men_n1498_), .Y(men_men_n1499_));
  AOI210     u1471(.A0(men_men_n1499_), .A1(men_men_n1476_), .B0(men_men_n1106_), .Y(men_men_n1500_));
  INV        u1472(.A(men_men_n49_), .Y(men_men_n1501_));
  NA2        u1473(.A(men_men_n1501_), .B(men_men_n1231_), .Y(men_men_n1502_));
  INV        u1474(.A(men_men_n1502_), .Y(men_men_n1503_));
  OAI220     u1475(.A0(men_men_n694_), .A1(g), .B0(men_men_n231_), .B1(c), .Y(men_men_n1504_));
  AOI210     u1476(.A0(men_men_n1469_), .A1(men_men_n41_), .B0(men_men_n1504_), .Y(men_men_n1505_));
  NO2        u1477(.A(men_men_n136_), .B(l), .Y(men_men_n1506_));
  NO2        u1478(.A(men_men_n231_), .B(k), .Y(men_men_n1507_));
  OAI210     u1479(.A0(men_men_n1507_), .A1(men_men_n1450_), .B0(men_men_n1506_), .Y(men_men_n1508_));
  OAI220     u1480(.A0(men_men_n1508_), .A1(men_men_n31_), .B0(men_men_n1505_), .B1(men_men_n183_), .Y(men_men_n1509_));
  NO3        u1481(.A(men_men_n1484_), .B(men_men_n490_), .C(men_men_n369_), .Y(men_men_n1510_));
  NO4        u1482(.A(men_men_n1510_), .B(men_men_n1509_), .C(men_men_n1503_), .D(men_men_n1500_), .Y(men_men_n1511_));
  NO3        u1483(.A(men_men_n1148_), .B(men_men_n1411_), .C(men_men_n49_), .Y(men_men_n1512_));
  AOI220     u1484(.A0(men_men_n1512_), .A1(men_men_n221_), .B0(men_men_n1149_), .B1(men_men_n1601_), .Y(men_men_n1513_));
  NO2        u1485(.A(men_men_n1133_), .B(h), .Y(men_men_n1514_));
  NA3        u1486(.A(men_men_n1514_), .B(d), .C(men_men_n1098_), .Y(men_men_n1515_));
  OAI220     u1487(.A0(men_men_n1515_), .A1(c), .B0(men_men_n1513_), .B1(j), .Y(men_men_n1516_));
  NA3        u1488(.A(men_men_n1490_), .B(men_men_n490_), .C(f), .Y(men_men_n1517_));
  NO2        u1489(.A(men_men_n1407_), .B(men_men_n42_), .Y(men_men_n1518_));
  AOI210     u1490(.A0(men_men_n116_), .A1(men_men_n40_), .B0(men_men_n1518_), .Y(men_men_n1519_));
  NO2        u1491(.A(men_men_n1519_), .B(men_men_n1517_), .Y(men_men_n1520_));
  AOI210     u1492(.A0(men_men_n552_), .A1(h), .B0(men_men_n68_), .Y(men_men_n1521_));
  NA2        u1493(.A(men_men_n1521_), .B(men_men_n1448_), .Y(men_men_n1522_));
  NO2        u1494(.A(j), .B(men_men_n182_), .Y(men_men_n1523_));
  NOi21      u1495(.An(d), .B(f), .Y(men_men_n1524_));
  NO3        u1496(.A(men_men_n1456_), .B(men_men_n1524_), .C(men_men_n40_), .Y(men_men_n1525_));
  NA2        u1497(.A(men_men_n1525_), .B(men_men_n1523_), .Y(men_men_n1526_));
  NO2        u1498(.A(men_men_n1411_), .B(f), .Y(men_men_n1527_));
  NA2        u1499(.A(men_men_n1448_), .B(men_men_n1518_), .Y(men_men_n1528_));
  NO2        u1500(.A(men_men_n310_), .B(c), .Y(men_men_n1529_));
  NA2        u1501(.A(men_men_n1529_), .B(men_men_n568_), .Y(men_men_n1530_));
  NA4        u1502(.A(men_men_n1530_), .B(men_men_n1528_), .C(men_men_n1526_), .D(men_men_n1522_), .Y(men_men_n1531_));
  NO3        u1503(.A(men_men_n1531_), .B(men_men_n1520_), .C(men_men_n1516_), .Y(men_men_n1532_));
  NA4        u1504(.A(men_men_n1532_), .B(men_men_n1511_), .C(men_men_n1497_), .D(men_men_n1496_), .Y(men_men_n1533_));
  OAI220     u1505(.A0(men_men_n490_), .A1(men_men_n310_), .B0(men_men_n135_), .B1(men_men_n59_), .Y(men_men_n1534_));
  NA2        u1506(.A(men_men_n1534_), .B(men_men_n1423_), .Y(men_men_n1535_));
  OAI210     u1507(.A0(men_men_n1474_), .A1(men_men_n1412_), .B0(men_men_n928_), .Y(men_men_n1536_));
  OAI220     u1508(.A0(men_men_n1094_), .A1(men_men_n136_), .B0(men_men_n694_), .B1(men_men_n182_), .Y(men_men_n1537_));
  NA2        u1509(.A(men_men_n1537_), .B(men_men_n648_), .Y(men_men_n1538_));
  NA3        u1510(.A(men_men_n1538_), .B(men_men_n1536_), .C(men_men_n1535_), .Y(men_men_n1539_));
  NA2        u1511(.A(men_men_n1443_), .B(men_men_n1524_), .Y(men_men_n1540_));
  NO2        u1512(.A(men_men_n1540_), .B(m), .Y(men_men_n1541_));
  NA3        u1513(.A(men_men_n1146_), .B(men_men_n111_), .C(men_men_n228_), .Y(men_men_n1542_));
  NA2        u1514(.A(men_men_n113_), .B(men_men_n1455_), .Y(men_men_n1543_));
  NA2        u1515(.A(men_men_n1543_), .B(men_men_n1542_), .Y(men_men_n1544_));
  NO3        u1516(.A(men_men_n1544_), .B(men_men_n1541_), .C(men_men_n1539_), .Y(men_men_n1545_));
  NO2        u1517(.A(men_men_n1410_), .B(e), .Y(men_men_n1546_));
  NA2        u1518(.A(men_men_n1546_), .B(men_men_n424_), .Y(men_men_n1547_));
  OR3        u1519(.A(men_men_n1507_), .B(men_men_n1270_), .C(men_men_n136_), .Y(men_men_n1548_));
  NO2        u1520(.A(men_men_n1548_), .B(men_men_n1547_), .Y(men_men_n1549_));
  NO3        u1521(.A(men_men_n1484_), .B(men_men_n369_), .C(a), .Y(men_men_n1550_));
  NO2        u1522(.A(men_men_n1550_), .B(men_men_n1549_), .Y(men_men_n1551_));
  NA2        u1523(.A(men_men_n566_), .B(g), .Y(men_men_n1552_));
  AOI210     u1524(.A0(men_men_n1552_), .A1(men_men_n1440_), .B0(men_men_n1512_), .Y(men_men_n1553_));
  NO2        u1525(.A(men_men_n1477_), .B(f), .Y(men_men_n1554_));
  AOI210     u1526(.A0(men_men_n1178_), .A1(a), .B0(men_men_n1554_), .Y(men_men_n1555_));
  OAI220     u1527(.A0(men_men_n1555_), .A1(men_men_n68_), .B0(men_men_n1553_), .B1(men_men_n220_), .Y(men_men_n1556_));
  NA4        u1528(.A(men_men_n1146_), .B(men_men_n1143_), .C(men_men_n228_), .D(men_men_n67_), .Y(men_men_n1557_));
  NO2        u1529(.A(men_men_n49_), .B(l), .Y(men_men_n1558_));
  INV        u1530(.A(men_men_n508_), .Y(men_men_n1559_));
  OAI210     u1531(.A0(men_men_n1559_), .A1(men_men_n1149_), .B0(men_men_n1558_), .Y(men_men_n1560_));
  NO2        u1532(.A(men_men_n259_), .B(g), .Y(men_men_n1561_));
  NO2        u1533(.A(m), .B(i), .Y(men_men_n1562_));
  AOI220     u1534(.A0(men_men_n1562_), .A1(men_men_n1442_), .B0(men_men_n1125_), .B1(men_men_n1561_), .Y(men_men_n1563_));
  NA3        u1535(.A(men_men_n1563_), .B(men_men_n1560_), .C(men_men_n1557_), .Y(men_men_n1564_));
  NO2        u1536(.A(men_men_n1564_), .B(men_men_n1556_), .Y(men_men_n1565_));
  NA3        u1537(.A(men_men_n1565_), .B(men_men_n1551_), .C(men_men_n1545_), .Y(men_men_n1566_));
  NA3        u1538(.A(men_men_n1009_), .B(men_men_n143_), .C(men_men_n46_), .Y(men_men_n1567_));
  AOI210     u1539(.A0(men_men_n154_), .A1(c), .B0(men_men_n1567_), .Y(men_men_n1568_));
  AO210      u1540(.A0(men_men_n137_), .A1(l), .B0(men_men_n1467_), .Y(men_men_n1569_));
  NO2        u1541(.A(men_men_n71_), .B(c), .Y(men_men_n1570_));
  NO4        u1542(.A(men_men_n1428_), .B(men_men_n192_), .C(men_men_n471_), .D(men_men_n45_), .Y(men_men_n1571_));
  AOI210     u1543(.A0(men_men_n1523_), .A1(men_men_n1570_), .B0(men_men_n1571_), .Y(men_men_n1572_));
  NA2        u1544(.A(men_men_n1572_), .B(men_men_n1569_), .Y(men_men_n1573_));
  NO2        u1545(.A(men_men_n1573_), .B(men_men_n1568_), .Y(men_men_n1574_));
  NO4        u1546(.A(men_men_n231_), .B(men_men_n192_), .C(men_men_n263_), .D(k), .Y(men_men_n1575_));
  NO2        u1547(.A(men_men_n1567_), .B(men_men_n113_), .Y(men_men_n1576_));
  NOi21      u1548(.An(men_men_n1413_), .B(e), .Y(men_men_n1577_));
  NO3        u1549(.A(men_men_n1577_), .B(men_men_n1576_), .C(men_men_n1575_), .Y(men_men_n1578_));
  AO220      u1550(.A0(men_men_n1146_), .A1(men_men_n1132_), .B0(men_men_n1419_), .B1(men_men_n799_), .Y(men_men_n1579_));
  AOI220     u1551(.A0(men_men_n1562_), .A1(men_men_n669_), .B0(men_men_n1110_), .B1(men_men_n166_), .Y(men_men_n1580_));
  NOi31      u1552(.An(men_men_n30_), .B(men_men_n1580_), .C(n), .Y(men_men_n1581_));
  AOI210     u1553(.A0(men_men_n1579_), .A1(men_men_n1223_), .B0(men_men_n1581_), .Y(men_men_n1582_));
  NO2        u1554(.A(men_men_n1517_), .B(men_men_n68_), .Y(men_men_n1583_));
  NO2        u1555(.A(men_men_n1422_), .B(men_men_n121_), .Y(men_men_n1584_));
  NO2        u1556(.A(men_men_n1584_), .B(men_men_n1467_), .Y(men_men_n1585_));
  NO2        u1557(.A(men_men_n1585_), .B(men_men_n1583_), .Y(men_men_n1586_));
  NA4        u1558(.A(men_men_n1586_), .B(men_men_n1582_), .C(men_men_n1578_), .D(men_men_n1574_), .Y(men_men_n1587_));
  OR4        u1559(.A(men_men_n1587_), .B(men_men_n1566_), .C(men_men_n1533_), .D(men_men_n1489_), .Y(men04));
  NOi31      u1560(.An(men_men_n1474_), .B(men_men_n1475_), .C(men_men_n1100_), .Y(men_men_n1589_));
  NA2        u1561(.A(men_men_n1527_), .B(men_men_n867_), .Y(men_men_n1590_));
  NO4        u1562(.A(men_men_n1590_), .B(men_men_n1090_), .C(men_men_n509_), .D(j), .Y(men_men_n1591_));
  OR3        u1563(.A(men_men_n1591_), .B(men_men_n1589_), .C(men_men_n1116_), .Y(men_men_n1592_));
  NO2        u1564(.A(men_men_n92_), .B(k), .Y(men_men_n1593_));
  AOI210     u1565(.A0(men_men_n1593_), .A1(men_men_n1109_), .B0(men_men_n1244_), .Y(men_men_n1594_));
  NA2        u1566(.A(men_men_n1594_), .B(men_men_n1274_), .Y(men_men_n1595_));
  NO4        u1567(.A(men_men_n1595_), .B(men_men_n1592_), .C(men_men_n1123_), .D(men_men_n1105_), .Y(men_men_n1596_));
  NA4        u1568(.A(men_men_n1596_), .B(men_men_n1180_), .C(men_men_n1165_), .D(men_men_n1152_), .Y(men05));
  INV        u1569(.A(l), .Y(men_men_n1600_));
  INV        u1570(.A(n), .Y(men_men_n1601_));
  INV        u1571(.A(men_men_n727_), .Y(men_men_n1602_));
  INV        u1572(.A(m), .Y(men_men_n1603_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule