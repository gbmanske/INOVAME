// Benchmark "top" written by ABC on Fri Jun 21 17:49:29 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n135_,
    new_new_n136_, new_new_n137_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n987_,
    new_new_n988_, new_new_n989_, new_new_n990_, new_new_n991_,
    new_new_n992_, new_new_n993_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g021(.A(new_new_n35_), .Y(men1));
  INV        g022(.A(i_11_), .Y(new_new_n45_));
  NO2        g023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g024(.A(i_2_), .Y(new_new_n47_));
  NA2        g025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g026(.A(i_5_), .Y(new_new_n49_));
  NO2        g027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g041(.A(i_1_), .Y(new_new_n64_));
  INV        g042(.A(new_new_n62_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n51_), .B(i_2_), .Y(new_new_n66_));
  AOI210     g044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n67_));
  NA2        g045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n74_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n75_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  NA2        g055(.A(i_2_), .B(i_8_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_9_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_7_), .Y(new_new_n80_));
  NO2        g058(.A(new_new_n79_), .B(new_new_n64_), .Y(new_new_n81_));
  INV        g059(.A(i_6_), .Y(new_new_n82_));
  NO2        g060(.A(i_2_), .B(i_7_), .Y(new_new_n83_));
  NA2        g061(.A(new_new_n81_), .B(i_7_), .Y(new_new_n84_));
  NAi21      g062(.An(i_6_), .B(i_10_), .Y(new_new_n85_));
  NA2        g063(.A(i_6_), .B(i_9_), .Y(new_new_n86_));
  AOI210     g064(.A0(new_new_n86_), .A1(new_new_n85_), .B0(new_new_n64_), .Y(new_new_n87_));
  NA2        g065(.A(i_2_), .B(i_6_), .Y(new_new_n88_));
  NO3        g066(.A(new_new_n88_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n89_));
  NO2        g067(.A(new_new_n89_), .B(new_new_n87_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n84_), .B0(new_new_n77_), .Y(new_new_n91_));
  AN3        g069(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n92_));
  NAi21      g070(.An(i_6_), .B(i_11_), .Y(new_new_n93_));
  NO2        g071(.A(i_5_), .B(i_8_), .Y(new_new_n94_));
  NOi21      g072(.An(new_new_n94_), .B(new_new_n93_), .Y(new_new_n95_));
  AOI220     g073(.A0(new_new_n95_), .A1(new_new_n63_), .B0(new_new_n92_), .B1(new_new_n32_), .Y(new_new_n96_));
  INV        g074(.A(i_7_), .Y(new_new_n97_));
  NA2        g075(.A(new_new_n47_), .B(new_new_n97_), .Y(new_new_n98_));
  NO2        g076(.A(i_0_), .B(i_5_), .Y(new_new_n99_));
  NO2        g077(.A(new_new_n99_), .B(new_new_n82_), .Y(new_new_n100_));
  NA2        g078(.A(i_12_), .B(i_3_), .Y(new_new_n101_));
  INV        g079(.A(new_new_n101_), .Y(new_new_n102_));
  NA3        g080(.A(new_new_n102_), .B(new_new_n100_), .C(new_new_n98_), .Y(new_new_n103_));
  NAi21      g081(.An(i_7_), .B(i_11_), .Y(new_new_n104_));
  NO3        g082(.A(new_new_n104_), .B(new_new_n85_), .C(new_new_n54_), .Y(new_new_n105_));
  AN2        g083(.A(i_2_), .B(i_10_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(i_7_), .Y(new_new_n107_));
  OR2        g085(.A(new_new_n77_), .B(new_new_n59_), .Y(new_new_n108_));
  NO2        g086(.A(i_8_), .B(new_new_n97_), .Y(new_new_n109_));
  NO3        g087(.A(new_new_n109_), .B(new_new_n108_), .C(new_new_n107_), .Y(new_new_n110_));
  NA2        g088(.A(i_12_), .B(i_7_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n112_), .B(i_0_), .Y(new_new_n113_));
  NA2        g091(.A(i_11_), .B(i_12_), .Y(new_new_n114_));
  OAI210     g092(.A0(new_new_n113_), .A1(new_new_n111_), .B0(new_new_n114_), .Y(new_new_n115_));
  NO2        g093(.A(new_new_n115_), .B(new_new_n110_), .Y(new_new_n116_));
  NAi41      g094(.An(new_new_n105_), .B(new_new_n116_), .C(new_new_n103_), .D(new_new_n96_), .Y(new_new_n117_));
  NOi21      g095(.An(i_1_), .B(i_5_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n118_), .B(i_11_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n120_));
  NA2        g098(.A(i_7_), .B(new_new_n25_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n121_), .B(new_new_n120_), .Y(new_new_n122_));
  NO2        g100(.A(new_new_n122_), .B(new_new_n47_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n86_), .B(new_new_n85_), .Y(new_new_n124_));
  NAi21      g102(.An(i_3_), .B(i_8_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n125_), .B(new_new_n63_), .Y(new_new_n126_));
  NOi31      g104(.An(new_new_n126_), .B(new_new_n124_), .C(new_new_n123_), .Y(new_new_n127_));
  NO2        g105(.A(i_1_), .B(new_new_n82_), .Y(new_new_n128_));
  NO2        g106(.A(i_6_), .B(i_5_), .Y(new_new_n129_));
  NA2        g107(.A(new_new_n129_), .B(i_3_), .Y(new_new_n130_));
  AO210      g108(.A0(new_new_n130_), .A1(new_new_n48_), .B0(new_new_n128_), .Y(new_new_n131_));
  OAI220     g109(.A0(new_new_n131_), .A1(new_new_n104_), .B0(new_new_n127_), .B1(new_new_n119_), .Y(new_new_n132_));
  NO3        g110(.A(new_new_n132_), .B(new_new_n117_), .C(new_new_n91_), .Y(new_new_n133_));
  NA3        g111(.A(new_new_n133_), .B(new_new_n76_), .C(new_new_n57_), .Y(men2));
  NO2        g112(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n135_));
  NA2        g113(.A(i_6_), .B(new_new_n25_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(new_new_n135_), .Y(new_new_n137_));
  NA4        g115(.A(new_new_n137_), .B(new_new_n74_), .C(new_new_n66_), .D(new_new_n30_), .Y(men0));
  AN2        g116(.A(i_8_), .B(i_7_), .Y(new_new_n139_));
  NA2        g117(.A(new_new_n139_), .B(i_6_), .Y(new_new_n140_));
  NO2        g118(.A(i_12_), .B(i_13_), .Y(new_new_n141_));
  NAi21      g119(.An(i_5_), .B(i_11_), .Y(new_new_n142_));
  NOi21      g120(.An(new_new_n141_), .B(new_new_n142_), .Y(new_new_n143_));
  NO2        g121(.A(i_0_), .B(i_1_), .Y(new_new_n144_));
  NA2        g122(.A(i_2_), .B(i_3_), .Y(new_new_n145_));
  NO2        g123(.A(new_new_n145_), .B(i_4_), .Y(new_new_n146_));
  NA3        g124(.A(new_new_n146_), .B(new_new_n144_), .C(new_new_n143_), .Y(new_new_n147_));
  OR2        g125(.A(new_new_n147_), .B(new_new_n25_), .Y(new_new_n148_));
  AN2        g126(.A(new_new_n141_), .B(new_new_n79_), .Y(new_new_n149_));
  NA2        g127(.A(i_1_), .B(i_5_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n70_), .B(new_new_n47_), .Y(new_new_n151_));
  NA2        g129(.A(new_new_n151_), .B(new_new_n36_), .Y(new_new_n152_));
  NO3        g130(.A(new_new_n152_), .B(new_new_n150_), .C(i_13_), .Y(new_new_n153_));
  OR2        g131(.A(i_0_), .B(i_1_), .Y(new_new_n154_));
  NO3        g132(.A(new_new_n154_), .B(new_new_n77_), .C(i_13_), .Y(new_new_n155_));
  NAi32      g133(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n156_));
  NAi21      g134(.An(new_new_n156_), .B(new_new_n155_), .Y(new_new_n157_));
  NOi21      g135(.An(i_4_), .B(i_10_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n40_), .Y(new_new_n159_));
  NO2        g137(.A(i_3_), .B(i_5_), .Y(new_new_n160_));
  NO3        g138(.A(new_new_n70_), .B(i_2_), .C(i_1_), .Y(new_new_n161_));
  NA2        g139(.A(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  OAI210     g140(.A0(new_new_n162_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n163_), .B(new_new_n153_), .Y(new_new_n164_));
  AOI210     g142(.A0(new_new_n164_), .A1(new_new_n148_), .B0(new_new_n140_), .Y(new_new_n165_));
  NA2        g143(.A(i_3_), .B(new_new_n49_), .Y(new_new_n166_));
  NOi21      g144(.An(i_4_), .B(i_9_), .Y(new_new_n167_));
  NOi21      g145(.An(i_11_), .B(i_13_), .Y(new_new_n168_));
  NA2        g146(.A(new_new_n168_), .B(new_new_n167_), .Y(new_new_n169_));
  NO2        g147(.A(i_4_), .B(i_5_), .Y(new_new_n170_));
  NAi21      g148(.An(i_12_), .B(i_11_), .Y(new_new_n171_));
  NO2        g149(.A(new_new_n171_), .B(i_13_), .Y(new_new_n172_));
  NA3        g150(.A(new_new_n172_), .B(new_new_n170_), .C(new_new_n79_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n173_), .B(new_new_n989_), .Y(new_new_n174_));
  NO2        g152(.A(new_new_n70_), .B(new_new_n64_), .Y(new_new_n175_));
  NA2        g153(.A(new_new_n175_), .B(new_new_n47_), .Y(new_new_n176_));
  NA2        g154(.A(new_new_n36_), .B(i_5_), .Y(new_new_n177_));
  NAi31      g155(.An(new_new_n177_), .B(new_new_n149_), .C(i_11_), .Y(new_new_n178_));
  NA2        g156(.A(i_3_), .B(i_5_), .Y(new_new_n179_));
  AOI210     g157(.A0(new_new_n169_), .A1(new_new_n178_), .B0(new_new_n176_), .Y(new_new_n180_));
  NO2        g158(.A(new_new_n70_), .B(i_5_), .Y(new_new_n181_));
  NO2        g159(.A(i_13_), .B(i_10_), .Y(new_new_n182_));
  NA3        g160(.A(new_new_n182_), .B(new_new_n181_), .C(new_new_n45_), .Y(new_new_n183_));
  NO2        g161(.A(i_2_), .B(i_1_), .Y(new_new_n184_));
  NA2        g162(.A(new_new_n184_), .B(i_3_), .Y(new_new_n185_));
  NAi21      g163(.An(i_4_), .B(i_12_), .Y(new_new_n186_));
  NO4        g164(.A(new_new_n186_), .B(new_new_n185_), .C(new_new_n183_), .D(new_new_n25_), .Y(new_new_n187_));
  NO3        g165(.A(new_new_n187_), .B(new_new_n180_), .C(new_new_n174_), .Y(new_new_n188_));
  INV        g166(.A(i_8_), .Y(new_new_n189_));
  NA2        g167(.A(i_8_), .B(i_6_), .Y(new_new_n190_));
  NO3        g168(.A(i_3_), .B(new_new_n82_), .C(new_new_n49_), .Y(new_new_n191_));
  NA2        g169(.A(new_new_n191_), .B(new_new_n109_), .Y(new_new_n192_));
  NO3        g170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n193_));
  NA3        g171(.A(new_new_n193_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n194_));
  NO3        g172(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n195_));
  NA2        g173(.A(new_new_n92_), .B(new_new_n195_), .Y(new_new_n196_));
  AOI210     g174(.A0(new_new_n196_), .A1(new_new_n194_), .B0(new_new_n192_), .Y(new_new_n197_));
  NO2        g175(.A(i_3_), .B(i_8_), .Y(new_new_n198_));
  NO3        g176(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n199_));
  NA3        g177(.A(new_new_n199_), .B(new_new_n198_), .C(new_new_n40_), .Y(new_new_n200_));
  NO2        g178(.A(i_13_), .B(i_9_), .Y(new_new_n201_));
  NA3        g179(.A(new_new_n201_), .B(i_6_), .C(new_new_n189_), .Y(new_new_n202_));
  NAi21      g180(.An(i_12_), .B(i_3_), .Y(new_new_n203_));
  OR2        g181(.A(new_new_n203_), .B(new_new_n202_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n45_), .B(i_5_), .Y(new_new_n205_));
  NO3        g183(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n206_));
  INV        g184(.A(new_new_n206_), .Y(new_new_n207_));
  OAI220     g185(.A0(new_new_n207_), .A1(new_new_n204_), .B0(new_new_n59_), .B1(new_new_n200_), .Y(new_new_n208_));
  AOI210     g186(.A0(new_new_n208_), .A1(i_7_), .B0(new_new_n197_), .Y(new_new_n209_));
  OAI220     g187(.A0(new_new_n209_), .A1(i_4_), .B0(new_new_n190_), .B1(new_new_n188_), .Y(new_new_n210_));
  NAi21      g188(.An(i_12_), .B(i_7_), .Y(new_new_n211_));
  NA3        g189(.A(i_13_), .B(new_new_n189_), .C(i_10_), .Y(new_new_n212_));
  NO2        g190(.A(new_new_n212_), .B(new_new_n211_), .Y(new_new_n213_));
  NA2        g191(.A(i_0_), .B(i_5_), .Y(new_new_n214_));
  NA2        g192(.A(new_new_n214_), .B(new_new_n100_), .Y(new_new_n215_));
  OAI220     g193(.A0(new_new_n215_), .A1(new_new_n185_), .B0(new_new_n176_), .B1(new_new_n130_), .Y(new_new_n216_));
  NAi31      g194(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n217_));
  NO2        g195(.A(new_new_n36_), .B(i_13_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n70_), .B(new_new_n26_), .Y(new_new_n219_));
  NO2        g197(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n220_));
  NA3        g198(.A(new_new_n220_), .B(new_new_n219_), .C(new_new_n218_), .Y(new_new_n221_));
  INV        g199(.A(i_13_), .Y(new_new_n222_));
  NO2        g200(.A(i_12_), .B(new_new_n222_), .Y(new_new_n223_));
  NA3        g201(.A(new_new_n223_), .B(new_new_n193_), .C(new_new_n191_), .Y(new_new_n224_));
  OAI210     g202(.A0(new_new_n221_), .A1(new_new_n217_), .B0(new_new_n224_), .Y(new_new_n225_));
  AOI220     g203(.A0(new_new_n225_), .A1(new_new_n139_), .B0(new_new_n216_), .B1(new_new_n213_), .Y(new_new_n226_));
  NO2        g204(.A(i_12_), .B(new_new_n37_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n179_), .B(i_4_), .Y(new_new_n228_));
  NA2        g206(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n229_));
  OR2        g207(.A(i_8_), .B(i_7_), .Y(new_new_n230_));
  NO2        g208(.A(new_new_n230_), .B(new_new_n82_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n54_), .B(i_1_), .Y(new_new_n232_));
  INV        g210(.A(i_12_), .Y(new_new_n233_));
  NO3        g211(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n234_));
  NA2        g212(.A(i_2_), .B(i_1_), .Y(new_new_n235_));
  NO3        g213(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n236_));
  NAi21      g214(.An(i_4_), .B(i_3_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n237_), .B(new_new_n72_), .Y(new_new_n238_));
  NO2        g216(.A(i_0_), .B(i_6_), .Y(new_new_n239_));
  NOi41      g217(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n240_));
  NA2        g218(.A(new_new_n240_), .B(new_new_n239_), .Y(new_new_n241_));
  NO2        g219(.A(new_new_n235_), .B(new_new_n179_), .Y(new_new_n242_));
  NAi21      g220(.An(new_new_n241_), .B(new_new_n242_), .Y(new_new_n243_));
  NO2        g221(.A(i_11_), .B(new_new_n222_), .Y(new_new_n244_));
  NAi21      g222(.An(i_3_), .B(i_7_), .Y(new_new_n245_));
  NO2        g223(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n246_));
  NO2        g224(.A(i_12_), .B(i_3_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n70_), .B(i_5_), .Y(new_new_n248_));
  NA3        g226(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n249_));
  INV        g227(.A(new_new_n140_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n233_), .B(i_13_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n251_), .B(new_new_n72_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n252_), .B(new_new_n250_), .Y(new_new_n253_));
  NO2        g231(.A(new_new_n230_), .B(new_new_n37_), .Y(new_new_n254_));
  NA2        g232(.A(i_12_), .B(i_6_), .Y(new_new_n255_));
  OR2        g233(.A(i_13_), .B(i_9_), .Y(new_new_n256_));
  NO3        g234(.A(new_new_n256_), .B(new_new_n255_), .C(new_new_n49_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n237_), .B(i_2_), .Y(new_new_n258_));
  NA3        g236(.A(new_new_n258_), .B(new_new_n257_), .C(new_new_n45_), .Y(new_new_n259_));
  NA2        g237(.A(new_new_n244_), .B(i_9_), .Y(new_new_n260_));
  OAI210     g238(.A0(new_new_n70_), .A1(new_new_n260_), .B0(new_new_n259_), .Y(new_new_n261_));
  NO3        g239(.A(i_11_), .B(new_new_n222_), .C(new_new_n25_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n245_), .B(i_8_), .Y(new_new_n263_));
  NO2        g241(.A(i_6_), .B(new_new_n49_), .Y(new_new_n264_));
  NA3        g242(.A(new_new_n264_), .B(new_new_n263_), .C(new_new_n262_), .Y(new_new_n265_));
  NO3        g243(.A(new_new_n26_), .B(new_new_n82_), .C(i_5_), .Y(new_new_n266_));
  NA3        g244(.A(new_new_n266_), .B(new_new_n254_), .C(new_new_n223_), .Y(new_new_n267_));
  AOI210     g245(.A0(new_new_n267_), .A1(new_new_n265_), .B0(i_1_), .Y(new_new_n268_));
  AOI210     g246(.A0(new_new_n261_), .A1(new_new_n254_), .B0(new_new_n268_), .Y(new_new_n269_));
  NA4        g247(.A(new_new_n269_), .B(new_new_n253_), .C(new_new_n243_), .D(new_new_n226_), .Y(new_new_n270_));
  NO3        g248(.A(i_12_), .B(new_new_n222_), .C(new_new_n37_), .Y(new_new_n271_));
  INV        g249(.A(new_new_n271_), .Y(new_new_n272_));
  NA2        g250(.A(i_8_), .B(new_new_n97_), .Y(new_new_n273_));
  NO3        g251(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n274_));
  AOI220     g252(.A0(new_new_n274_), .A1(new_new_n191_), .B0(new_new_n160_), .B1(new_new_n232_), .Y(new_new_n275_));
  NO2        g253(.A(new_new_n275_), .B(new_new_n273_), .Y(new_new_n276_));
  NO2        g254(.A(new_new_n235_), .B(i_0_), .Y(new_new_n277_));
  AOI220     g255(.A0(new_new_n277_), .A1(i_8_), .B0(i_1_), .B1(new_new_n139_), .Y(new_new_n278_));
  NA2        g256(.A(new_new_n264_), .B(new_new_n26_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n279_), .B(new_new_n278_), .Y(new_new_n280_));
  NA2        g258(.A(i_0_), .B(i_1_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n281_), .B(i_2_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n60_), .B(i_6_), .Y(new_new_n283_));
  NA3        g261(.A(new_new_n283_), .B(new_new_n282_), .C(new_new_n160_), .Y(new_new_n284_));
  OAI210     g262(.A0(new_new_n162_), .A1(new_new_n140_), .B0(new_new_n284_), .Y(new_new_n285_));
  NO3        g263(.A(new_new_n285_), .B(new_new_n280_), .C(new_new_n276_), .Y(new_new_n286_));
  NO2        g264(.A(i_3_), .B(i_10_), .Y(new_new_n287_));
  NA3        g265(.A(new_new_n287_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n288_));
  NO2        g266(.A(i_2_), .B(new_new_n97_), .Y(new_new_n289_));
  NA2        g267(.A(i_1_), .B(new_new_n36_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n290_), .B(i_8_), .Y(new_new_n291_));
  NA2        g269(.A(new_new_n291_), .B(new_new_n289_), .Y(new_new_n292_));
  AN2        g270(.A(i_3_), .B(i_10_), .Y(new_new_n293_));
  NA3        g271(.A(new_new_n293_), .B(new_new_n172_), .C(new_new_n170_), .Y(new_new_n294_));
  NO2        g272(.A(i_5_), .B(new_new_n37_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n296_));
  OR2        g274(.A(new_new_n292_), .B(new_new_n288_), .Y(new_new_n297_));
  OAI220     g275(.A0(new_new_n297_), .A1(i_6_), .B0(new_new_n286_), .B1(new_new_n272_), .Y(new_new_n298_));
  NO4        g276(.A(new_new_n298_), .B(new_new_n270_), .C(new_new_n210_), .D(new_new_n165_), .Y(new_new_n299_));
  NO3        g277(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n300_));
  NO3        g278(.A(i_6_), .B(new_new_n189_), .C(i_7_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n189_), .B(new_new_n166_), .Y(new_new_n302_));
  NO2        g280(.A(i_2_), .B(i_3_), .Y(new_new_n303_));
  OR2        g281(.A(i_0_), .B(i_5_), .Y(new_new_n304_));
  NA2        g282(.A(new_new_n214_), .B(new_new_n304_), .Y(new_new_n305_));
  NA4        g283(.A(new_new_n305_), .B(new_new_n231_), .C(new_new_n303_), .D(i_1_), .Y(new_new_n306_));
  NA3        g284(.A(new_new_n277_), .B(new_new_n160_), .C(new_new_n109_), .Y(new_new_n307_));
  NAi21      g285(.An(i_8_), .B(i_7_), .Y(new_new_n308_));
  NO2        g286(.A(new_new_n308_), .B(i_6_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n154_), .B(new_new_n47_), .Y(new_new_n310_));
  NA3        g288(.A(new_new_n310_), .B(new_new_n309_), .C(new_new_n160_), .Y(new_new_n311_));
  NA3        g289(.A(new_new_n311_), .B(new_new_n307_), .C(new_new_n306_), .Y(new_new_n312_));
  OAI210     g290(.A0(new_new_n312_), .A1(new_new_n302_), .B0(i_4_), .Y(new_new_n313_));
  NO2        g291(.A(i_12_), .B(i_10_), .Y(new_new_n314_));
  NOi21      g292(.An(i_5_), .B(i_0_), .Y(new_new_n315_));
  NO2        g293(.A(new_new_n290_), .B(new_new_n125_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n316_), .B(new_new_n314_), .Y(new_new_n317_));
  NO2        g295(.A(i_6_), .B(i_8_), .Y(new_new_n318_));
  NOi21      g296(.An(i_0_), .B(i_2_), .Y(new_new_n319_));
  AN2        g297(.A(new_new_n319_), .B(new_new_n318_), .Y(new_new_n320_));
  NO2        g298(.A(i_1_), .B(i_7_), .Y(new_new_n321_));
  AO220      g299(.A0(new_new_n321_), .A1(new_new_n320_), .B0(new_new_n309_), .B1(new_new_n232_), .Y(new_new_n322_));
  NA2        g300(.A(new_new_n322_), .B(new_new_n42_), .Y(new_new_n323_));
  NA3        g301(.A(new_new_n323_), .B(new_new_n317_), .C(new_new_n313_), .Y(new_new_n324_));
  NO3        g302(.A(new_new_n230_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n325_));
  NO3        g303(.A(new_new_n308_), .B(i_2_), .C(i_1_), .Y(new_new_n326_));
  OAI210     g304(.A0(new_new_n326_), .A1(new_new_n325_), .B0(i_6_), .Y(new_new_n327_));
  NA2        g305(.A(i_1_), .B(new_new_n289_), .Y(new_new_n328_));
  AOI210     g306(.A0(new_new_n328_), .A1(new_new_n327_), .B0(new_new_n305_), .Y(new_new_n329_));
  NOi21      g307(.An(new_new_n150_), .B(new_new_n100_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n330_), .B(new_new_n121_), .Y(new_new_n331_));
  OAI210     g309(.A0(new_new_n331_), .A1(new_new_n329_), .B0(i_3_), .Y(new_new_n332_));
  INV        g310(.A(new_new_n80_), .Y(new_new_n333_));
  NO2        g311(.A(new_new_n281_), .B(new_new_n78_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n334_), .B(new_new_n129_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n88_), .B(new_new_n189_), .Y(new_new_n336_));
  NA2        g314(.A(new_new_n336_), .B(new_new_n64_), .Y(new_new_n337_));
  AOI210     g315(.A0(new_new_n337_), .A1(new_new_n335_), .B0(new_new_n333_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n189_), .B(i_9_), .Y(new_new_n339_));
  NA2        g317(.A(new_new_n339_), .B(i_6_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n338_), .B(new_new_n280_), .Y(new_new_n341_));
  AOI210     g319(.A0(new_new_n341_), .A1(new_new_n332_), .B0(new_new_n159_), .Y(new_new_n342_));
  AOI210     g320(.A0(new_new_n324_), .A1(new_new_n300_), .B0(new_new_n342_), .Y(new_new_n343_));
  NOi32      g321(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n344_));
  INV        g322(.A(new_new_n344_), .Y(new_new_n345_));
  NAi21      g323(.An(i_0_), .B(i_6_), .Y(new_new_n346_));
  NAi21      g324(.An(i_1_), .B(i_5_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n347_), .B(new_new_n346_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n348_), .B(new_new_n25_), .Y(new_new_n349_));
  OAI210     g327(.A0(new_new_n349_), .A1(new_new_n156_), .B0(new_new_n241_), .Y(new_new_n350_));
  NAi41      g328(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n351_));
  AOI210     g329(.A0(new_new_n351_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n352_));
  NOi32      g330(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n353_));
  NO2        g331(.A(i_1_), .B(new_new_n97_), .Y(new_new_n354_));
  NAi21      g332(.An(i_3_), .B(i_4_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n355_), .B(i_9_), .Y(new_new_n356_));
  AN2        g334(.A(i_6_), .B(i_7_), .Y(new_new_n357_));
  OAI210     g335(.A0(new_new_n357_), .A1(new_new_n354_), .B0(new_new_n356_), .Y(new_new_n358_));
  NA2        g336(.A(i_2_), .B(i_7_), .Y(new_new_n359_));
  NO2        g337(.A(new_new_n355_), .B(i_10_), .Y(new_new_n360_));
  NA3        g338(.A(new_new_n360_), .B(new_new_n359_), .C(new_new_n239_), .Y(new_new_n361_));
  AOI210     g339(.A0(new_new_n361_), .A1(new_new_n358_), .B0(new_new_n181_), .Y(new_new_n362_));
  AOI210     g340(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n363_));
  OAI210     g341(.A0(new_new_n363_), .A1(new_new_n184_), .B0(new_new_n360_), .Y(new_new_n364_));
  AOI220     g342(.A0(new_new_n360_), .A1(new_new_n321_), .B0(new_new_n234_), .B1(new_new_n184_), .Y(new_new_n365_));
  AOI210     g343(.A0(new_new_n365_), .A1(new_new_n364_), .B0(i_5_), .Y(new_new_n366_));
  NO4        g344(.A(new_new_n366_), .B(new_new_n362_), .C(new_new_n352_), .D(new_new_n350_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n367_), .B(new_new_n345_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n369_));
  AN2        g347(.A(i_12_), .B(i_5_), .Y(new_new_n370_));
  NO2        g348(.A(i_4_), .B(new_new_n26_), .Y(new_new_n371_));
  NA2        g349(.A(new_new_n371_), .B(new_new_n370_), .Y(new_new_n372_));
  NO2        g350(.A(i_11_), .B(i_6_), .Y(new_new_n373_));
  NA3        g351(.A(new_new_n373_), .B(new_new_n310_), .C(new_new_n222_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n374_), .B(new_new_n372_), .Y(new_new_n375_));
  NO2        g353(.A(new_new_n237_), .B(i_5_), .Y(new_new_n376_));
  NO2        g354(.A(i_5_), .B(i_10_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n376_), .B(new_new_n193_), .Y(new_new_n378_));
  NO2        g356(.A(i_12_), .B(new_new_n378_), .Y(new_new_n379_));
  OAI210     g357(.A0(new_new_n379_), .A1(new_new_n375_), .B0(new_new_n369_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n381_));
  INV        g359(.A(new_new_n147_), .Y(new_new_n382_));
  OAI210     g360(.A0(new_new_n382_), .A1(new_new_n375_), .B0(new_new_n381_), .Y(new_new_n383_));
  NO3        g361(.A(new_new_n82_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n384_));
  NO2        g362(.A(i_11_), .B(i_12_), .Y(new_new_n385_));
  NA2        g363(.A(new_new_n377_), .B(new_new_n233_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n109_), .B(new_new_n42_), .Y(new_new_n387_));
  NO2        g365(.A(new_new_n387_), .B(new_new_n217_), .Y(new_new_n388_));
  NAi21      g366(.An(i_13_), .B(i_0_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n389_), .B(new_new_n235_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n388_), .B(new_new_n390_), .Y(new_new_n391_));
  NA3        g369(.A(new_new_n391_), .B(new_new_n383_), .C(new_new_n380_), .Y(new_new_n392_));
  NO3        g370(.A(i_1_), .B(i_12_), .C(new_new_n82_), .Y(new_new_n393_));
  NO2        g371(.A(i_0_), .B(i_11_), .Y(new_new_n394_));
  INV        g372(.A(i_5_), .Y(new_new_n395_));
  AN2        g373(.A(i_1_), .B(i_6_), .Y(new_new_n396_));
  NOi21      g374(.An(i_2_), .B(i_12_), .Y(new_new_n397_));
  NA2        g375(.A(new_new_n397_), .B(new_new_n396_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n395_), .Y(new_new_n399_));
  NA2        g377(.A(new_new_n139_), .B(i_9_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n400_), .B(i_4_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n399_), .B(new_new_n401_), .Y(new_new_n402_));
  NAi21      g380(.An(i_9_), .B(i_4_), .Y(new_new_n403_));
  OR2        g381(.A(i_13_), .B(i_10_), .Y(new_new_n404_));
  NO3        g382(.A(new_new_n404_), .B(new_new_n114_), .C(new_new_n403_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n169_), .B(new_new_n120_), .Y(new_new_n406_));
  BUFFER     g384(.A(new_new_n212_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n97_), .B(new_new_n25_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n271_), .B(new_new_n408_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n264_), .B(new_new_n206_), .Y(new_new_n410_));
  OAI220     g388(.A0(new_new_n410_), .A1(new_new_n407_), .B0(new_new_n409_), .B1(new_new_n330_), .Y(new_new_n411_));
  INV        g389(.A(new_new_n411_), .Y(new_new_n412_));
  AOI210     g390(.A0(new_new_n412_), .A1(new_new_n402_), .B0(new_new_n26_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n307_), .B(new_new_n306_), .Y(new_new_n414_));
  AOI220     g392(.A0(new_new_n283_), .A1(new_new_n274_), .B0(new_new_n277_), .B1(i_6_), .Y(new_new_n415_));
  NO2        g393(.A(new_new_n415_), .B(new_new_n166_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n179_), .B(new_new_n82_), .Y(new_new_n417_));
  AOI220     g395(.A0(new_new_n417_), .A1(new_new_n282_), .B0(new_new_n266_), .B1(new_new_n206_), .Y(new_new_n418_));
  NO2        g396(.A(new_new_n418_), .B(new_new_n273_), .Y(new_new_n419_));
  NO3        g397(.A(new_new_n419_), .B(new_new_n416_), .C(new_new_n414_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n191_), .B(new_new_n92_), .Y(new_new_n421_));
  NA3        g399(.A(new_new_n310_), .B(new_new_n160_), .C(new_new_n82_), .Y(new_new_n422_));
  AOI210     g400(.A0(new_new_n422_), .A1(new_new_n421_), .B0(new_new_n308_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n283_), .B(new_new_n232_), .Y(new_new_n424_));
  NO2        g402(.A(new_new_n424_), .B(new_new_n179_), .Y(new_new_n425_));
  NA3        g403(.A(new_new_n321_), .B(new_new_n320_), .C(i_5_), .Y(new_new_n426_));
  INV        g404(.A(new_new_n301_), .Y(new_new_n427_));
  OAI210     g405(.A0(new_new_n427_), .A1(new_new_n185_), .B0(new_new_n426_), .Y(new_new_n428_));
  NO3        g406(.A(new_new_n428_), .B(new_new_n425_), .C(new_new_n423_), .Y(new_new_n429_));
  AOI210     g407(.A0(new_new_n429_), .A1(new_new_n420_), .B0(new_new_n260_), .Y(new_new_n430_));
  NO4        g408(.A(new_new_n430_), .B(new_new_n413_), .C(new_new_n392_), .D(new_new_n368_), .Y(new_new_n431_));
  NO2        g409(.A(new_new_n64_), .B(i_4_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n70_), .B(i_13_), .Y(new_new_n433_));
  NO2        g411(.A(i_10_), .B(i_9_), .Y(new_new_n434_));
  NAi21      g412(.An(i_12_), .B(i_8_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n296_), .B(i_0_), .Y(new_new_n436_));
  NO3        g414(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n255_), .B(new_new_n93_), .Y(new_new_n438_));
  NA2        g416(.A(i_8_), .B(i_9_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n244_), .B(new_new_n295_), .Y(new_new_n440_));
  NO3        g418(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n441_));
  INV        g419(.A(new_new_n441_), .Y(new_new_n442_));
  NA3        g420(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n443_));
  NA4        g421(.A(new_new_n142_), .B(new_new_n112_), .C(new_new_n77_), .D(new_new_n23_), .Y(new_new_n444_));
  OAI220     g422(.A0(new_new_n444_), .A1(new_new_n443_), .B0(new_new_n442_), .B1(new_new_n440_), .Y(new_new_n445_));
  INV        g423(.A(new_new_n445_), .Y(new_new_n446_));
  OA210      g424(.A0(new_new_n340_), .A1(new_new_n97_), .B0(new_new_n284_), .Y(new_new_n447_));
  OA220      g425(.A0(new_new_n447_), .A1(new_new_n159_), .B0(new_new_n202_), .B1(new_new_n229_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n92_), .B(i_13_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n417_), .B(new_new_n369_), .Y(new_new_n450_));
  NO2        g428(.A(i_2_), .B(i_13_), .Y(new_new_n451_));
  NO2        g429(.A(new_new_n450_), .B(new_new_n449_), .Y(new_new_n452_));
  NO3        g430(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n453_));
  NO2        g431(.A(i_6_), .B(i_7_), .Y(new_new_n454_));
  NA2        g432(.A(new_new_n454_), .B(new_new_n453_), .Y(new_new_n455_));
  NO2        g433(.A(i_11_), .B(i_1_), .Y(new_new_n456_));
  NOi21      g434(.An(i_2_), .B(i_7_), .Y(new_new_n457_));
  NAi31      g435(.An(i_11_), .B(new_new_n457_), .C(new_new_n993_), .Y(new_new_n458_));
  INV        g436(.A(new_new_n404_), .Y(new_new_n459_));
  NA3        g437(.A(new_new_n459_), .B(new_new_n432_), .C(new_new_n72_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n460_), .B(new_new_n458_), .Y(new_new_n461_));
  NO2        g439(.A(i_6_), .B(i_10_), .Y(new_new_n462_));
  NA4        g440(.A(new_new_n462_), .B(new_new_n300_), .C(i_8_), .D(new_new_n233_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n463_), .B(new_new_n152_), .Y(new_new_n464_));
  NA3        g442(.A(new_new_n240_), .B(new_new_n168_), .C(new_new_n129_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n466_));
  NO2        g444(.A(new_new_n154_), .B(i_3_), .Y(new_new_n467_));
  NAi31      g445(.An(new_new_n466_), .B(new_new_n467_), .C(new_new_n223_), .Y(new_new_n468_));
  NA3        g446(.A(new_new_n381_), .B(new_new_n175_), .C(new_new_n146_), .Y(new_new_n469_));
  NA3        g447(.A(new_new_n469_), .B(new_new_n468_), .C(new_new_n465_), .Y(new_new_n470_));
  NO4        g448(.A(new_new_n470_), .B(new_new_n464_), .C(new_new_n461_), .D(new_new_n452_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n441_), .B(new_new_n377_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n472_), .B(new_new_n221_), .Y(new_new_n473_));
  NAi21      g451(.An(new_new_n212_), .B(new_new_n385_), .Y(new_new_n474_));
  NA3        g452(.A(new_new_n992_), .B(i_3_), .C(new_new_n139_), .Y(new_new_n475_));
  OR3        g453(.A(new_new_n290_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n476_));
  NO2        g454(.A(new_new_n476_), .B(new_new_n475_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n27_), .B(i_10_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n478_), .B(new_new_n449_), .Y(new_new_n479_));
  NA3        g457(.A(new_new_n293_), .B(new_new_n220_), .C(new_new_n70_), .Y(new_new_n480_));
  NO2        g458(.A(new_new_n480_), .B(new_new_n455_), .Y(new_new_n481_));
  NO4        g459(.A(new_new_n481_), .B(new_new_n479_), .C(new_new_n477_), .D(new_new_n473_), .Y(new_new_n482_));
  NA4        g460(.A(new_new_n482_), .B(new_new_n471_), .C(new_new_n448_), .D(new_new_n446_), .Y(new_new_n483_));
  AN2        g461(.A(new_new_n274_), .B(new_new_n231_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n484_), .B(new_new_n172_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n119_), .B(new_new_n108_), .Y(new_new_n486_));
  AN2        g464(.A(new_new_n486_), .B(new_new_n437_), .Y(new_new_n487_));
  OAI210     g465(.A0(i_2_), .A1(new_new_n229_), .B0(new_new_n294_), .Y(new_new_n488_));
  AOI220     g466(.A0(new_new_n488_), .A1(new_new_n309_), .B0(new_new_n487_), .B1(new_new_n296_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n344_), .B(new_new_n70_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n357_), .B(new_new_n353_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n36_), .B(i_8_), .Y(new_new_n492_));
  NAi41      g470(.An(new_new_n490_), .B(new_new_n462_), .C(new_new_n492_), .D(new_new_n47_), .Y(new_new_n493_));
  AOI210     g471(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n405_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n494_), .B(new_new_n493_), .Y(new_new_n495_));
  INV        g473(.A(new_new_n495_), .Y(new_new_n496_));
  INV        g474(.A(new_new_n248_), .Y(new_new_n497_));
  OAI210     g475(.A0(i_8_), .A1(new_new_n497_), .B0(new_new_n131_), .Y(new_new_n498_));
  NO2        g476(.A(i_7_), .B(new_new_n194_), .Y(new_new_n499_));
  OR2        g477(.A(new_new_n179_), .B(i_4_), .Y(new_new_n500_));
  INV        g478(.A(new_new_n500_), .Y(new_new_n501_));
  AOI220     g479(.A0(new_new_n501_), .A1(new_new_n499_), .B0(new_new_n498_), .B1(new_new_n406_), .Y(new_new_n502_));
  NA4        g480(.A(new_new_n502_), .B(new_new_n496_), .C(new_new_n489_), .D(new_new_n485_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n376_), .B(new_new_n282_), .Y(new_new_n504_));
  NA2        g482(.A(new_new_n372_), .B(new_new_n504_), .Y(new_new_n505_));
  NO2        g483(.A(i_12_), .B(new_new_n189_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n506_), .B(new_new_n222_), .Y(new_new_n507_));
  NA2        g485(.A(new_new_n462_), .B(new_new_n27_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n508_), .B(new_new_n507_), .Y(new_new_n509_));
  NOi31      g487(.An(new_new_n301_), .B(new_new_n404_), .C(new_new_n38_), .Y(new_new_n510_));
  OAI210     g488(.A0(new_new_n510_), .A1(new_new_n509_), .B0(new_new_n505_), .Y(new_new_n511_));
  NO2        g489(.A(i_8_), .B(i_7_), .Y(new_new_n512_));
  INV        g490(.A(new_new_n220_), .Y(new_new_n513_));
  OAI220     g491(.A0(new_new_n47_), .A1(new_new_n500_), .B0(new_new_n513_), .B1(new_new_n237_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n45_), .B(i_10_), .Y(new_new_n515_));
  NO2        g493(.A(new_new_n515_), .B(i_6_), .Y(new_new_n516_));
  NA3        g494(.A(new_new_n516_), .B(new_new_n514_), .C(new_new_n512_), .Y(new_new_n517_));
  AOI210     g495(.A0(new_new_n417_), .A1(new_new_n310_), .B0(new_new_n242_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n518_), .B(new_new_n251_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n519_), .B(new_new_n254_), .Y(new_new_n520_));
  NOi31      g498(.An(new_new_n277_), .B(new_new_n288_), .C(new_new_n177_), .Y(new_new_n521_));
  NA3        g499(.A(new_new_n293_), .B(new_new_n170_), .C(new_new_n92_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n218_), .B(new_new_n45_), .Y(new_new_n523_));
  NO2        g501(.A(new_new_n154_), .B(i_5_), .Y(new_new_n524_));
  NA2        g502(.A(new_new_n524_), .B(new_new_n303_), .Y(new_new_n525_));
  OAI210     g503(.A0(new_new_n525_), .A1(new_new_n523_), .B0(new_new_n522_), .Y(new_new_n526_));
  OAI210     g504(.A0(new_new_n526_), .A1(new_new_n521_), .B0(new_new_n441_), .Y(new_new_n527_));
  NA4        g505(.A(new_new_n527_), .B(new_new_n520_), .C(new_new_n517_), .D(new_new_n511_), .Y(new_new_n528_));
  NA3        g506(.A(new_new_n214_), .B(new_new_n68_), .C(new_new_n45_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n271_), .B(new_new_n80_), .Y(new_new_n530_));
  AOI210     g508(.A0(new_new_n529_), .A1(new_new_n335_), .B0(new_new_n530_), .Y(new_new_n531_));
  NA2        g509(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n434_), .B(new_new_n218_), .Y(new_new_n533_));
  NO2        g511(.A(new_new_n532_), .B(new_new_n533_), .Y(new_new_n534_));
  NA2        g512(.A(i_0_), .B(new_new_n49_), .Y(new_new_n535_));
  NA3        g513(.A(new_new_n506_), .B(new_new_n262_), .C(new_new_n535_), .Y(new_new_n536_));
  NO2        g514(.A(i_1_), .B(new_new_n536_), .Y(new_new_n537_));
  NO3        g515(.A(new_new_n537_), .B(new_new_n534_), .C(new_new_n531_), .Y(new_new_n538_));
  NO4        g516(.A(i_1_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n539_));
  NO3        g517(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n230_), .B(new_new_n36_), .Y(new_new_n541_));
  AN2        g519(.A(new_new_n541_), .B(new_new_n540_), .Y(new_new_n542_));
  OA210      g520(.A0(new_new_n542_), .A1(new_new_n539_), .B0(new_new_n344_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n404_), .B(i_1_), .Y(new_new_n544_));
  NOi31      g522(.An(new_new_n544_), .B(new_new_n438_), .C(new_new_n70_), .Y(new_new_n545_));
  AN3        g523(.A(new_new_n545_), .B(new_new_n401_), .C(i_3_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n415_), .B(new_new_n173_), .Y(new_new_n547_));
  NO3        g525(.A(new_new_n547_), .B(new_new_n546_), .C(new_new_n543_), .Y(new_new_n548_));
  NOi21      g526(.An(i_10_), .B(i_6_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n82_), .B(new_new_n25_), .Y(new_new_n550_));
  AOI220     g528(.A0(new_new_n271_), .A1(new_new_n550_), .B0(new_new_n262_), .B1(new_new_n549_), .Y(new_new_n551_));
  NO2        g529(.A(new_new_n551_), .B(new_new_n436_), .Y(new_new_n552_));
  NO2        g530(.A(new_new_n111_), .B(new_new_n23_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n301_), .B(new_new_n161_), .Y(new_new_n554_));
  AOI220     g532(.A0(new_new_n554_), .A1(new_new_n424_), .B0(new_new_n169_), .B1(new_new_n178_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n555_), .B(new_new_n552_), .Y(new_new_n556_));
  NO2        g534(.A(new_new_n490_), .B(new_new_n365_), .Y(new_new_n557_));
  INV        g535(.A(new_new_n303_), .Y(new_new_n558_));
  NO2        g536(.A(i_12_), .B(new_new_n82_), .Y(new_new_n559_));
  NA3        g537(.A(new_new_n559_), .B(new_new_n262_), .C(new_new_n535_), .Y(new_new_n560_));
  NA3        g538(.A(new_new_n373_), .B(new_new_n271_), .C(new_new_n214_), .Y(new_new_n561_));
  AOI210     g539(.A0(new_new_n561_), .A1(new_new_n560_), .B0(new_new_n558_), .Y(new_new_n562_));
  NO3        g540(.A(i_4_), .B(new_new_n327_), .C(new_new_n288_), .Y(new_new_n563_));
  OR2        g541(.A(i_2_), .B(i_5_), .Y(new_new_n564_));
  OR2        g542(.A(new_new_n564_), .B(new_new_n396_), .Y(new_new_n565_));
  NO2        g543(.A(new_new_n565_), .B(new_new_n474_), .Y(new_new_n566_));
  NO4        g544(.A(new_new_n566_), .B(new_new_n563_), .C(new_new_n562_), .D(new_new_n557_), .Y(new_new_n567_));
  NA4        g545(.A(new_new_n567_), .B(new_new_n556_), .C(new_new_n548_), .D(new_new_n538_), .Y(new_new_n568_));
  NO4        g546(.A(new_new_n568_), .B(new_new_n528_), .C(new_new_n503_), .D(new_new_n483_), .Y(new_new_n569_));
  NA4        g547(.A(new_new_n569_), .B(new_new_n431_), .C(new_new_n343_), .D(new_new_n299_), .Y(men7));
  NO2        g548(.A(new_new_n88_), .B(new_new_n55_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n104_), .B(new_new_n85_), .Y(new_new_n572_));
  NA2        g550(.A(new_new_n462_), .B(new_new_n80_), .Y(new_new_n573_));
  NA2        g551(.A(i_11_), .B(new_new_n189_), .Y(new_new_n574_));
  NA3        g552(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n575_));
  NO2        g553(.A(new_new_n233_), .B(i_4_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n576_), .B(i_8_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n101_), .B(new_new_n575_), .Y(new_new_n578_));
  NA2        g556(.A(i_2_), .B(new_new_n82_), .Y(new_new_n579_));
  OAI210     g557(.A0(new_new_n83_), .A1(new_new_n198_), .B0(new_new_n199_), .Y(new_new_n580_));
  NA2        g558(.A(i_4_), .B(i_8_), .Y(new_new_n581_));
  OAI220     g559(.A0(new_new_n991_), .A1(new_new_n579_), .B0(new_new_n580_), .B1(i_13_), .Y(new_new_n582_));
  NO4        g560(.A(new_new_n582_), .B(new_new_n578_), .C(new_new_n572_), .D(new_new_n571_), .Y(new_new_n583_));
  INV        g561(.A(new_new_n158_), .Y(new_new_n584_));
  OR2        g562(.A(i_6_), .B(i_10_), .Y(new_new_n585_));
  NO2        g563(.A(new_new_n585_), .B(new_new_n23_), .Y(new_new_n586_));
  OR3        g564(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n587_));
  NO3        g565(.A(new_new_n587_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n588_));
  INV        g566(.A(new_new_n195_), .Y(new_new_n589_));
  NO2        g567(.A(new_new_n588_), .B(new_new_n586_), .Y(new_new_n590_));
  OA220      g568(.A0(new_new_n590_), .A1(new_new_n558_), .B0(new_new_n584_), .B1(new_new_n256_), .Y(new_new_n591_));
  AOI210     g569(.A0(new_new_n591_), .A1(new_new_n583_), .B0(new_new_n64_), .Y(new_new_n592_));
  NOi21      g570(.An(i_11_), .B(i_7_), .Y(new_new_n593_));
  AO210      g571(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n594_));
  NO2        g572(.A(new_new_n594_), .B(new_new_n593_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n595_), .B(new_new_n201_), .Y(new_new_n596_));
  NA3        g574(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n597_));
  NAi31      g575(.An(new_new_n597_), .B(new_new_n211_), .C(i_11_), .Y(new_new_n598_));
  AOI210     g576(.A0(new_new_n598_), .A1(new_new_n596_), .B0(new_new_n64_), .Y(new_new_n599_));
  NA2        g577(.A(new_new_n223_), .B(new_new_n64_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n397_), .B(new_new_n31_), .Y(new_new_n601_));
  OR2        g579(.A(new_new_n203_), .B(new_new_n104_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n602_), .B(new_new_n601_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n64_), .B(i_9_), .Y(new_new_n604_));
  NA2        g582(.A(new_new_n64_), .B(new_new_n603_), .Y(new_new_n605_));
  NO2        g583(.A(i_1_), .B(i_12_), .Y(new_new_n606_));
  NA2        g584(.A(new_new_n605_), .B(new_new_n600_), .Y(new_new_n607_));
  OAI210     g585(.A0(new_new_n607_), .A1(new_new_n599_), .B0(i_6_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n233_), .B(new_new_n82_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n609_), .B(i_11_), .Y(new_new_n610_));
  NO4        g588(.A(new_new_n211_), .B(new_new_n125_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n611_), .B(new_new_n604_), .Y(new_new_n612_));
  NA2        g590(.A(new_new_n233_), .B(i_6_), .Y(new_new_n613_));
  NO3        g591(.A(new_new_n585_), .B(new_new_n230_), .C(new_new_n23_), .Y(new_new_n614_));
  INV        g592(.A(new_new_n614_), .Y(new_new_n615_));
  OAI210     g593(.A0(new_new_n615_), .A1(new_new_n45_), .B0(new_new_n612_), .Y(new_new_n616_));
  NA3        g594(.A(new_new_n512_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n617_));
  NA2        g595(.A(new_new_n135_), .B(i_9_), .Y(new_new_n618_));
  NA3        g596(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n47_), .B(i_1_), .Y(new_new_n620_));
  NA3        g598(.A(new_new_n620_), .B(new_new_n255_), .C(new_new_n45_), .Y(new_new_n621_));
  OAI220     g599(.A0(new_new_n621_), .A1(new_new_n619_), .B0(new_new_n618_), .B1(new_new_n987_), .Y(new_new_n622_));
  NA3        g600(.A(new_new_n604_), .B(new_new_n303_), .C(i_6_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n623_), .B(new_new_n23_), .Y(new_new_n624_));
  AOI210     g602(.A0(new_new_n456_), .A1(new_new_n408_), .B0(new_new_n236_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(new_new_n579_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n620_), .B(new_new_n255_), .Y(new_new_n627_));
  NO2        g605(.A(i_11_), .B(new_new_n37_), .Y(new_new_n628_));
  NA2        g606(.A(new_new_n628_), .B(new_new_n24_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n629_), .B(new_new_n627_), .Y(new_new_n630_));
  OR4        g608(.A(new_new_n630_), .B(new_new_n626_), .C(new_new_n624_), .D(new_new_n622_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n631_), .B(new_new_n616_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n233_), .B(new_new_n97_), .Y(new_new_n633_));
  NO2        g611(.A(new_new_n633_), .B(new_new_n593_), .Y(new_new_n634_));
  NA2        g612(.A(new_new_n634_), .B(i_1_), .Y(new_new_n635_));
  NO2        g613(.A(new_new_n635_), .B(new_new_n587_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n403_), .B(new_new_n82_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n636_), .B(new_new_n47_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n114_), .B(new_new_n37_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n82_), .B(i_9_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n640_), .B(new_new_n64_), .Y(new_new_n641_));
  NA2        g619(.A(i_1_), .B(i_3_), .Y(new_new_n642_));
  NA3        g620(.A(new_new_n638_), .B(new_new_n632_), .C(new_new_n608_), .Y(new_new_n643_));
  NO3        g621(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n644_));
  NOi21      g622(.An(new_new_n644_), .B(i_10_), .Y(new_new_n645_));
  OA210      g623(.A0(new_new_n645_), .A1(new_new_n240_), .B0(new_new_n82_), .Y(new_new_n646_));
  NO3        g624(.A(new_new_n457_), .B(new_new_n581_), .C(new_new_n82_), .Y(new_new_n647_));
  NA2        g625(.A(new_new_n647_), .B(new_new_n25_), .Y(new_new_n648_));
  INV        g626(.A(new_new_n648_), .Y(new_new_n649_));
  OAI210     g627(.A0(new_new_n649_), .A1(new_new_n646_), .B0(i_1_), .Y(new_new_n650_));
  AOI210     g628(.A0(new_new_n255_), .A1(new_new_n93_), .B0(i_1_), .Y(new_new_n651_));
  NO2        g629(.A(new_new_n355_), .B(i_2_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n652_), .B(new_new_n651_), .Y(new_new_n653_));
  OAI210     g631(.A0(new_new_n623_), .A1(new_new_n435_), .B0(new_new_n653_), .Y(new_new_n654_));
  INV        g632(.A(new_new_n654_), .Y(new_new_n655_));
  AOI210     g633(.A0(new_new_n655_), .A1(new_new_n650_), .B0(i_13_), .Y(new_new_n656_));
  OR2        g634(.A(i_11_), .B(i_7_), .Y(new_new_n657_));
  NA3        g635(.A(new_new_n657_), .B(new_new_n102_), .C(new_new_n135_), .Y(new_new_n658_));
  AOI220     g636(.A0(new_new_n451_), .A1(new_new_n158_), .B0(i_2_), .B1(new_new_n135_), .Y(new_new_n659_));
  OAI210     g637(.A0(new_new_n659_), .A1(new_new_n45_), .B0(new_new_n658_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n457_), .B(new_new_n24_), .Y(new_new_n661_));
  AOI220     g639(.A0(new_new_n661_), .A1(new_new_n637_), .B0(new_new_n240_), .B1(new_new_n128_), .Y(new_new_n662_));
  NO2        g640(.A(new_new_n662_), .B(new_new_n41_), .Y(new_new_n663_));
  AOI210     g641(.A0(new_new_n660_), .A1(new_new_n318_), .B0(new_new_n663_), .Y(new_new_n664_));
  AOI210     g642(.A0(new_new_n435_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n665_));
  NOi31      g643(.An(new_new_n665_), .B(new_new_n573_), .C(new_new_n45_), .Y(new_new_n666_));
  NA2        g644(.A(new_new_n124_), .B(i_13_), .Y(new_new_n667_));
  NO2        g645(.A(new_new_n619_), .B(new_new_n111_), .Y(new_new_n668_));
  INV        g646(.A(new_new_n668_), .Y(new_new_n669_));
  OAI220     g647(.A0(new_new_n669_), .A1(new_new_n68_), .B0(new_new_n667_), .B1(new_new_n651_), .Y(new_new_n670_));
  NO3        g648(.A(new_new_n68_), .B(new_new_n32_), .C(new_new_n97_), .Y(new_new_n671_));
  NA2        g649(.A(new_new_n26_), .B(new_new_n189_), .Y(new_new_n672_));
  NA2        g650(.A(new_new_n672_), .B(i_7_), .Y(new_new_n673_));
  NO3        g651(.A(new_new_n457_), .B(new_new_n233_), .C(new_new_n82_), .Y(new_new_n674_));
  AOI210     g652(.A0(new_new_n674_), .A1(new_new_n673_), .B0(new_new_n671_), .Y(new_new_n675_));
  AOI220     g653(.A0(new_new_n373_), .A1(new_new_n620_), .B0(new_new_n87_), .B1(new_new_n98_), .Y(new_new_n676_));
  OAI220     g654(.A0(new_new_n676_), .A1(new_new_n577_), .B0(new_new_n675_), .B1(new_new_n589_), .Y(new_new_n677_));
  NO3        g655(.A(new_new_n677_), .B(new_new_n670_), .C(new_new_n666_), .Y(new_new_n678_));
  OR2        g656(.A(i_11_), .B(i_6_), .Y(new_new_n679_));
  NA3        g657(.A(new_new_n576_), .B(new_new_n672_), .C(i_7_), .Y(new_new_n680_));
  AOI210     g658(.A0(new_new_n680_), .A1(new_new_n669_), .B0(new_new_n679_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n610_), .B(i_13_), .Y(new_new_n682_));
  NAi21      g660(.An(i_11_), .B(i_12_), .Y(new_new_n683_));
  NO2        g661(.A(new_new_n559_), .B(new_new_n581_), .Y(new_new_n684_));
  NA2        g662(.A(new_new_n684_), .B(new_new_n300_), .Y(new_new_n685_));
  NA2        g663(.A(new_new_n685_), .B(new_new_n682_), .Y(new_new_n686_));
  OAI210     g664(.A0(new_new_n686_), .A1(new_new_n681_), .B0(new_new_n64_), .Y(new_new_n687_));
  NO2        g665(.A(i_2_), .B(i_12_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n354_), .B(new_new_n688_), .Y(new_new_n689_));
  NO2        g667(.A(new_new_n125_), .B(i_2_), .Y(new_new_n690_));
  NA2        g668(.A(new_new_n690_), .B(new_new_n606_), .Y(new_new_n691_));
  NA2        g669(.A(new_new_n691_), .B(new_new_n689_), .Y(new_new_n692_));
  NA3        g670(.A(new_new_n692_), .B(new_new_n46_), .C(new_new_n222_), .Y(new_new_n693_));
  NA4        g671(.A(new_new_n693_), .B(new_new_n687_), .C(new_new_n678_), .D(new_new_n664_), .Y(new_new_n694_));
  OR4        g672(.A(new_new_n694_), .B(new_new_n656_), .C(new_new_n643_), .D(new_new_n592_), .Y(men5));
  AOI210     g673(.A0(new_new_n634_), .A1(new_new_n258_), .B0(new_new_n406_), .Y(new_new_n696_));
  AN2        g674(.A(new_new_n24_), .B(i_10_), .Y(new_new_n697_));
  NA3        g675(.A(new_new_n697_), .B(new_new_n688_), .C(new_new_n104_), .Y(new_new_n698_));
  NO2        g676(.A(new_new_n577_), .B(i_11_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n83_), .B(new_new_n699_), .Y(new_new_n700_));
  NA3        g678(.A(new_new_n700_), .B(new_new_n698_), .C(new_new_n696_), .Y(new_new_n701_));
  NO3        g679(.A(i_11_), .B(new_new_n233_), .C(i_13_), .Y(new_new_n702_));
  NO2        g680(.A(new_new_n121_), .B(new_new_n23_), .Y(new_new_n703_));
  NA2        g681(.A(i_12_), .B(i_8_), .Y(new_new_n704_));
  OAI210     g682(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n704_), .Y(new_new_n705_));
  INV        g683(.A(new_new_n434_), .Y(new_new_n706_));
  AOI220     g684(.A0(new_new_n303_), .A1(new_new_n553_), .B0(new_new_n705_), .B1(new_new_n703_), .Y(new_new_n707_));
  INV        g685(.A(new_new_n707_), .Y(new_new_n708_));
  NO2        g686(.A(new_new_n708_), .B(new_new_n701_), .Y(new_new_n709_));
  INV        g687(.A(new_new_n168_), .Y(new_new_n710_));
  NA2        g688(.A(new_new_n652_), .B(new_new_n107_), .Y(new_new_n711_));
  NO2        g689(.A(new_new_n711_), .B(new_new_n710_), .Y(new_new_n712_));
  NO2        g690(.A(new_new_n439_), .B(new_new_n26_), .Y(new_new_n713_));
  NO2        g691(.A(new_new_n713_), .B(new_new_n408_), .Y(new_new_n714_));
  NA2        g692(.A(new_new_n714_), .B(i_2_), .Y(new_new_n715_));
  INV        g693(.A(new_new_n715_), .Y(new_new_n716_));
  AOI210     g694(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n404_), .Y(new_new_n717_));
  AOI210     g695(.A0(new_new_n717_), .A1(new_new_n716_), .B0(new_new_n712_), .Y(new_new_n718_));
  NO2        g696(.A(new_new_n186_), .B(new_new_n122_), .Y(new_new_n719_));
  OAI210     g697(.A0(new_new_n719_), .A1(new_new_n703_), .B0(i_2_), .Y(new_new_n720_));
  NO3        g698(.A(new_new_n594_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n721_));
  AOI210     g699(.A0(new_new_n990_), .A1(new_new_n720_), .B0(new_new_n189_), .Y(new_new_n722_));
  OA210      g700(.A0(new_new_n595_), .A1(new_new_n123_), .B0(i_13_), .Y(new_new_n723_));
  NA2        g701(.A(new_new_n149_), .B(new_new_n574_), .Y(new_new_n724_));
  NO2        g702(.A(new_new_n724_), .B(new_new_n359_), .Y(new_new_n725_));
  AOI210     g703(.A0(new_new_n203_), .A1(new_new_n145_), .B0(new_new_n492_), .Y(new_new_n726_));
  NA2        g704(.A(new_new_n726_), .B(new_new_n408_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n98_), .B(new_new_n45_), .Y(new_new_n728_));
  INV        g706(.A(new_new_n289_), .Y(new_new_n729_));
  NA4        g707(.A(new_new_n729_), .B(new_new_n293_), .C(new_new_n121_), .D(new_new_n43_), .Y(new_new_n730_));
  OAI210     g708(.A0(new_new_n730_), .A1(new_new_n728_), .B0(new_new_n727_), .Y(new_new_n731_));
  NO4        g709(.A(new_new_n731_), .B(new_new_n725_), .C(new_new_n723_), .D(new_new_n722_), .Y(new_new_n732_));
  NA2        g710(.A(new_new_n553_), .B(new_new_n28_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n702_), .B(new_new_n263_), .Y(new_new_n734_));
  NA2        g712(.A(new_new_n734_), .B(new_new_n733_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n63_), .B(i_12_), .Y(new_new_n736_));
  NO2        g714(.A(new_new_n736_), .B(new_new_n123_), .Y(new_new_n737_));
  NO2        g715(.A(new_new_n737_), .B(new_new_n574_), .Y(new_new_n738_));
  AOI220     g716(.A0(new_new_n738_), .A1(new_new_n36_), .B0(new_new_n735_), .B1(new_new_n47_), .Y(new_new_n739_));
  NA4        g717(.A(new_new_n739_), .B(new_new_n732_), .C(new_new_n718_), .D(new_new_n709_), .Y(men6));
  NO3        g718(.A(new_new_n246_), .B(new_new_n295_), .C(i_1_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n181_), .B(new_new_n136_), .Y(new_new_n742_));
  OAI210     g720(.A0(new_new_n742_), .A1(new_new_n741_), .B0(new_new_n690_), .Y(new_new_n743_));
  NO2        g721(.A(new_new_n217_), .B(new_new_n466_), .Y(new_new_n744_));
  AO210      g722(.A0(new_new_n988_), .A1(new_new_n743_), .B0(i_12_), .Y(new_new_n745_));
  NA2        g723(.A(new_new_n645_), .B(new_new_n70_), .Y(new_new_n746_));
  INV        g724(.A(new_new_n314_), .Y(new_new_n747_));
  NA2        g725(.A(new_new_n72_), .B(new_new_n128_), .Y(new_new_n748_));
  INV        g726(.A(new_new_n121_), .Y(new_new_n749_));
  NA2        g727(.A(new_new_n749_), .B(new_new_n47_), .Y(new_new_n750_));
  AOI210     g728(.A0(new_new_n750_), .A1(new_new_n748_), .B0(new_new_n747_), .Y(new_new_n751_));
  NO2        g729(.A(new_new_n32_), .B(i_11_), .Y(new_new_n752_));
  NA3        g730(.A(new_new_n752_), .B(new_new_n454_), .C(new_new_n377_), .Y(new_new_n753_));
  NAi32      g731(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n679_), .B(new_new_n754_), .Y(new_new_n755_));
  OAI210     g733(.A0(new_new_n644_), .A1(new_new_n541_), .B0(new_new_n540_), .Y(new_new_n756_));
  NAi31      g734(.An(new_new_n755_), .B(new_new_n756_), .C(new_new_n753_), .Y(new_new_n757_));
  OR2        g735(.A(new_new_n757_), .B(new_new_n751_), .Y(new_new_n758_));
  NO2        g736(.A(new_new_n657_), .B(i_2_), .Y(new_new_n759_));
  NA2        g737(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n760_));
  NO2        g738(.A(new_new_n760_), .B(new_new_n396_), .Y(new_new_n761_));
  NA2        g739(.A(new_new_n761_), .B(new_new_n759_), .Y(new_new_n762_));
  AO210      g740(.A0(new_new_n348_), .A1(new_new_n339_), .B0(new_new_n384_), .Y(new_new_n763_));
  NA3        g741(.A(new_new_n763_), .B(new_new_n247_), .C(i_7_), .Y(new_new_n764_));
  BUFFER     g742(.A(new_new_n595_), .Y(new_new_n765_));
  NA2        g743(.A(new_new_n765_), .B(new_new_n144_), .Y(new_new_n766_));
  AO210      g744(.A0(new_new_n472_), .A1(new_new_n706_), .B0(new_new_n36_), .Y(new_new_n767_));
  NA4        g745(.A(new_new_n767_), .B(new_new_n766_), .C(new_new_n764_), .D(new_new_n762_), .Y(new_new_n768_));
  NO2        g746(.A(new_new_n609_), .B(i_11_), .Y(new_new_n769_));
  AOI220     g747(.A0(new_new_n769_), .A1(new_new_n540_), .B0(new_new_n744_), .B1(new_new_n673_), .Y(new_new_n770_));
  NA3        g748(.A(new_new_n359_), .B(new_new_n234_), .C(new_new_n144_), .Y(new_new_n771_));
  NA2        g749(.A(new_new_n384_), .B(new_new_n67_), .Y(new_new_n772_));
  NA4        g750(.A(new_new_n772_), .B(new_new_n771_), .C(new_new_n770_), .D(new_new_n580_), .Y(new_new_n773_));
  NO2        g751(.A(new_new_n585_), .B(new_new_n98_), .Y(new_new_n774_));
  OAI210     g752(.A0(new_new_n774_), .A1(new_new_n108_), .B0(new_new_n394_), .Y(new_new_n775_));
  INV        g753(.A(new_new_n565_), .Y(new_new_n776_));
  NA3        g754(.A(new_new_n776_), .B(new_new_n314_), .C(i_7_), .Y(new_new_n777_));
  NA2        g755(.A(new_new_n777_), .B(new_new_n775_), .Y(new_new_n778_));
  NO4        g756(.A(new_new_n778_), .B(new_new_n773_), .C(new_new_n768_), .D(new_new_n758_), .Y(new_new_n779_));
  NA4        g757(.A(new_new_n779_), .B(new_new_n746_), .C(new_new_n745_), .D(new_new_n367_), .Y(men3));
  NA2        g758(.A(i_6_), .B(i_7_), .Y(new_new_n781_));
  NO2        g759(.A(new_new_n781_), .B(i_0_), .Y(new_new_n782_));
  NO2        g760(.A(i_11_), .B(new_new_n233_), .Y(new_new_n783_));
  OAI210     g761(.A0(new_new_n782_), .A1(new_new_n277_), .B0(new_new_n783_), .Y(new_new_n784_));
  INV        g762(.A(new_new_n784_), .Y(new_new_n785_));
  NO3        g763(.A(new_new_n436_), .B(new_new_n85_), .C(new_new_n45_), .Y(new_new_n786_));
  OA210      g764(.A0(new_new_n786_), .A1(new_new_n785_), .B0(new_new_n170_), .Y(new_new_n787_));
  NA3        g765(.A(new_new_n771_), .B(new_new_n580_), .C(new_new_n358_), .Y(new_new_n788_));
  NA2        g766(.A(new_new_n788_), .B(new_new_n40_), .Y(new_new_n789_));
  NO3        g767(.A(new_new_n602_), .B(new_new_n439_), .C(new_new_n128_), .Y(new_new_n790_));
  AN2        g768(.A(new_new_n438_), .B(new_new_n56_), .Y(new_new_n791_));
  NO2        g769(.A(new_new_n791_), .B(new_new_n790_), .Y(new_new_n792_));
  AOI210     g770(.A0(new_new_n792_), .A1(new_new_n789_), .B0(new_new_n49_), .Y(new_new_n793_));
  NO4        g771(.A(new_new_n363_), .B(new_new_n370_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n181_), .B(new_new_n549_), .Y(new_new_n795_));
  NOi21      g773(.An(new_new_n795_), .B(new_new_n794_), .Y(new_new_n796_));
  NA2        g774(.A(new_new_n665_), .B(new_new_n640_), .Y(new_new_n797_));
  NA2        g775(.A(new_new_n319_), .B(i_5_), .Y(new_new_n798_));
  OAI220     g776(.A0(new_new_n798_), .A1(new_new_n797_), .B0(new_new_n796_), .B1(new_new_n64_), .Y(new_new_n799_));
  NOi21      g777(.An(i_5_), .B(i_9_), .Y(new_new_n800_));
  NA2        g778(.A(new_new_n800_), .B(new_new_n433_), .Y(new_new_n801_));
  AOI210     g779(.A0(new_new_n255_), .A1(new_new_n456_), .B0(new_new_n647_), .Y(new_new_n802_));
  NO3        g780(.A(new_new_n400_), .B(new_new_n255_), .C(new_new_n70_), .Y(new_new_n803_));
  NO2        g781(.A(new_new_n171_), .B(new_new_n145_), .Y(new_new_n804_));
  INV        g782(.A(new_new_n803_), .Y(new_new_n805_));
  OAI220     g783(.A0(new_new_n805_), .A1(new_new_n177_), .B0(new_new_n802_), .B1(new_new_n801_), .Y(new_new_n806_));
  NO4        g784(.A(new_new_n806_), .B(new_new_n799_), .C(new_new_n793_), .D(new_new_n787_), .Y(new_new_n807_));
  NA2        g785(.A(new_new_n181_), .B(new_new_n24_), .Y(new_new_n808_));
  NO2        g786(.A(new_new_n639_), .B(new_new_n572_), .Y(new_new_n809_));
  NO2        g787(.A(new_new_n809_), .B(new_new_n808_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n300_), .B(new_new_n126_), .Y(new_new_n811_));
  NAi21      g789(.An(new_new_n159_), .B(i_5_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n811_), .B(new_new_n386_), .Y(new_new_n813_));
  NO2        g791(.A(new_new_n813_), .B(new_new_n810_), .Y(new_new_n814_));
  NO2        g792(.A(new_new_n377_), .B(new_new_n281_), .Y(new_new_n815_));
  NA2        g793(.A(new_new_n815_), .B(new_new_n668_), .Y(new_new_n816_));
  NA2        g794(.A(new_new_n550_), .B(i_0_), .Y(new_new_n817_));
  NO2        g795(.A(new_new_n817_), .B(new_new_n372_), .Y(new_new_n818_));
  INV        g796(.A(new_new_n818_), .Y(new_new_n819_));
  AN2        g797(.A(new_new_n92_), .B(new_new_n238_), .Y(new_new_n820_));
  NA2        g798(.A(new_new_n702_), .B(new_new_n315_), .Y(new_new_n821_));
  AOI210     g799(.A0(new_new_n462_), .A1(new_new_n83_), .B0(new_new_n59_), .Y(new_new_n822_));
  OAI220     g800(.A0(new_new_n822_), .A1(new_new_n821_), .B0(new_new_n629_), .B1(new_new_n513_), .Y(new_new_n823_));
  NA2        g801(.A(i_0_), .B(i_10_), .Y(new_new_n824_));
  NA2        g802(.A(new_new_n319_), .B(new_new_n94_), .Y(new_new_n825_));
  NA2        g803(.A(new_new_n544_), .B(i_4_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n184_), .B(new_new_n198_), .Y(new_new_n827_));
  OAI220     g805(.A0(new_new_n827_), .A1(new_new_n821_), .B0(new_new_n826_), .B1(new_new_n825_), .Y(new_new_n828_));
  NO3        g806(.A(new_new_n828_), .B(new_new_n823_), .C(new_new_n820_), .Y(new_new_n829_));
  NA4        g807(.A(new_new_n829_), .B(new_new_n819_), .C(new_new_n816_), .D(new_new_n814_), .Y(new_new_n830_));
  NO2        g808(.A(new_new_n99_), .B(new_new_n37_), .Y(new_new_n831_));
  NA2        g809(.A(i_11_), .B(i_9_), .Y(new_new_n832_));
  NO3        g810(.A(i_12_), .B(new_new_n832_), .C(new_new_n579_), .Y(new_new_n833_));
  AN2        g811(.A(new_new_n833_), .B(new_new_n831_), .Y(new_new_n834_));
  NO2        g812(.A(new_new_n49_), .B(i_7_), .Y(new_new_n835_));
  NA2        g813(.A(new_new_n381_), .B(new_new_n175_), .Y(new_new_n836_));
  NA2        g814(.A(new_new_n836_), .B(new_new_n157_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n171_), .B(i_0_), .Y(new_new_n838_));
  INV        g816(.A(new_new_n838_), .Y(new_new_n839_));
  NA2        g817(.A(new_new_n454_), .B(new_new_n228_), .Y(new_new_n840_));
  AOI210     g818(.A0(new_new_n357_), .A1(new_new_n42_), .B0(new_new_n393_), .Y(new_new_n841_));
  OAI220     g819(.A0(new_new_n841_), .A1(new_new_n801_), .B0(new_new_n840_), .B1(new_new_n839_), .Y(new_new_n842_));
  NO3        g820(.A(new_new_n842_), .B(new_new_n837_), .C(new_new_n834_), .Y(new_new_n843_));
  NA2        g821(.A(new_new_n628_), .B(new_new_n118_), .Y(new_new_n844_));
  NO2        g822(.A(i_6_), .B(new_new_n844_), .Y(new_new_n845_));
  AOI210     g823(.A0(new_new_n435_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n846_));
  NA2        g824(.A(new_new_n168_), .B(new_new_n99_), .Y(new_new_n847_));
  NOi32      g825(.An(new_new_n846_), .Bn(new_new_n184_), .C(new_new_n847_), .Y(new_new_n848_));
  NO2        g826(.A(new_new_n848_), .B(new_new_n845_), .Y(new_new_n849_));
  NOi21      g827(.An(i_7_), .B(i_5_), .Y(new_new_n850_));
  NOi31      g828(.An(new_new_n850_), .B(i_0_), .C(new_new_n683_), .Y(new_new_n851_));
  OR2        g829(.A(new_new_n847_), .B(new_new_n491_), .Y(new_new_n852_));
  NO3        g830(.A(new_new_n389_), .B(new_new_n351_), .C(new_new_n347_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n249_), .B(new_new_n304_), .Y(new_new_n854_));
  INV        g832(.A(new_new_n683_), .Y(new_new_n855_));
  AOI210     g833(.A0(new_new_n855_), .A1(new_new_n854_), .B0(new_new_n853_), .Y(new_new_n856_));
  NA4        g834(.A(new_new_n856_), .B(new_new_n852_), .C(new_new_n849_), .D(new_new_n843_), .Y(new_new_n857_));
  NO2        g835(.A(new_new_n808_), .B(new_new_n235_), .Y(new_new_n858_));
  AN2        g836(.A(new_new_n318_), .B(new_new_n315_), .Y(new_new_n859_));
  AN2        g837(.A(new_new_n859_), .B(new_new_n804_), .Y(new_new_n860_));
  OAI210     g838(.A0(new_new_n860_), .A1(new_new_n858_), .B0(i_10_), .Y(new_new_n861_));
  OA210      g839(.A0(new_new_n454_), .A1(new_new_n220_), .B0(new_new_n453_), .Y(new_new_n862_));
  NA3        g840(.A(new_new_n453_), .B(new_new_n397_), .C(new_new_n46_), .Y(new_new_n863_));
  OAI210     g841(.A0(new_new_n812_), .A1(i_6_), .B0(new_new_n863_), .Y(new_new_n864_));
  NO2        g842(.A(new_new_n247_), .B(new_new_n47_), .Y(new_new_n865_));
  NO2        g843(.A(new_new_n865_), .B(new_new_n183_), .Y(new_new_n866_));
  AOI220     g844(.A0(new_new_n866_), .A1(new_new_n454_), .B0(new_new_n864_), .B1(new_new_n70_), .Y(new_new_n867_));
  NA3        g845(.A(new_new_n760_), .B(new_new_n369_), .C(new_new_n609_), .Y(new_new_n868_));
  NA2        g846(.A(new_new_n88_), .B(new_new_n45_), .Y(new_new_n869_));
  NO2        g847(.A(new_new_n72_), .B(new_new_n704_), .Y(new_new_n870_));
  AOI220     g848(.A0(new_new_n870_), .A1(new_new_n869_), .B0(new_new_n170_), .B1(new_new_n572_), .Y(new_new_n871_));
  AOI210     g849(.A0(new_new_n871_), .A1(new_new_n868_), .B0(new_new_n48_), .Y(new_new_n872_));
  NO3        g850(.A(new_new_n564_), .B(new_new_n346_), .C(new_new_n24_), .Y(new_new_n873_));
  AOI210     g851(.A0(new_new_n661_), .A1(new_new_n524_), .B0(new_new_n873_), .Y(new_new_n874_));
  NO2        g852(.A(new_new_n575_), .B(new_new_n101_), .Y(new_new_n875_));
  NA2        g853(.A(new_new_n875_), .B(i_0_), .Y(new_new_n876_));
  OAI220     g854(.A0(new_new_n876_), .A1(new_new_n82_), .B0(new_new_n874_), .B1(new_new_n169_), .Y(new_new_n877_));
  NO3        g855(.A(new_new_n877_), .B(new_new_n872_), .C(new_new_n495_), .Y(new_new_n878_));
  NA3        g856(.A(new_new_n878_), .B(new_new_n867_), .C(new_new_n861_), .Y(new_new_n879_));
  NO3        g857(.A(new_new_n879_), .B(new_new_n857_), .C(new_new_n830_), .Y(new_new_n880_));
  NO2        g858(.A(i_0_), .B(new_new_n683_), .Y(new_new_n881_));
  NO3        g859(.A(new_new_n101_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n882_));
  AO220      g860(.A0(new_new_n882_), .A1(new_new_n70_), .B0(new_new_n881_), .B1(new_new_n170_), .Y(new_new_n883_));
  NA2        g861(.A(new_new_n883_), .B(new_new_n336_), .Y(new_new_n884_));
  NA2        g862(.A(new_new_n690_), .B(new_new_n143_), .Y(new_new_n885_));
  INV        g863(.A(new_new_n885_), .Y(new_new_n886_));
  NA2        g864(.A(new_new_n886_), .B(new_new_n640_), .Y(new_new_n887_));
  NO2        g865(.A(new_new_n756_), .B(new_new_n389_), .Y(new_new_n888_));
  NA2        g866(.A(new_new_n782_), .B(new_new_n49_), .Y(new_new_n889_));
  NA2        g867(.A(new_new_n783_), .B(i_9_), .Y(new_new_n890_));
  NO2        g868(.A(new_new_n889_), .B(new_new_n890_), .Y(new_new_n891_));
  NA2        g869(.A(new_new_n239_), .B(new_new_n227_), .Y(new_new_n892_));
  AOI210     g870(.A0(new_new_n892_), .A1(new_new_n817_), .B0(new_new_n150_), .Y(new_new_n893_));
  NO3        g871(.A(new_new_n893_), .B(new_new_n891_), .C(new_new_n888_), .Y(new_new_n894_));
  NA3        g872(.A(new_new_n894_), .B(new_new_n887_), .C(new_new_n884_), .Y(new_new_n895_));
  NA2        g873(.A(new_new_n859_), .B(new_new_n359_), .Y(new_new_n896_));
  AOI210     g874(.A0(new_new_n288_), .A1(new_new_n159_), .B0(new_new_n896_), .Y(new_new_n897_));
  NA2        g875(.A(new_new_n40_), .B(new_new_n45_), .Y(new_new_n898_));
  NA2        g876(.A(new_new_n835_), .B(new_new_n467_), .Y(new_new_n899_));
  AOI210     g877(.A0(new_new_n898_), .A1(new_new_n159_), .B0(new_new_n899_), .Y(new_new_n900_));
  NO2        g878(.A(new_new_n900_), .B(new_new_n897_), .Y(new_new_n901_));
  NO3        g879(.A(new_new_n824_), .B(new_new_n800_), .C(new_new_n186_), .Y(new_new_n902_));
  AOI220     g880(.A0(new_new_n902_), .A1(i_11_), .B0(new_new_n545_), .B1(new_new_n72_), .Y(new_new_n903_));
  NO3        g881(.A(new_new_n205_), .B(new_new_n370_), .C(i_0_), .Y(new_new_n904_));
  OAI210     g882(.A0(new_new_n904_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n905_));
  INV        g883(.A(new_new_n214_), .Y(new_new_n906_));
  OAI220     g884(.A0(new_new_n507_), .A1(new_new_n136_), .B0(new_new_n613_), .B1(new_new_n589_), .Y(new_new_n907_));
  NA3        g885(.A(new_new_n907_), .B(i_7_), .C(new_new_n906_), .Y(new_new_n908_));
  NA4        g886(.A(new_new_n908_), .B(new_new_n905_), .C(new_new_n903_), .D(new_new_n901_), .Y(new_new_n909_));
  NO2        g887(.A(new_new_n237_), .B(new_new_n88_), .Y(new_new_n910_));
  AOI210     g888(.A0(new_new_n910_), .A1(new_new_n881_), .B0(new_new_n105_), .Y(new_new_n911_));
  AOI220     g889(.A0(new_new_n850_), .A1(new_new_n467_), .B0(new_new_n782_), .B1(new_new_n160_), .Y(new_new_n912_));
  NA2        g890(.A(new_new_n339_), .B(new_new_n172_), .Y(new_new_n913_));
  OA220      g891(.A0(new_new_n913_), .A1(new_new_n912_), .B0(new_new_n911_), .B1(i_5_), .Y(new_new_n914_));
  AOI210     g892(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n171_), .Y(new_new_n915_));
  NA2        g893(.A(new_new_n915_), .B(new_new_n862_), .Y(new_new_n916_));
  NA3        g894(.A(new_new_n586_), .B(new_new_n181_), .C(new_new_n80_), .Y(new_new_n917_));
  NA2        g895(.A(new_new_n917_), .B(new_new_n522_), .Y(new_new_n918_));
  INV        g896(.A(new_new_n465_), .Y(new_new_n919_));
  NO2        g897(.A(new_new_n919_), .B(new_new_n918_), .Y(new_new_n920_));
  NA3        g898(.A(new_new_n377_), .B(new_new_n320_), .C(new_new_n218_), .Y(new_new_n921_));
  NA4        g899(.A(new_new_n921_), .B(new_new_n920_), .C(new_new_n916_), .D(new_new_n914_), .Y(new_new_n922_));
  INV        g900(.A(new_new_n588_), .Y(new_new_n923_));
  NO3        g901(.A(new_new_n923_), .B(new_new_n535_), .C(new_new_n333_), .Y(new_new_n924_));
  NO2        g902(.A(new_new_n82_), .B(i_5_), .Y(new_new_n925_));
  NA3        g903(.A(new_new_n783_), .B(new_new_n106_), .C(new_new_n121_), .Y(new_new_n926_));
  INV        g904(.A(new_new_n926_), .Y(new_new_n927_));
  AOI210     g905(.A0(new_new_n927_), .A1(new_new_n925_), .B0(new_new_n924_), .Y(new_new_n928_));
  NA3        g906(.A(new_new_n293_), .B(i_5_), .C(new_new_n189_), .Y(new_new_n929_));
  NAi31      g907(.An(new_new_n236_), .B(new_new_n929_), .C(new_new_n237_), .Y(new_new_n930_));
  NO4        g908(.A(new_new_n235_), .B(new_new_n205_), .C(i_0_), .D(i_12_), .Y(new_new_n931_));
  NA2        g909(.A(new_new_n931_), .B(new_new_n930_), .Y(new_new_n932_));
  AN2        g910(.A(new_new_n824_), .B(new_new_n150_), .Y(new_new_n933_));
  NO4        g911(.A(new_new_n933_), .B(i_12_), .C(new_new_n617_), .D(new_new_n128_), .Y(new_new_n934_));
  NA2        g912(.A(new_new_n934_), .B(new_new_n214_), .Y(new_new_n935_));
  NA3        g913(.A(new_new_n94_), .B(new_new_n549_), .C(i_11_), .Y(new_new_n936_));
  NO2        g914(.A(new_new_n936_), .B(new_new_n152_), .Y(new_new_n937_));
  NA2        g915(.A(new_new_n850_), .B(new_new_n451_), .Y(new_new_n938_));
  OAI220     g916(.A0(i_7_), .A1(new_new_n929_), .B0(new_new_n938_), .B1(new_new_n641_), .Y(new_new_n939_));
  AOI210     g917(.A0(new_new_n939_), .A1(new_new_n838_), .B0(new_new_n937_), .Y(new_new_n940_));
  NA4        g918(.A(new_new_n940_), .B(new_new_n935_), .C(new_new_n932_), .D(new_new_n928_), .Y(new_new_n941_));
  NO4        g919(.A(new_new_n941_), .B(new_new_n922_), .C(new_new_n909_), .D(new_new_n895_), .Y(new_new_n942_));
  OAI210     g920(.A0(new_new_n759_), .A1(new_new_n752_), .B0(new_new_n37_), .Y(new_new_n943_));
  NA3        g921(.A(new_new_n846_), .B(new_new_n354_), .C(i_5_), .Y(new_new_n944_));
  NA3        g922(.A(new_new_n944_), .B(new_new_n943_), .C(new_new_n584_), .Y(new_new_n945_));
  NA2        g923(.A(new_new_n945_), .B(new_new_n201_), .Y(new_new_n946_));
  BUFFER     g924(.A(new_new_n355_), .Y(new_new_n947_));
  NA2        g925(.A(new_new_n182_), .B(new_new_n184_), .Y(new_new_n948_));
  AO210      g926(.A0(new_new_n947_), .A1(new_new_n33_), .B0(new_new_n948_), .Y(new_new_n949_));
  OAI210     g927(.A0(new_new_n588_), .A1(new_new_n586_), .B0(new_new_n303_), .Y(new_new_n950_));
  INV        g928(.A(new_new_n614_), .Y(new_new_n951_));
  NA3        g929(.A(new_new_n951_), .B(new_new_n950_), .C(new_new_n949_), .Y(new_new_n952_));
  NO2        g930(.A(new_new_n443_), .B(new_new_n255_), .Y(new_new_n953_));
  NO4        g931(.A(new_new_n230_), .B(new_new_n142_), .C(new_new_n642_), .D(new_new_n37_), .Y(new_new_n954_));
  NO2        g932(.A(new_new_n954_), .B(new_new_n953_), .Y(new_new_n955_));
  OAI210     g933(.A0(new_new_n936_), .A1(new_new_n145_), .B0(new_new_n955_), .Y(new_new_n956_));
  AOI210     g934(.A0(new_new_n952_), .A1(new_new_n49_), .B0(new_new_n956_), .Y(new_new_n957_));
  AOI210     g935(.A0(new_new_n957_), .A1(new_new_n946_), .B0(new_new_n70_), .Y(new_new_n958_));
  NO2        g936(.A(new_new_n542_), .B(new_new_n366_), .Y(new_new_n959_));
  NO2        g937(.A(new_new_n959_), .B(new_new_n710_), .Y(new_new_n960_));
  OAI210     g938(.A0(new_new_n77_), .A1(new_new_n55_), .B0(new_new_n104_), .Y(new_new_n961_));
  NA2        g939(.A(new_new_n961_), .B(new_new_n73_), .Y(new_new_n962_));
  AOI210     g940(.A0(new_new_n915_), .A1(new_new_n835_), .B0(new_new_n851_), .Y(new_new_n963_));
  AOI210     g941(.A0(new_new_n963_), .A1(new_new_n962_), .B0(new_new_n642_), .Y(new_new_n964_));
  NA2        g942(.A(new_new_n249_), .B(new_new_n58_), .Y(new_new_n965_));
  AOI220     g943(.A0(new_new_n965_), .A1(new_new_n73_), .B0(new_new_n334_), .B1(new_new_n246_), .Y(new_new_n966_));
  NO2        g944(.A(new_new_n966_), .B(new_new_n233_), .Y(new_new_n967_));
  NA3        g945(.A(new_new_n92_), .B(new_new_n295_), .C(new_new_n31_), .Y(new_new_n968_));
  INV        g946(.A(new_new_n968_), .Y(new_new_n969_));
  NO3        g947(.A(new_new_n969_), .B(new_new_n967_), .C(new_new_n964_), .Y(new_new_n970_));
  OAI210     g948(.A0(new_new_n257_), .A1(new_new_n155_), .B0(new_new_n83_), .Y(new_new_n971_));
  NA3        g949(.A(new_new_n713_), .B(new_new_n277_), .C(new_new_n77_), .Y(new_new_n972_));
  AOI210     g950(.A0(new_new_n972_), .A1(new_new_n971_), .B0(i_11_), .Y(new_new_n973_));
  NA2        g951(.A(new_new_n581_), .B(new_new_n211_), .Y(new_new_n974_));
  OAI210     g952(.A0(new_new_n974_), .A1(new_new_n846_), .B0(new_new_n201_), .Y(new_new_n975_));
  NA2        g953(.A(new_new_n161_), .B(i_5_), .Y(new_new_n976_));
  NO2        g954(.A(new_new_n975_), .B(new_new_n976_), .Y(new_new_n977_));
  NO3        g955(.A(new_new_n60_), .B(new_new_n59_), .C(i_4_), .Y(new_new_n978_));
  OAI210     g956(.A0(new_new_n854_), .A1(new_new_n295_), .B0(new_new_n978_), .Y(new_new_n979_));
  NO2        g957(.A(new_new_n979_), .B(new_new_n683_), .Y(new_new_n980_));
  NO3        g958(.A(new_new_n980_), .B(new_new_n977_), .C(new_new_n973_), .Y(new_new_n981_));
  OAI210     g959(.A0(new_new_n970_), .A1(i_4_), .B0(new_new_n981_), .Y(new_new_n982_));
  NO3        g960(.A(new_new_n982_), .B(new_new_n960_), .C(new_new_n958_), .Y(new_new_n983_));
  NA4        g961(.A(new_new_n983_), .B(new_new_n942_), .C(new_new_n880_), .D(new_new_n807_), .Y(men4));
  INV        g962(.A(i_2_), .Y(new_new_n987_));
  INV        g963(.A(new_new_n315_), .Y(new_new_n988_));
  INV        g964(.A(i_1_), .Y(new_new_n989_));
  INV        g965(.A(new_new_n721_), .Y(new_new_n990_));
  INV        g966(.A(new_new_n293_), .Y(new_new_n991_));
  INV        g967(.A(i_0_), .Y(new_new_n992_));
  INV        g968(.A(i_3_), .Y(new_new_n993_));
endmodule


