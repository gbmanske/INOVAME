//Benchmark atmr_alu4_1266_0.25

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n106_, ori_ori_n107_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n128_, mai_mai_n129_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NAi31      o017(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n35_), .Y(ori1));
  INV        o019(.A(i_11_), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(i_6_), .Y(ori_ori_n43_));
  INV        o021(.A(i_2_), .Y(ori_ori_n44_));
  INV        o022(.A(i_5_), .Y(ori_ori_n45_));
  NO2        o023(.A(i_7_), .B(i_10_), .Y(ori_ori_n46_));
  AOI210     o024(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n46_), .Y(ori_ori_n47_));
  NO2        o025(.A(i_5_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NA2        o026(.A(i_7_), .B(i_9_), .Y(ori_ori_n49_));
  NA2        o027(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n50_));
  NO2        o028(.A(i_1_), .B(i_6_), .Y(ori_ori_n51_));
  NAi21      o029(.An(i_2_), .B(i_7_), .Y(ori_ori_n52_));
  INV        o030(.A(i_1_), .Y(ori_ori_n53_));
  NA3        o031(.A(ori_ori_n327_), .B(ori_ori_n52_), .C(ori_ori_n31_), .Y(ori_ori_n54_));
  NA2        o032(.A(i_1_), .B(i_10_), .Y(ori_ori_n55_));
  INV        o033(.A(ori_ori_n55_), .Y(ori_ori_n56_));
  NAi21      o034(.An(ori_ori_n56_), .B(ori_ori_n54_), .Y(ori_ori_n57_));
  NA2        o035(.A(ori_ori_n47_), .B(i_2_), .Y(ori_ori_n58_));
  AOI210     o036(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n59_));
  NA2        o037(.A(i_1_), .B(i_6_), .Y(ori_ori_n60_));
  NO2        o038(.A(ori_ori_n60_), .B(ori_ori_n25_), .Y(ori_ori_n61_));
  INV        o039(.A(i_0_), .Y(ori_ori_n62_));
  NAi21      o040(.An(i_5_), .B(i_10_), .Y(ori_ori_n63_));
  NA2        o041(.A(i_5_), .B(i_9_), .Y(ori_ori_n64_));
  AOI210     o042(.A0(ori_ori_n64_), .A1(ori_ori_n63_), .B0(ori_ori_n62_), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n65_), .B(ori_ori_n61_), .Y(ori_ori_n66_));
  INV        o044(.A(ori_ori_n66_), .Y(ori_ori_n67_));
  OAI210     o045(.A0(ori_ori_n67_), .A1(ori_ori_n57_), .B0(i_0_), .Y(ori_ori_n68_));
  NA2        o046(.A(i_12_), .B(i_5_), .Y(ori_ori_n69_));
  INV        o047(.A(i_6_), .Y(ori_ori_n70_));
  NO2        o048(.A(i_2_), .B(i_7_), .Y(ori_ori_n71_));
  INV        o049(.A(ori_ori_n71_), .Y(ori_ori_n72_));
  NA2        o050(.A(i_1_), .B(ori_ori_n72_), .Y(ori_ori_n73_));
  NAi21      o051(.An(i_6_), .B(i_10_), .Y(ori_ori_n74_));
  NA2        o052(.A(i_6_), .B(i_9_), .Y(ori_ori_n75_));
  AOI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n53_), .Y(ori_ori_n76_));
  NA2        o054(.A(i_2_), .B(i_6_), .Y(ori_ori_n77_));
  INV        o055(.A(ori_ori_n76_), .Y(ori_ori_n78_));
  AOI210     o056(.A0(ori_ori_n78_), .A1(ori_ori_n73_), .B0(ori_ori_n69_), .Y(ori_ori_n79_));
  AN3        o057(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n80_));
  NAi21      o058(.An(i_6_), .B(i_11_), .Y(ori_ori_n81_));
  NA2        o059(.A(ori_ori_n80_), .B(ori_ori_n32_), .Y(ori_ori_n82_));
  INV        o060(.A(i_7_), .Y(ori_ori_n83_));
  NA2        o061(.A(ori_ori_n44_), .B(ori_ori_n83_), .Y(ori_ori_n84_));
  NO2        o062(.A(i_0_), .B(i_5_), .Y(ori_ori_n85_));
  NO2        o063(.A(ori_ori_n85_), .B(ori_ori_n70_), .Y(ori_ori_n86_));
  NA3        o064(.A(i_12_), .B(ori_ori_n86_), .C(ori_ori_n84_), .Y(ori_ori_n87_));
  INV        o065(.A(i_7_), .Y(ori_ori_n88_));
  OR2        o066(.A(ori_ori_n69_), .B(ori_ori_n51_), .Y(ori_ori_n89_));
  NA2        o067(.A(i_12_), .B(i_7_), .Y(ori_ori_n90_));
  NA2        o068(.A(i_11_), .B(i_12_), .Y(ori_ori_n91_));
  NA3        o069(.A(ori_ori_n91_), .B(ori_ori_n87_), .C(ori_ori_n82_), .Y(ori_ori_n92_));
  NOi21      o070(.An(i_1_), .B(i_5_), .Y(ori_ori_n93_));
  NA2        o071(.A(ori_ori_n93_), .B(i_11_), .Y(ori_ori_n94_));
  NA2        o072(.A(ori_ori_n83_), .B(ori_ori_n37_), .Y(ori_ori_n95_));
  NA2        o073(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n96_));
  NA2        o074(.A(ori_ori_n96_), .B(ori_ori_n95_), .Y(ori_ori_n97_));
  NO2        o075(.A(ori_ori_n97_), .B(ori_ori_n44_), .Y(ori_ori_n98_));
  NA2        o076(.A(ori_ori_n75_), .B(ori_ori_n74_), .Y(ori_ori_n99_));
  INV        o077(.A(ori_ori_n52_), .Y(ori_ori_n100_));
  NOi21      o078(.An(ori_ori_n100_), .B(ori_ori_n99_), .Y(ori_ori_n101_));
  NO2        o079(.A(i_1_), .B(ori_ori_n70_), .Y(ori_ori_n102_));
  NO2        o080(.A(ori_ori_n101_), .B(ori_ori_n94_), .Y(ori_ori_n103_));
  NO3        o081(.A(ori_ori_n103_), .B(ori_ori_n92_), .C(ori_ori_n79_), .Y(ori_ori_n104_));
  NA3        o082(.A(ori_ori_n104_), .B(ori_ori_n68_), .C(ori_ori_n50_), .Y(ori2));
  NO2        o083(.A(ori_ori_n53_), .B(ori_ori_n37_), .Y(ori_ori_n106_));
  NA2        o084(.A(ori_ori_n325_), .B(ori_ori_n106_), .Y(ori_ori_n107_));
  NA4        o085(.A(ori_ori_n107_), .B(ori_ori_n66_), .C(ori_ori_n58_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o086(.A(i_0_), .B(i_1_), .Y(ori_ori_n109_));
  NA2        o087(.A(i_2_), .B(i_3_), .Y(ori_ori_n110_));
  NO2        o088(.A(ori_ori_n110_), .B(i_4_), .Y(ori_ori_n111_));
  NA2        o089(.A(i_1_), .B(i_5_), .Y(ori_ori_n112_));
  NOi21      o090(.An(i_4_), .B(i_10_), .Y(ori_ori_n113_));
  NOi21      o091(.An(i_4_), .B(i_9_), .Y(ori_ori_n114_));
  NOi21      o092(.An(i_11_), .B(i_13_), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n62_), .B(ori_ori_n53_), .Y(ori_ori_n116_));
  NAi21      o094(.An(i_4_), .B(i_12_), .Y(ori_ori_n117_));
  INV        o095(.A(i_8_), .Y(ori_ori_n118_));
  NO3        o096(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n119_));
  NO2        o097(.A(i_13_), .B(i_9_), .Y(ori_ori_n120_));
  NAi21      o098(.An(i_12_), .B(i_3_), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n42_), .B(i_5_), .Y(ori_ori_n122_));
  INV        o100(.A(i_13_), .Y(ori_ori_n123_));
  NO2        o101(.A(i_12_), .B(ori_ori_n123_), .Y(ori_ori_n124_));
  NO2        o102(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n125_));
  INV        o103(.A(i_12_), .Y(ori_ori_n126_));
  NO3        o104(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n127_));
  NAi21      o105(.An(i_4_), .B(i_3_), .Y(ori_ori_n128_));
  INV        o106(.A(i_0_), .Y(ori_ori_n129_));
  NO2        o107(.A(i_11_), .B(ori_ori_n123_), .Y(ori_ori_n130_));
  NA2        o108(.A(i_12_), .B(i_6_), .Y(ori_ori_n131_));
  OR2        o109(.A(i_13_), .B(i_9_), .Y(ori_ori_n132_));
  NO2        o110(.A(ori_ori_n128_), .B(i_2_), .Y(ori_ori_n133_));
  NO2        o111(.A(i_2_), .B(ori_ori_n83_), .Y(ori_ori_n134_));
  AN2        o112(.A(i_3_), .B(i_10_), .Y(ori_ori_n135_));
  NO2        o113(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n136_));
  NO2        o114(.A(ori_ori_n44_), .B(ori_ori_n26_), .Y(ori_ori_n137_));
  NO2        o115(.A(i_2_), .B(i_3_), .Y(ori_ori_n138_));
  NO2        o116(.A(i_12_), .B(i_10_), .Y(ori_ori_n139_));
  NOi21      o117(.An(i_5_), .B(i_0_), .Y(ori_ori_n140_));
  NAi21      o118(.An(i_3_), .B(i_4_), .Y(ori_ori_n141_));
  AN2        o119(.A(i_12_), .B(i_5_), .Y(ori_ori_n142_));
  NO2        o120(.A(i_5_), .B(i_10_), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n144_));
  NO3        o122(.A(ori_ori_n70_), .B(ori_ori_n45_), .C(i_9_), .Y(ori_ori_n145_));
  NO2        o123(.A(i_0_), .B(i_11_), .Y(ori_ori_n146_));
  NOi21      o124(.An(i_2_), .B(i_12_), .Y(ori_ori_n147_));
  NAi21      o125(.An(i_9_), .B(i_4_), .Y(ori_ori_n148_));
  OR2        o126(.A(i_13_), .B(i_10_), .Y(ori_ori_n149_));
  NO3        o127(.A(ori_ori_n149_), .B(ori_ori_n91_), .C(ori_ori_n148_), .Y(ori_ori_n150_));
  NO2        o128(.A(ori_ori_n83_), .B(ori_ori_n25_), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n62_), .B(i_13_), .Y(ori_ori_n152_));
  NO2        o130(.A(i_10_), .B(i_9_), .Y(ori_ori_n153_));
  NO3        o131(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n154_));
  NA2        o132(.A(ori_ori_n131_), .B(ori_ori_n81_), .Y(ori_ori_n155_));
  NA2        o133(.A(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n130_), .B(ori_ori_n136_), .Y(ori_ori_n157_));
  NO3        o135(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n158_));
  INV        o136(.A(ori_ori_n158_), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n159_), .B(ori_ori_n157_), .Y(ori_ori_n160_));
  INV        o138(.A(ori_ori_n160_), .Y(ori_ori_n161_));
  NO2        o139(.A(i_11_), .B(i_1_), .Y(ori_ori_n162_));
  NA3        o140(.A(ori_ori_n144_), .B(ori_ori_n116_), .C(ori_ori_n111_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n154_), .B(ori_ori_n142_), .Y(ori_ori_n164_));
  NA2        o142(.A(ori_ori_n158_), .B(ori_ori_n143_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n163_), .B(ori_ori_n161_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n167_));
  AOI210     o145(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n150_), .Y(ori_ori_n168_));
  INV        o146(.A(ori_ori_n168_), .Y(ori_ori_n169_));
  NO3        o147(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n170_));
  NO2        o148(.A(ori_ori_n149_), .B(i_1_), .Y(ori_ori_n171_));
  NOi31      o149(.An(ori_ori_n171_), .B(ori_ori_n155_), .C(ori_ori_n62_), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n90_), .B(ori_ori_n23_), .Y(ori_ori_n173_));
  NO2        o151(.A(i_12_), .B(ori_ori_n70_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n169_), .B(ori_ori_n166_), .Y(ori_ori_n175_));
  INV        o153(.A(ori_ori_n175_), .Y(ori7));
  NO2        o154(.A(ori_ori_n77_), .B(ori_ori_n49_), .Y(ori_ori_n177_));
  NA2        o155(.A(i_11_), .B(ori_ori_n118_), .Y(ori_ori_n178_));
  NA2        o156(.A(i_2_), .B(ori_ori_n70_), .Y(ori_ori_n179_));
  NA2        o157(.A(ori_ori_n71_), .B(ori_ori_n119_), .Y(ori_ori_n180_));
  NO2        o158(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n135_), .B(ori_ori_n181_), .Y(ori_ori_n182_));
  OAI220     o160(.A0(ori_ori_n182_), .A1(ori_ori_n179_), .B0(ori_ori_n180_), .B1(i_13_), .Y(ori_ori_n183_));
  NO2        o161(.A(ori_ori_n183_), .B(ori_ori_n177_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n52_), .B(i_10_), .Y(ori_ori_n185_));
  AOI210     o163(.A0(ori_ori_n185_), .A1(ori_ori_n126_), .B0(ori_ori_n113_), .Y(ori_ori_n186_));
  OR2        o164(.A(ori_ori_n186_), .B(ori_ori_n132_), .Y(ori_ori_n187_));
  AOI210     o165(.A0(ori_ori_n187_), .A1(ori_ori_n184_), .B0(ori_ori_n53_), .Y(ori_ori_n188_));
  NOi21      o166(.An(i_11_), .B(i_7_), .Y(ori_ori_n189_));
  AO210      o167(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n190_));
  NO2        o168(.A(ori_ori_n190_), .B(ori_ori_n189_), .Y(ori_ori_n191_));
  NA2        o169(.A(ori_ori_n124_), .B(ori_ori_n53_), .Y(ori_ori_n192_));
  NO2        o170(.A(i_1_), .B(i_12_), .Y(ori_ori_n193_));
  INV        o171(.A(ori_ori_n192_), .Y(ori_ori_n194_));
  NA2        o172(.A(ori_ori_n194_), .B(i_6_), .Y(ori_ori_n195_));
  NO2        o173(.A(i_6_), .B(i_11_), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n156_), .Y(ori_ori_n197_));
  INV        o175(.A(i_2_), .Y(ori_ori_n198_));
  NA2        o176(.A(ori_ori_n106_), .B(i_9_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n199_), .B(ori_ori_n198_), .Y(ori_ori_n200_));
  AOI210     o178(.A0(ori_ori_n162_), .A1(ori_ori_n151_), .B0(ori_ori_n127_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n201_), .B(ori_ori_n179_), .Y(ori_ori_n202_));
  NO2        o180(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n203_));
  OR2        o181(.A(ori_ori_n202_), .B(ori_ori_n200_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n204_), .B(ori_ori_n197_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n126_), .B(ori_ori_n83_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n206_), .B(ori_ori_n189_), .Y(ori_ori_n207_));
  NO2        o185(.A(i_7_), .B(ori_ori_n42_), .Y(ori_ori_n208_));
  NO3        o186(.A(ori_ori_n208_), .B(ori_ori_n137_), .C(i_12_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n91_), .B(ori_ori_n37_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n210_), .B(i_6_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n70_), .B(i_9_), .Y(ori_ori_n212_));
  NO2        o190(.A(ori_ori_n212_), .B(ori_ori_n53_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n213_), .B(ori_ori_n193_), .Y(ori_ori_n214_));
  NO4        o192(.A(ori_ori_n214_), .B(ori_ori_n211_), .C(ori_ori_n209_), .D(i_4_), .Y(ori_ori_n215_));
  INV        o193(.A(ori_ori_n215_), .Y(ori_ori_n216_));
  NA3        o194(.A(ori_ori_n216_), .B(ori_ori_n205_), .C(ori_ori_n195_), .Y(ori_ori_n217_));
  AOI210     o195(.A0(ori_ori_n131_), .A1(ori_ori_n81_), .B0(i_1_), .Y(ori_ori_n218_));
  NO2        o196(.A(ori_ori_n141_), .B(i_2_), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n219_), .B(ori_ori_n218_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n220_), .B(i_13_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n49_), .B(i_12_), .Y(ori_ori_n222_));
  INV        o200(.A(ori_ori_n222_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n223_), .B(ori_ori_n77_), .Y(ori_ori_n224_));
  INV        o202(.A(ori_ori_n224_), .Y(ori_ori_n225_));
  NA2        o203(.A(ori_ori_n99_), .B(i_13_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n226_), .B(ori_ori_n218_), .Y(ori_ori_n227_));
  INV        o205(.A(ori_ori_n227_), .Y(ori_ori_n228_));
  OR2        o206(.A(i_11_), .B(i_6_), .Y(ori_ori_n229_));
  NA3        o207(.A(ori_ori_n147_), .B(ori_ori_n181_), .C(ori_ori_n81_), .Y(ori_ori_n230_));
  NA2        o208(.A(ori_ori_n196_), .B(i_13_), .Y(ori_ori_n231_));
  NA2        o209(.A(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NA2        o210(.A(ori_ori_n232_), .B(ori_ori_n53_), .Y(ori_ori_n233_));
  NA3        o211(.A(ori_ori_n233_), .B(ori_ori_n228_), .C(ori_ori_n225_), .Y(ori_ori_n234_));
  OR4        o212(.A(ori_ori_n234_), .B(ori_ori_n221_), .C(ori_ori_n217_), .D(ori_ori_n188_), .Y(ori5));
  NA2        o213(.A(ori_ori_n207_), .B(ori_ori_n133_), .Y(ori_ori_n236_));
  INV        o214(.A(ori_ori_n236_), .Y(ori_ori_n237_));
  NO2        o215(.A(ori_ori_n96_), .B(ori_ori_n23_), .Y(ori_ori_n238_));
  INV        o216(.A(ori_ori_n153_), .Y(ori_ori_n239_));
  AOI220     o217(.A0(ori_ori_n138_), .A1(ori_ori_n173_), .B0(i_12_), .B1(ori_ori_n238_), .Y(ori_ori_n240_));
  INV        o218(.A(ori_ori_n240_), .Y(ori_ori_n241_));
  NO2        o219(.A(ori_ori_n241_), .B(ori_ori_n237_), .Y(ori_ori_n242_));
  INV        o220(.A(ori_ori_n115_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n219_), .B(ori_ori_n88_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n244_), .B(ori_ori_n243_), .Y(ori_ori_n245_));
  INV        o223(.A(ori_ori_n151_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n246_), .B(i_2_), .Y(ori_ori_n247_));
  INV        o225(.A(ori_ori_n247_), .Y(ori_ori_n248_));
  AOI210     o226(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n149_), .Y(ori_ori_n249_));
  AOI210     o227(.A0(ori_ori_n249_), .A1(ori_ori_n248_), .B0(ori_ori_n245_), .Y(ori_ori_n250_));
  NO2        o228(.A(ori_ori_n117_), .B(ori_ori_n97_), .Y(ori_ori_n251_));
  OAI210     o229(.A0(ori_ori_n251_), .A1(ori_ori_n238_), .B0(i_2_), .Y(ori_ori_n252_));
  NO2        o230(.A(ori_ori_n252_), .B(ori_ori_n118_), .Y(ori_ori_n253_));
  OA210      o231(.A0(ori_ori_n191_), .A1(ori_ori_n98_), .B0(i_13_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n121_), .A1(ori_ori_n110_), .B0(ori_ori_n167_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n255_), .B(ori_ori_n151_), .Y(ori_ori_n256_));
  NO2        o234(.A(ori_ori_n84_), .B(ori_ori_n42_), .Y(ori_ori_n257_));
  INV        o235(.A(ori_ori_n134_), .Y(ori_ori_n258_));
  NA4        o236(.A(ori_ori_n258_), .B(ori_ori_n135_), .C(ori_ori_n96_), .D(ori_ori_n40_), .Y(ori_ori_n259_));
  OAI210     o237(.A0(ori_ori_n259_), .A1(ori_ori_n257_), .B0(ori_ori_n256_), .Y(ori_ori_n260_));
  NO3        o238(.A(ori_ori_n260_), .B(ori_ori_n254_), .C(ori_ori_n253_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n52_), .B(i_12_), .Y(ori_ori_n262_));
  NO2        o240(.A(ori_ori_n262_), .B(ori_ori_n98_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n263_), .B(ori_ori_n178_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n264_), .B(ori_ori_n36_), .Y(ori_ori_n265_));
  NA4        o243(.A(ori_ori_n265_), .B(ori_ori_n261_), .C(ori_ori_n250_), .D(ori_ori_n242_), .Y(ori6));
  INV        o244(.A(ori_ori_n140_), .Y(ori_ori_n267_));
  OR2        o245(.A(ori_ori_n267_), .B(i_12_), .Y(ori_ori_n268_));
  NA2        o246(.A(ori_ori_n174_), .B(ori_ori_n53_), .Y(ori_ori_n269_));
  INV        o247(.A(ori_ori_n269_), .Y(ori_ori_n270_));
  NA2        o248(.A(ori_ori_n270_), .B(ori_ori_n62_), .Y(ori_ori_n271_));
  INV        o249(.A(ori_ori_n139_), .Y(ori_ori_n272_));
  NA2        o250(.A(ori_ori_n64_), .B(ori_ori_n102_), .Y(ori_ori_n273_));
  INV        o251(.A(ori_ori_n96_), .Y(ori_ori_n274_));
  NA2        o252(.A(ori_ori_n274_), .B(ori_ori_n44_), .Y(ori_ori_n275_));
  AOI210     o253(.A0(ori_ori_n275_), .A1(ori_ori_n273_), .B0(ori_ori_n272_), .Y(ori_ori_n276_));
  NAi32      o254(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n277_));
  NO2        o255(.A(ori_ori_n229_), .B(ori_ori_n277_), .Y(ori_ori_n278_));
  OR2        o256(.A(ori_ori_n278_), .B(ori_ori_n276_), .Y(ori_ori_n279_));
  BUFFER     o257(.A(ori_ori_n191_), .Y(ori_ori_n280_));
  NA2        o258(.A(ori_ori_n280_), .B(ori_ori_n109_), .Y(ori_ori_n281_));
  AO210      o259(.A0(ori_ori_n165_), .A1(ori_ori_n239_), .B0(ori_ori_n36_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n282_), .B(ori_ori_n281_), .Y(ori_ori_n283_));
  NO2        o261(.A(i_6_), .B(i_11_), .Y(ori_ori_n284_));
  NA2        o262(.A(ori_ori_n284_), .B(ori_ori_n170_), .Y(ori_ori_n285_));
  NA2        o263(.A(ori_ori_n145_), .B(ori_ori_n59_), .Y(ori_ori_n286_));
  NA3        o264(.A(ori_ori_n286_), .B(ori_ori_n285_), .C(ori_ori_n180_), .Y(ori_ori_n287_));
  NA2        o265(.A(ori_ori_n89_), .B(ori_ori_n146_), .Y(ori_ori_n288_));
  INV        o266(.A(ori_ori_n288_), .Y(ori_ori_n289_));
  NO4        o267(.A(ori_ori_n289_), .B(ori_ori_n287_), .C(ori_ori_n283_), .D(ori_ori_n279_), .Y(ori_ori_n290_));
  NA3        o268(.A(ori_ori_n290_), .B(ori_ori_n271_), .C(ori_ori_n268_), .Y(ori3));
  NO3        o269(.A(ori_ori_n142_), .B(ori_ori_n38_), .C(i_0_), .Y(ori_ori_n292_));
  NO2        o270(.A(ori_ori_n326_), .B(ori_ori_n53_), .Y(ori_ori_n293_));
  NOi21      o271(.An(i_5_), .B(i_9_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n294_), .B(ori_ori_n152_), .Y(ori_ori_n295_));
  BUFFER     o273(.A(ori_ori_n131_), .Y(ori_ori_n296_));
  NA2        o274(.A(ori_ori_n296_), .B(ori_ori_n162_), .Y(ori_ori_n297_));
  NO2        o275(.A(ori_ori_n297_), .B(ori_ori_n295_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n298_), .B(ori_ori_n293_), .Y(ori_ori_n299_));
  NA2        o277(.A(i_9_), .B(i_0_), .Y(ori_ori_n300_));
  NA2        o278(.A(i_0_), .B(i_10_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n203_), .B(ori_ori_n93_), .Y(ori_ori_n302_));
  NA2        o280(.A(ori_ori_n115_), .B(ori_ori_n85_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n269_), .B(ori_ori_n303_), .Y(ori_ori_n304_));
  INV        o282(.A(ori_ori_n304_), .Y(ori_ori_n305_));
  NA2        o283(.A(ori_ori_n129_), .B(ori_ori_n125_), .Y(ori_ori_n306_));
  AOI210     o284(.A0(ori_ori_n306_), .A1(ori_ori_n300_), .B0(ori_ori_n112_), .Y(ori_ori_n307_));
  INV        o285(.A(ori_ori_n307_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n308_), .B(ori_ori_n305_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n301_), .B(ori_ori_n294_), .Y(ori_ori_n310_));
  AOI220     o288(.A0(ori_ori_n310_), .A1(i_11_), .B0(ori_ori_n172_), .B1(ori_ori_n64_), .Y(ori_ori_n311_));
  NO3        o289(.A(ori_ori_n122_), .B(ori_ori_n142_), .C(i_0_), .Y(ori_ori_n312_));
  OAI210     o290(.A0(ori_ori_n312_), .A1(ori_ori_n65_), .B0(i_13_), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n313_), .B(ori_ori_n311_), .Y(ori_ori_n314_));
  NA3        o292(.A(ori_ori_n143_), .B(ori_ori_n115_), .C(ori_ori_n114_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n315_), .B(ori_ori_n164_), .Y(ori_ori_n316_));
  NO3        o294(.A(ori_ori_n316_), .B(ori_ori_n314_), .C(ori_ori_n309_), .Y(ori_ori_n317_));
  INV        o295(.A(ori_ori_n186_), .Y(ori_ori_n318_));
  NA2        o296(.A(ori_ori_n318_), .B(ori_ori_n120_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n319_), .B(ori_ori_n62_), .Y(ori_ori_n320_));
  INV        o298(.A(ori_ori_n320_), .Y(ori_ori_n321_));
  NA4        o299(.A(ori_ori_n321_), .B(ori_ori_n317_), .C(ori_ori_n302_), .D(ori_ori_n299_), .Y(ori4));
  INV        o300(.A(i_6_), .Y(ori_ori_n325_));
  INV        o301(.A(ori_ori_n292_), .Y(ori_ori_n326_));
  INV        o302(.A(i_6_), .Y(ori_ori_n327_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NOi21      m016(.An(i_12_), .B(i_13_), .Y(mai_mai_n39_));
  INV        m017(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NAi31      m018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n41_));
  INV        m019(.A(mai_mai_n35_), .Y(mai1));
  INV        m020(.A(i_11_), .Y(mai_mai_n43_));
  NO2        m021(.A(mai_mai_n43_), .B(i_6_), .Y(mai_mai_n44_));
  INV        m022(.A(i_2_), .Y(mai_mai_n45_));
  NA2        m023(.A(i_0_), .B(i_3_), .Y(mai_mai_n46_));
  INV        m024(.A(i_5_), .Y(mai_mai_n47_));
  NO2        m025(.A(i_7_), .B(i_10_), .Y(mai_mai_n48_));
  AOI210     m026(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n48_), .Y(mai_mai_n49_));
  NO2        m027(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n50_));
  NA2        m028(.A(i_0_), .B(i_2_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_7_), .B(i_9_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NA2        m031(.A(mai_mai_n50_), .B(mai_mai_n44_), .Y(mai_mai_n54_));
  NA3        m032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n55_));
  NO2        m033(.A(i_1_), .B(i_6_), .Y(mai_mai_n56_));
  NA2        m034(.A(i_8_), .B(i_7_), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  NA2        m036(.A(mai_mai_n58_), .B(i_12_), .Y(mai_mai_n59_));
  NAi21      m037(.An(i_2_), .B(i_7_), .Y(mai_mai_n60_));
  INV        m038(.A(i_1_), .Y(mai_mai_n61_));
  NA3        m039(.A(i_1_), .B(mai_mai_n60_), .C(mai_mai_n31_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n62_), .B(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n49_), .B(i_2_), .Y(mai_mai_n64_));
  NA2        m042(.A(i_1_), .B(i_6_), .Y(mai_mai_n65_));
  NO2        m043(.A(mai_mai_n65_), .B(mai_mai_n25_), .Y(mai_mai_n66_));
  INV        m044(.A(i_0_), .Y(mai_mai_n67_));
  NAi21      m045(.An(i_5_), .B(i_10_), .Y(mai_mai_n68_));
  NA2        m046(.A(i_5_), .B(i_9_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n68_), .B0(mai_mai_n67_), .Y(mai_mai_n70_));
  NO2        m048(.A(mai_mai_n70_), .B(mai_mai_n66_), .Y(mai_mai_n71_));
  NA2        m049(.A(mai_mai_n64_), .B(mai_mai_n71_), .Y(mai_mai_n72_));
  OAI210     m050(.A0(mai_mai_n72_), .A1(mai_mai_n63_), .B0(i_0_), .Y(mai_mai_n73_));
  NA2        m051(.A(i_12_), .B(i_5_), .Y(mai_mai_n74_));
  NO2        m052(.A(i_3_), .B(i_9_), .Y(mai_mai_n75_));
  NO2        m053(.A(i_3_), .B(i_7_), .Y(mai_mai_n76_));
  INV        m054(.A(i_6_), .Y(mai_mai_n77_));
  OR4        m055(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n78_));
  INV        m056(.A(mai_mai_n78_), .Y(mai_mai_n79_));
  NO2        m057(.A(i_2_), .B(i_7_), .Y(mai_mai_n80_));
  NAi21      m058(.An(i_6_), .B(i_10_), .Y(mai_mai_n81_));
  NA2        m059(.A(i_6_), .B(i_9_), .Y(mai_mai_n82_));
  AOI210     m060(.A0(mai_mai_n82_), .A1(mai_mai_n81_), .B0(mai_mai_n61_), .Y(mai_mai_n83_));
  NA2        m061(.A(i_2_), .B(i_6_), .Y(mai_mai_n84_));
  INV        m062(.A(mai_mai_n83_), .Y(mai_mai_n85_));
  NO2        m063(.A(mai_mai_n85_), .B(mai_mai_n74_), .Y(mai_mai_n86_));
  AN3        m064(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n87_));
  NAi21      m065(.An(i_6_), .B(i_11_), .Y(mai_mai_n88_));
  NO2        m066(.A(i_5_), .B(i_8_), .Y(mai_mai_n89_));
  NOi21      m067(.An(mai_mai_n89_), .B(mai_mai_n88_), .Y(mai_mai_n90_));
  AOI220     m068(.A0(mai_mai_n90_), .A1(mai_mai_n60_), .B0(mai_mai_n87_), .B1(mai_mai_n32_), .Y(mai_mai_n91_));
  INV        m069(.A(i_7_), .Y(mai_mai_n92_));
  NA2        m070(.A(mai_mai_n45_), .B(mai_mai_n92_), .Y(mai_mai_n93_));
  NO2        m071(.A(i_0_), .B(i_5_), .Y(mai_mai_n94_));
  NO2        m072(.A(mai_mai_n94_), .B(mai_mai_n77_), .Y(mai_mai_n95_));
  NA2        m073(.A(i_12_), .B(i_3_), .Y(mai_mai_n96_));
  INV        m074(.A(mai_mai_n96_), .Y(mai_mai_n97_));
  NA3        m075(.A(mai_mai_n97_), .B(mai_mai_n95_), .C(mai_mai_n93_), .Y(mai_mai_n98_));
  NAi21      m076(.An(i_7_), .B(i_11_), .Y(mai_mai_n99_));
  AN2        m077(.A(i_2_), .B(i_10_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(i_7_), .Y(mai_mai_n101_));
  OR2        m079(.A(mai_mai_n74_), .B(mai_mai_n56_), .Y(mai_mai_n102_));
  NO2        m080(.A(i_8_), .B(mai_mai_n92_), .Y(mai_mai_n103_));
  NO3        m081(.A(mai_mai_n103_), .B(mai_mai_n102_), .C(mai_mai_n101_), .Y(mai_mai_n104_));
  NA2        m082(.A(i_12_), .B(i_7_), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n61_), .B(mai_mai_n26_), .Y(mai_mai_n106_));
  NA2        m084(.A(mai_mai_n106_), .B(i_0_), .Y(mai_mai_n107_));
  NA2        m085(.A(i_11_), .B(i_12_), .Y(mai_mai_n108_));
  OAI210     m086(.A0(mai_mai_n107_), .A1(mai_mai_n105_), .B0(mai_mai_n108_), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n109_), .B(mai_mai_n104_), .Y(mai_mai_n110_));
  NA3        m088(.A(mai_mai_n110_), .B(mai_mai_n98_), .C(mai_mai_n91_), .Y(mai_mai_n111_));
  NOi21      m089(.An(i_1_), .B(i_5_), .Y(mai_mai_n112_));
  NA2        m090(.A(mai_mai_n112_), .B(i_11_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n92_), .B(mai_mai_n37_), .Y(mai_mai_n114_));
  NA2        m092(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n115_));
  NA2        m093(.A(mai_mai_n115_), .B(mai_mai_n114_), .Y(mai_mai_n116_));
  NO2        m094(.A(mai_mai_n116_), .B(mai_mai_n45_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n82_), .B(mai_mai_n81_), .Y(mai_mai_n118_));
  NAi21      m096(.An(i_3_), .B(i_8_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(mai_mai_n60_), .Y(mai_mai_n120_));
  NO2        m098(.A(i_1_), .B(mai_mai_n77_), .Y(mai_mai_n121_));
  NO2        m099(.A(i_6_), .B(i_5_), .Y(mai_mai_n122_));
  NA2        m100(.A(mai_mai_n122_), .B(i_3_), .Y(mai_mai_n123_));
  AO210      m101(.A0(mai_mai_n123_), .A1(mai_mai_n46_), .B0(mai_mai_n121_), .Y(mai_mai_n124_));
  OAI220     m102(.A0(mai_mai_n124_), .A1(mai_mai_n99_), .B0(mai_mai_n120_), .B1(mai_mai_n113_), .Y(mai_mai_n125_));
  NO3        m103(.A(mai_mai_n125_), .B(mai_mai_n111_), .C(mai_mai_n86_), .Y(mai_mai_n126_));
  NA3        m104(.A(mai_mai_n126_), .B(mai_mai_n73_), .C(mai_mai_n54_), .Y(mai2));
  NO2        m105(.A(mai_mai_n61_), .B(mai_mai_n37_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n868_), .B(mai_mai_n128_), .Y(mai_mai_n129_));
  NA4        m107(.A(mai_mai_n129_), .B(mai_mai_n71_), .C(mai_mai_n64_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m108(.A(i_8_), .B(i_7_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n131_), .B(i_6_), .Y(mai_mai_n132_));
  NO2        m110(.A(i_12_), .B(i_13_), .Y(mai_mai_n133_));
  NAi21      m111(.An(i_5_), .B(i_11_), .Y(mai_mai_n134_));
  NOi21      m112(.An(mai_mai_n133_), .B(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m113(.A(i_0_), .B(i_1_), .Y(mai_mai_n136_));
  AN2        m114(.A(mai_mai_n133_), .B(mai_mai_n75_), .Y(mai_mai_n137_));
  NA2        m115(.A(i_1_), .B(i_5_), .Y(mai_mai_n138_));
  NO2        m116(.A(mai_mai_n67_), .B(mai_mai_n45_), .Y(mai_mai_n139_));
  NA2        m117(.A(mai_mai_n139_), .B(mai_mai_n36_), .Y(mai_mai_n140_));
  NO3        m118(.A(mai_mai_n140_), .B(mai_mai_n138_), .C(i_13_), .Y(mai_mai_n141_));
  OR2        m119(.A(i_0_), .B(i_1_), .Y(mai_mai_n142_));
  NO3        m120(.A(mai_mai_n142_), .B(mai_mai_n74_), .C(i_13_), .Y(mai_mai_n143_));
  NAi32      m121(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n144_));
  NAi21      m122(.An(mai_mai_n144_), .B(mai_mai_n143_), .Y(mai_mai_n145_));
  NOi21      m123(.An(i_4_), .B(i_10_), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n146_), .B(mai_mai_n39_), .Y(mai_mai_n147_));
  NO2        m125(.A(i_3_), .B(i_5_), .Y(mai_mai_n148_));
  NA2        m126(.A(i_0_), .B(mai_mai_n148_), .Y(mai_mai_n149_));
  OAI210     m127(.A0(mai_mai_n149_), .A1(mai_mai_n147_), .B0(mai_mai_n145_), .Y(mai_mai_n150_));
  NO2        m128(.A(mai_mai_n150_), .B(mai_mai_n141_), .Y(mai_mai_n151_));
  NO2        m129(.A(mai_mai_n151_), .B(mai_mai_n132_), .Y(mai_mai_n152_));
  NOi21      m130(.An(i_4_), .B(i_9_), .Y(mai_mai_n153_));
  NOi21      m131(.An(i_11_), .B(i_13_), .Y(mai_mai_n154_));
  NA2        m132(.A(mai_mai_n154_), .B(mai_mai_n153_), .Y(mai_mai_n155_));
  NO2        m133(.A(i_4_), .B(i_5_), .Y(mai_mai_n156_));
  NAi21      m134(.An(i_12_), .B(i_11_), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n157_), .B(i_13_), .Y(mai_mai_n158_));
  NO2        m136(.A(mai_mai_n67_), .B(mai_mai_n61_), .Y(mai_mai_n159_));
  NAi31      m137(.An(i_4_), .B(mai_mai_n137_), .C(i_11_), .Y(mai_mai_n160_));
  NA2        m138(.A(i_3_), .B(i_5_), .Y(mai_mai_n161_));
  BUFFER     m139(.A(mai_mai_n155_), .Y(mai_mai_n162_));
  AOI210     m140(.A0(mai_mai_n162_), .A1(mai_mai_n160_), .B0(mai_mai_n61_), .Y(mai_mai_n163_));
  NO2        m141(.A(mai_mai_n67_), .B(i_5_), .Y(mai_mai_n164_));
  NO2        m142(.A(i_13_), .B(i_10_), .Y(mai_mai_n165_));
  NA3        m143(.A(mai_mai_n165_), .B(mai_mai_n164_), .C(mai_mai_n43_), .Y(mai_mai_n166_));
  NO2        m144(.A(i_2_), .B(i_1_), .Y(mai_mai_n167_));
  NA2        m145(.A(mai_mai_n167_), .B(i_3_), .Y(mai_mai_n168_));
  NAi21      m146(.An(i_4_), .B(i_12_), .Y(mai_mai_n169_));
  NO4        m147(.A(mai_mai_n169_), .B(mai_mai_n168_), .C(mai_mai_n166_), .D(mai_mai_n25_), .Y(mai_mai_n170_));
  NO2        m148(.A(mai_mai_n170_), .B(mai_mai_n163_), .Y(mai_mai_n171_));
  INV        m149(.A(i_8_), .Y(mai_mai_n172_));
  NA2        m150(.A(i_8_), .B(i_6_), .Y(mai_mai_n173_));
  NO3        m151(.A(i_3_), .B(mai_mai_n77_), .C(mai_mai_n47_), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n174_), .B(mai_mai_n103_), .Y(mai_mai_n175_));
  NO3        m153(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n176_));
  NA3        m154(.A(mai_mai_n176_), .B(mai_mai_n39_), .C(mai_mai_n43_), .Y(mai_mai_n177_));
  NO3        m155(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n178_));
  NA2        m156(.A(i_12_), .B(mai_mai_n178_), .Y(mai_mai_n179_));
  AOI210     m157(.A0(mai_mai_n179_), .A1(mai_mai_n177_), .B0(mai_mai_n175_), .Y(mai_mai_n180_));
  NO2        m158(.A(i_3_), .B(i_8_), .Y(mai_mai_n181_));
  NO3        m159(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n94_), .B(mai_mai_n56_), .Y(mai_mai_n183_));
  NO2        m161(.A(i_13_), .B(i_9_), .Y(mai_mai_n184_));
  NA2        m162(.A(mai_mai_n184_), .B(mai_mai_n172_), .Y(mai_mai_n185_));
  NAi21      m163(.An(i_12_), .B(i_3_), .Y(mai_mai_n186_));
  NO2        m164(.A(mai_mai_n43_), .B(i_5_), .Y(mai_mai_n187_));
  NO3        m165(.A(i_0_), .B(i_2_), .C(mai_mai_n61_), .Y(mai_mai_n188_));
  INV        m166(.A(mai_mai_n180_), .Y(mai_mai_n189_));
  OAI220     m167(.A0(mai_mai_n189_), .A1(i_4_), .B0(mai_mai_n173_), .B1(mai_mai_n171_), .Y(mai_mai_n190_));
  NAi21      m168(.An(i_12_), .B(i_7_), .Y(mai_mai_n191_));
  NA3        m169(.A(i_13_), .B(mai_mai_n172_), .C(i_10_), .Y(mai_mai_n192_));
  NO2        m170(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n193_));
  NA2        m171(.A(i_0_), .B(i_5_), .Y(mai_mai_n194_));
  OAI220     m172(.A0(mai_mai_n77_), .A1(mai_mai_n168_), .B0(mai_mai_n61_), .B1(mai_mai_n123_), .Y(mai_mai_n195_));
  NAi31      m173(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n197_));
  NO2        m175(.A(mai_mai_n45_), .B(mai_mai_n61_), .Y(mai_mai_n198_));
  NA2        m176(.A(mai_mai_n198_), .B(mai_mai_n197_), .Y(mai_mai_n199_));
  INV        m177(.A(i_13_), .Y(mai_mai_n200_));
  NO2        m178(.A(i_12_), .B(mai_mai_n200_), .Y(mai_mai_n201_));
  NA3        m179(.A(mai_mai_n201_), .B(mai_mai_n176_), .C(mai_mai_n174_), .Y(mai_mai_n202_));
  INV        m180(.A(mai_mai_n202_), .Y(mai_mai_n203_));
  AOI220     m181(.A0(mai_mai_n203_), .A1(mai_mai_n131_), .B0(mai_mai_n195_), .B1(mai_mai_n193_), .Y(mai_mai_n204_));
  NO2        m182(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n161_), .B(i_4_), .Y(mai_mai_n206_));
  NA2        m184(.A(mai_mai_n206_), .B(mai_mai_n205_), .Y(mai_mai_n207_));
  OR2        m185(.A(i_8_), .B(i_7_), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n208_), .B(mai_mai_n77_), .Y(mai_mai_n209_));
  INV        m187(.A(i_12_), .Y(mai_mai_n210_));
  NO3        m188(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n211_));
  NA2        m189(.A(i_2_), .B(i_1_), .Y(mai_mai_n212_));
  NAi21      m190(.An(i_4_), .B(i_3_), .Y(mai_mai_n213_));
  NO2        m191(.A(i_0_), .B(i_6_), .Y(mai_mai_n214_));
  NOi41      m192(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n215_));
  NO2        m193(.A(i_11_), .B(mai_mai_n200_), .Y(mai_mai_n216_));
  NAi21      m194(.An(i_3_), .B(i_7_), .Y(mai_mai_n217_));
  NA2        m195(.A(mai_mai_n210_), .B(i_9_), .Y(mai_mai_n218_));
  OR2        m196(.A(mai_mai_n218_), .B(mai_mai_n217_), .Y(mai_mai_n219_));
  NO2        m197(.A(i_12_), .B(i_3_), .Y(mai_mai_n220_));
  NA2        m198(.A(i_3_), .B(i_9_), .Y(mai_mai_n221_));
  NAi21      m199(.An(i_7_), .B(i_10_), .Y(mai_mai_n222_));
  NO2        m200(.A(mai_mai_n222_), .B(mai_mai_n221_), .Y(mai_mai_n223_));
  INV        m201(.A(mai_mai_n219_), .Y(mai_mai_n224_));
  INV        m202(.A(mai_mai_n132_), .Y(mai_mai_n225_));
  NA2        m203(.A(mai_mai_n210_), .B(i_13_), .Y(mai_mai_n226_));
  NO2        m204(.A(mai_mai_n226_), .B(mai_mai_n69_), .Y(mai_mai_n227_));
  AOI220     m205(.A0(mai_mai_n227_), .A1(mai_mai_n225_), .B0(mai_mai_n224_), .B1(mai_mai_n216_), .Y(mai_mai_n228_));
  NO2        m206(.A(mai_mai_n208_), .B(mai_mai_n37_), .Y(mai_mai_n229_));
  NA2        m207(.A(i_12_), .B(i_6_), .Y(mai_mai_n230_));
  OR2        m208(.A(i_13_), .B(i_9_), .Y(mai_mai_n231_));
  NO3        m209(.A(mai_mai_n231_), .B(mai_mai_n230_), .C(mai_mai_n47_), .Y(mai_mai_n232_));
  NO2        m210(.A(mai_mai_n213_), .B(i_2_), .Y(mai_mai_n233_));
  NA3        m211(.A(mai_mai_n233_), .B(mai_mai_n232_), .C(mai_mai_n43_), .Y(mai_mai_n234_));
  NA2        m212(.A(mai_mai_n216_), .B(i_9_), .Y(mai_mai_n235_));
  OAI210     m213(.A0(mai_mai_n61_), .A1(mai_mai_n235_), .B0(mai_mai_n234_), .Y(mai_mai_n236_));
  NA2        m214(.A(mai_mai_n139_), .B(mai_mai_n61_), .Y(mai_mai_n237_));
  NO3        m215(.A(i_11_), .B(mai_mai_n200_), .C(mai_mai_n25_), .Y(mai_mai_n238_));
  NO2        m216(.A(mai_mai_n217_), .B(i_8_), .Y(mai_mai_n239_));
  NO2        m217(.A(i_6_), .B(mai_mai_n47_), .Y(mai_mai_n240_));
  NA2        m218(.A(mai_mai_n239_), .B(mai_mai_n238_), .Y(mai_mai_n241_));
  NA3        m219(.A(i_3_), .B(mai_mai_n229_), .C(mai_mai_n201_), .Y(mai_mai_n242_));
  AOI210     m220(.A0(mai_mai_n242_), .A1(mai_mai_n241_), .B0(mai_mai_n237_), .Y(mai_mai_n243_));
  AOI210     m221(.A0(mai_mai_n236_), .A1(mai_mai_n229_), .B0(mai_mai_n243_), .Y(mai_mai_n244_));
  NA3        m222(.A(mai_mai_n244_), .B(mai_mai_n228_), .C(mai_mai_n204_), .Y(mai_mai_n245_));
  NO3        m223(.A(i_12_), .B(mai_mai_n200_), .C(mai_mai_n37_), .Y(mai_mai_n246_));
  INV        m224(.A(mai_mai_n246_), .Y(mai_mai_n247_));
  NA2        m225(.A(i_8_), .B(mai_mai_n92_), .Y(mai_mai_n248_));
  NO2        m226(.A(i_3_), .B(mai_mai_n248_), .Y(mai_mai_n249_));
  NO2        m227(.A(mai_mai_n212_), .B(i_0_), .Y(mai_mai_n250_));
  AOI220     m228(.A0(mai_mai_n250_), .A1(i_8_), .B0(i_1_), .B1(mai_mai_n131_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n240_), .B(mai_mai_n26_), .Y(mai_mai_n252_));
  NO2        m230(.A(mai_mai_n252_), .B(mai_mai_n251_), .Y(mai_mai_n253_));
  NA2        m231(.A(i_0_), .B(i_1_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n254_), .B(i_2_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n57_), .B(i_6_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n256_), .B(mai_mai_n255_), .Y(mai_mai_n257_));
  OAI210     m235(.A0(mai_mai_n149_), .A1(mai_mai_n132_), .B0(mai_mai_n257_), .Y(mai_mai_n258_));
  NO3        m236(.A(mai_mai_n258_), .B(mai_mai_n253_), .C(mai_mai_n249_), .Y(mai_mai_n259_));
  NO2        m237(.A(i_3_), .B(i_10_), .Y(mai_mai_n260_));
  NA3        m238(.A(mai_mai_n260_), .B(mai_mai_n39_), .C(mai_mai_n43_), .Y(mai_mai_n261_));
  AN2        m239(.A(i_3_), .B(i_10_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n45_), .B(mai_mai_n26_), .Y(mai_mai_n263_));
  NO2        m241(.A(mai_mai_n259_), .B(mai_mai_n247_), .Y(mai_mai_n264_));
  NO4        m242(.A(mai_mai_n264_), .B(mai_mai_n245_), .C(mai_mai_n190_), .D(mai_mai_n152_), .Y(mai_mai_n265_));
  NO3        m243(.A(mai_mai_n43_), .B(i_13_), .C(i_9_), .Y(mai_mai_n266_));
  NO3        m244(.A(i_6_), .B(mai_mai_n172_), .C(i_7_), .Y(mai_mai_n267_));
  NO2        m245(.A(i_2_), .B(i_3_), .Y(mai_mai_n268_));
  INV        m246(.A(mai_mai_n194_), .Y(mai_mai_n269_));
  NA3        m247(.A(mai_mai_n209_), .B(mai_mai_n268_), .C(i_1_), .Y(mai_mai_n270_));
  NA2        m248(.A(mai_mai_n45_), .B(mai_mai_n270_), .Y(mai_mai_n271_));
  NA2        m249(.A(mai_mai_n271_), .B(i_4_), .Y(mai_mai_n272_));
  NO2        m250(.A(i_12_), .B(i_10_), .Y(mai_mai_n273_));
  NOi21      m251(.An(i_5_), .B(i_0_), .Y(mai_mai_n274_));
  NA4        m252(.A(mai_mai_n76_), .B(mai_mai_n36_), .C(mai_mai_n77_), .D(i_8_), .Y(mai_mai_n275_));
  NO2        m253(.A(i_6_), .B(i_8_), .Y(mai_mai_n276_));
  AN2        m254(.A(i_0_), .B(mai_mai_n276_), .Y(mai_mai_n277_));
  NO2        m255(.A(i_1_), .B(i_7_), .Y(mai_mai_n278_));
  NA2        m256(.A(mai_mai_n277_), .B(i_4_), .Y(mai_mai_n279_));
  NA2        m257(.A(mai_mai_n279_), .B(mai_mai_n272_), .Y(mai_mai_n280_));
  NO2        m258(.A(i_8_), .B(mai_mai_n269_), .Y(mai_mai_n281_));
  OAI210     m259(.A0(mai_mai_n25_), .A1(mai_mai_n281_), .B0(i_3_), .Y(mai_mai_n282_));
  NO2        m260(.A(mai_mai_n84_), .B(mai_mai_n172_), .Y(mai_mai_n283_));
  NO2        m261(.A(mai_mai_n172_), .B(i_9_), .Y(mai_mai_n284_));
  NO3        m262(.A(mai_mai_n284_), .B(mai_mai_n283_), .C(mai_mai_n253_), .Y(mai_mai_n285_));
  AOI210     m263(.A0(mai_mai_n285_), .A1(mai_mai_n282_), .B0(mai_mai_n147_), .Y(mai_mai_n286_));
  AOI210     m264(.A0(mai_mai_n280_), .A1(mai_mai_n266_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  NOi32      m265(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n288_));
  INV        m266(.A(mai_mai_n288_), .Y(mai_mai_n289_));
  NAi21      m267(.An(i_1_), .B(i_5_), .Y(mai_mai_n290_));
  NA2        m268(.A(mai_mai_n290_), .B(i_0_), .Y(mai_mai_n291_));
  NA2        m269(.A(mai_mai_n291_), .B(mai_mai_n25_), .Y(mai_mai_n292_));
  NO2        m270(.A(mai_mai_n292_), .B(mai_mai_n144_), .Y(mai_mai_n293_));
  NO2        m271(.A(mai_mai_n196_), .B(mai_mai_n144_), .Y(mai_mai_n294_));
  NO2        m272(.A(mai_mai_n144_), .B(mai_mai_n142_), .Y(mai_mai_n295_));
  NOi32      m273(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n296_));
  NA2        m274(.A(mai_mai_n296_), .B(mai_mai_n45_), .Y(mai_mai_n297_));
  NO2        m275(.A(mai_mai_n297_), .B(i_0_), .Y(mai_mai_n298_));
  OR3        m276(.A(mai_mai_n298_), .B(mai_mai_n295_), .C(mai_mai_n294_), .Y(mai_mai_n299_));
  NO2        m277(.A(i_1_), .B(mai_mai_n92_), .Y(mai_mai_n300_));
  NAi21      m278(.An(i_3_), .B(i_4_), .Y(mai_mai_n301_));
  NO2        m279(.A(mai_mai_n301_), .B(i_9_), .Y(mai_mai_n302_));
  NA2        m280(.A(i_7_), .B(mai_mai_n302_), .Y(mai_mai_n303_));
  NA2        m281(.A(i_2_), .B(i_7_), .Y(mai_mai_n304_));
  NO2        m282(.A(mai_mai_n301_), .B(i_10_), .Y(mai_mai_n305_));
  NA3        m283(.A(mai_mai_n305_), .B(mai_mai_n304_), .C(mai_mai_n214_), .Y(mai_mai_n306_));
  AOI210     m284(.A0(mai_mai_n306_), .A1(mai_mai_n303_), .B0(mai_mai_n164_), .Y(mai_mai_n307_));
  AOI210     m285(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n308_));
  OAI210     m286(.A0(mai_mai_n308_), .A1(mai_mai_n167_), .B0(mai_mai_n305_), .Y(mai_mai_n309_));
  AOI220     m287(.A0(mai_mai_n305_), .A1(mai_mai_n278_), .B0(mai_mai_n211_), .B1(mai_mai_n167_), .Y(mai_mai_n310_));
  AOI210     m288(.A0(mai_mai_n310_), .A1(mai_mai_n309_), .B0(i_5_), .Y(mai_mai_n311_));
  NO4        m289(.A(mai_mai_n311_), .B(mai_mai_n307_), .C(mai_mai_n299_), .D(mai_mai_n293_), .Y(mai_mai_n312_));
  NO2        m290(.A(mai_mai_n312_), .B(mai_mai_n289_), .Y(mai_mai_n313_));
  NO2        m291(.A(mai_mai_n57_), .B(mai_mai_n25_), .Y(mai_mai_n314_));
  AN2        m292(.A(i_12_), .B(i_5_), .Y(mai_mai_n315_));
  NO2        m293(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n316_), .B(mai_mai_n315_), .Y(mai_mai_n317_));
  NO2        m295(.A(i_11_), .B(i_6_), .Y(mai_mai_n318_));
  NA3        m296(.A(mai_mai_n318_), .B(i_2_), .C(mai_mai_n200_), .Y(mai_mai_n319_));
  NO2        m297(.A(mai_mai_n319_), .B(mai_mai_n317_), .Y(mai_mai_n320_));
  NO2        m298(.A(mai_mai_n213_), .B(i_5_), .Y(mai_mai_n321_));
  NO2        m299(.A(i_5_), .B(i_10_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n133_), .B(mai_mai_n44_), .Y(mai_mai_n323_));
  NO2        m301(.A(mai_mai_n323_), .B(mai_mai_n213_), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n324_), .B(mai_mai_n314_), .Y(mai_mai_n325_));
  NO2        m303(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n326_));
  INV        m304(.A(mai_mai_n320_), .Y(mai_mai_n327_));
  NO2        m305(.A(i_11_), .B(i_12_), .Y(mai_mai_n328_));
  NA2        m306(.A(mai_mai_n322_), .B(mai_mai_n210_), .Y(mai_mai_n329_));
  NO2        m307(.A(mai_mai_n92_), .B(mai_mai_n196_), .Y(mai_mai_n330_));
  NO2        m308(.A(i_13_), .B(mai_mai_n212_), .Y(mai_mai_n331_));
  NA2        m309(.A(mai_mai_n330_), .B(mai_mai_n331_), .Y(mai_mai_n332_));
  NA3        m310(.A(mai_mai_n332_), .B(mai_mai_n327_), .C(mai_mai_n325_), .Y(mai_mai_n333_));
  NO2        m311(.A(i_0_), .B(i_11_), .Y(mai_mai_n334_));
  NOi21      m312(.An(i_2_), .B(i_12_), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n131_), .B(i_9_), .Y(mai_mai_n336_));
  NO2        m314(.A(mai_mai_n336_), .B(i_4_), .Y(mai_mai_n337_));
  NA2        m315(.A(mai_mai_n335_), .B(mai_mai_n337_), .Y(mai_mai_n338_));
  NAi21      m316(.An(i_9_), .B(i_4_), .Y(mai_mai_n339_));
  OR2        m317(.A(i_13_), .B(i_10_), .Y(mai_mai_n340_));
  NO2        m318(.A(mai_mai_n155_), .B(mai_mai_n114_), .Y(mai_mai_n341_));
  BUFFER     m319(.A(mai_mai_n192_), .Y(mai_mai_n342_));
  NO2        m320(.A(mai_mai_n92_), .B(mai_mai_n25_), .Y(mai_mai_n343_));
  NA2        m321(.A(mai_mai_n246_), .B(mai_mai_n343_), .Y(mai_mai_n344_));
  NA2        m322(.A(mai_mai_n240_), .B(mai_mai_n188_), .Y(mai_mai_n345_));
  OAI220     m323(.A0(mai_mai_n345_), .A1(mai_mai_n342_), .B0(mai_mai_n344_), .B1(mai_mai_n94_), .Y(mai_mai_n346_));
  INV        m324(.A(mai_mai_n346_), .Y(mai_mai_n347_));
  AOI210     m325(.A0(mai_mai_n347_), .A1(mai_mai_n338_), .B0(mai_mai_n26_), .Y(mai_mai_n348_));
  INV        m326(.A(mai_mai_n270_), .Y(mai_mai_n349_));
  AOI220     m327(.A0(mai_mai_n256_), .A1(i_2_), .B0(mai_mai_n250_), .B1(i_7_), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n350_), .B(i_5_), .Y(mai_mai_n351_));
  AOI220     m329(.A0(i_3_), .A1(mai_mai_n255_), .B0(i_3_), .B1(mai_mai_n188_), .Y(mai_mai_n352_));
  NO2        m330(.A(mai_mai_n352_), .B(mai_mai_n248_), .Y(mai_mai_n353_));
  NO3        m331(.A(mai_mai_n353_), .B(mai_mai_n351_), .C(mai_mai_n349_), .Y(mai_mai_n354_));
  NA2        m332(.A(mai_mai_n174_), .B(mai_mai_n87_), .Y(mai_mai_n355_));
  NA3        m333(.A(i_2_), .B(mai_mai_n148_), .C(mai_mai_n77_), .Y(mai_mai_n356_));
  AOI210     m334(.A0(mai_mai_n356_), .A1(mai_mai_n355_), .B0(i_8_), .Y(mai_mai_n357_));
  NA2        m335(.A(mai_mai_n172_), .B(i_10_), .Y(mai_mai_n358_));
  NA2        m336(.A(i_1_), .B(i_2_), .Y(mai_mai_n359_));
  NA2        m337(.A(mai_mai_n256_), .B(i_2_), .Y(mai_mai_n360_));
  OAI220     m338(.A0(mai_mai_n360_), .A1(mai_mai_n161_), .B0(mai_mai_n359_), .B1(mai_mai_n358_), .Y(mai_mai_n361_));
  NA3        m339(.A(mai_mai_n278_), .B(mai_mai_n277_), .C(i_5_), .Y(mai_mai_n362_));
  INV        m340(.A(mai_mai_n267_), .Y(mai_mai_n363_));
  OAI210     m341(.A0(mai_mai_n363_), .A1(mai_mai_n168_), .B0(mai_mai_n362_), .Y(mai_mai_n364_));
  NO3        m342(.A(mai_mai_n364_), .B(mai_mai_n361_), .C(mai_mai_n357_), .Y(mai_mai_n365_));
  AOI210     m343(.A0(mai_mai_n365_), .A1(mai_mai_n354_), .B0(mai_mai_n235_), .Y(mai_mai_n366_));
  NO4        m344(.A(mai_mai_n366_), .B(mai_mai_n348_), .C(mai_mai_n333_), .D(mai_mai_n313_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n67_), .B(i_13_), .Y(mai_mai_n368_));
  NA3        m346(.A(mai_mai_n368_), .B(i_1_), .C(i_2_), .Y(mai_mai_n369_));
  NO2        m347(.A(i_10_), .B(i_9_), .Y(mai_mai_n370_));
  NAi21      m348(.An(i_12_), .B(i_8_), .Y(mai_mai_n371_));
  NO2        m349(.A(mai_mai_n371_), .B(i_3_), .Y(mai_mai_n372_));
  NA2        m350(.A(mai_mai_n372_), .B(mai_mai_n370_), .Y(mai_mai_n373_));
  NO2        m351(.A(mai_mai_n373_), .B(mai_mai_n369_), .Y(mai_mai_n374_));
  INV        m352(.A(mai_mai_n263_), .Y(mai_mai_n375_));
  NO3        m353(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n376_));
  NA2        m354(.A(mai_mai_n230_), .B(mai_mai_n88_), .Y(mai_mai_n377_));
  NA2        m355(.A(i_8_), .B(i_9_), .Y(mai_mai_n378_));
  NA2        m356(.A(mai_mai_n246_), .B(mai_mai_n183_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n379_), .B(mai_mai_n378_), .Y(mai_mai_n380_));
  NO3        m358(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n381_));
  NA3        m359(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n382_));
  NA4        m360(.A(mai_mai_n134_), .B(mai_mai_n106_), .C(mai_mai_n74_), .D(mai_mai_n23_), .Y(mai_mai_n383_));
  NO2        m361(.A(mai_mai_n383_), .B(mai_mai_n382_), .Y(mai_mai_n384_));
  NO3        m362(.A(mai_mai_n384_), .B(mai_mai_n380_), .C(mai_mai_n374_), .Y(mai_mai_n385_));
  BUFFER     m363(.A(mai_mai_n257_), .Y(mai_mai_n386_));
  OA220      m364(.A0(mai_mai_n386_), .A1(mai_mai_n147_), .B0(mai_mai_n185_), .B1(mai_mai_n207_), .Y(mai_mai_n387_));
  NA2        m365(.A(mai_mai_n87_), .B(i_13_), .Y(mai_mai_n388_));
  NA2        m366(.A(i_3_), .B(mai_mai_n314_), .Y(mai_mai_n389_));
  NO2        m367(.A(i_2_), .B(i_13_), .Y(mai_mai_n390_));
  NA3        m368(.A(mai_mai_n390_), .B(mai_mai_n146_), .C(mai_mai_n90_), .Y(mai_mai_n391_));
  NO2        m369(.A(mai_mai_n389_), .B(mai_mai_n388_), .Y(mai_mai_n392_));
  NO3        m370(.A(i_4_), .B(mai_mai_n47_), .C(i_8_), .Y(mai_mai_n393_));
  NO2        m371(.A(i_6_), .B(i_7_), .Y(mai_mai_n394_));
  NOi21      m372(.An(i_2_), .B(i_7_), .Y(mai_mai_n395_));
  NAi31      m373(.An(i_11_), .B(mai_mai_n395_), .C(i_0_), .Y(mai_mai_n396_));
  NO2        m374(.A(mai_mai_n340_), .B(i_6_), .Y(mai_mai_n397_));
  NA2        m375(.A(mai_mai_n397_), .B(i_1_), .Y(mai_mai_n398_));
  NO2        m376(.A(mai_mai_n398_), .B(mai_mai_n396_), .Y(mai_mai_n399_));
  NO2        m377(.A(i_3_), .B(mai_mai_n172_), .Y(mai_mai_n400_));
  NO2        m378(.A(i_6_), .B(i_10_), .Y(mai_mai_n401_));
  NA3        m379(.A(mai_mai_n215_), .B(mai_mai_n154_), .C(mai_mai_n122_), .Y(mai_mai_n402_));
  NA2        m380(.A(mai_mai_n45_), .B(mai_mai_n43_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n142_), .B(i_3_), .Y(mai_mai_n404_));
  NAi31      m382(.An(mai_mai_n403_), .B(mai_mai_n404_), .C(mai_mai_n201_), .Y(mai_mai_n405_));
  NA2        m383(.A(mai_mai_n405_), .B(mai_mai_n402_), .Y(mai_mai_n406_));
  NO3        m384(.A(mai_mai_n406_), .B(mai_mai_n399_), .C(mai_mai_n392_), .Y(mai_mai_n407_));
  NA2        m385(.A(mai_mai_n381_), .B(mai_mai_n322_), .Y(mai_mai_n408_));
  NO2        m386(.A(mai_mai_n408_), .B(mai_mai_n199_), .Y(mai_mai_n409_));
  NAi21      m387(.An(mai_mai_n192_), .B(mai_mai_n328_), .Y(mai_mai_n410_));
  NO2        m388(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n411_));
  NA3        m389(.A(i_6_), .B(mai_mai_n411_), .C(mai_mai_n131_), .Y(mai_mai_n412_));
  OAI220     m390(.A0(mai_mai_n38_), .A1(mai_mai_n412_), .B0(i_7_), .B1(mai_mai_n410_), .Y(mai_mai_n413_));
  NA2        m391(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n414_));
  NO2        m392(.A(mai_mai_n414_), .B(mai_mai_n388_), .Y(mai_mai_n415_));
  NO3        m393(.A(mai_mai_n415_), .B(mai_mai_n413_), .C(mai_mai_n409_), .Y(mai_mai_n416_));
  NA4        m394(.A(mai_mai_n416_), .B(mai_mai_n407_), .C(mai_mai_n387_), .D(mai_mai_n385_), .Y(mai_mai_n417_));
  NA3        m395(.A(mai_mai_n262_), .B(mai_mai_n158_), .C(mai_mai_n156_), .Y(mai_mai_n418_));
  NA2        m396(.A(mai_mai_n376_), .B(mai_mai_n263_), .Y(mai_mai_n419_));
  NA4        m397(.A(mai_mai_n368_), .B(i_1_), .C(mai_mai_n181_), .D(i_2_), .Y(mai_mai_n420_));
  INV        m398(.A(mai_mai_n420_), .Y(mai_mai_n421_));
  NA2        m399(.A(mai_mai_n315_), .B(mai_mai_n200_), .Y(mai_mai_n422_));
  NA2        m400(.A(mai_mai_n288_), .B(mai_mai_n67_), .Y(mai_mai_n423_));
  NA2        m401(.A(i_7_), .B(mai_mai_n296_), .Y(mai_mai_n424_));
  AO210      m402(.A0(mai_mai_n423_), .A1(mai_mai_n422_), .B0(mai_mai_n424_), .Y(mai_mai_n425_));
  NO2        m403(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n426_));
  INV        m404(.A(mai_mai_n425_), .Y(mai_mai_n427_));
  AOI210     m405(.A0(mai_mai_n421_), .A1(mai_mai_n182_), .B0(mai_mai_n427_), .Y(mai_mai_n428_));
  NO2        m406(.A(i_7_), .B(mai_mai_n177_), .Y(mai_mai_n429_));
  INV        m407(.A(mai_mai_n161_), .Y(mai_mai_n430_));
  AOI210     m408(.A0(mai_mai_n430_), .A1(mai_mai_n429_), .B0(mai_mai_n341_), .Y(mai_mai_n431_));
  NA4        m409(.A(mai_mai_n431_), .B(mai_mai_n428_), .C(mai_mai_n419_), .D(mai_mai_n418_), .Y(mai_mai_n432_));
  NA2        m410(.A(mai_mai_n321_), .B(mai_mai_n255_), .Y(mai_mai_n433_));
  NA2        m411(.A(mai_mai_n317_), .B(mai_mai_n433_), .Y(mai_mai_n434_));
  NO2        m412(.A(i_12_), .B(mai_mai_n172_), .Y(mai_mai_n435_));
  NOi31      m413(.An(mai_mai_n267_), .B(mai_mai_n340_), .C(mai_mai_n38_), .Y(mai_mai_n436_));
  OAI210     m414(.A0(mai_mai_n436_), .A1(mai_mai_n435_), .B0(mai_mai_n434_), .Y(mai_mai_n437_));
  NO2        m415(.A(i_8_), .B(i_7_), .Y(mai_mai_n438_));
  NA2        m416(.A(mai_mai_n43_), .B(i_10_), .Y(mai_mai_n439_));
  NO2        m417(.A(mai_mai_n439_), .B(i_6_), .Y(mai_mai_n440_));
  NA3        m418(.A(mai_mai_n440_), .B(mai_mai_n865_), .C(mai_mai_n438_), .Y(mai_mai_n441_));
  OAI220     m419(.A0(mai_mai_n161_), .A1(mai_mai_n226_), .B0(mai_mai_n388_), .B1(mai_mai_n123_), .Y(mai_mai_n442_));
  NA2        m420(.A(mai_mai_n442_), .B(mai_mai_n229_), .Y(mai_mai_n443_));
  NA3        m421(.A(mai_mai_n262_), .B(mai_mai_n156_), .C(mai_mai_n87_), .Y(mai_mai_n444_));
  NO2        m422(.A(mai_mai_n142_), .B(i_5_), .Y(mai_mai_n445_));
  NA2        m423(.A(mai_mai_n445_), .B(mai_mai_n268_), .Y(mai_mai_n446_));
  NA2        m424(.A(mai_mai_n446_), .B(mai_mai_n444_), .Y(mai_mai_n447_));
  NA2        m425(.A(mai_mai_n447_), .B(mai_mai_n381_), .Y(mai_mai_n448_));
  NA4        m426(.A(mai_mai_n448_), .B(mai_mai_n443_), .C(mai_mai_n441_), .D(mai_mai_n437_), .Y(mai_mai_n449_));
  NA2        m427(.A(mai_mai_n435_), .B(mai_mai_n238_), .Y(mai_mai_n450_));
  NO2        m428(.A(i_2_), .B(mai_mai_n450_), .Y(mai_mai_n451_));
  INV        m429(.A(mai_mai_n451_), .Y(mai_mai_n452_));
  NO3        m430(.A(mai_mai_n41_), .B(i_2_), .C(mai_mai_n47_), .Y(mai_mai_n453_));
  NO3        m431(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n454_));
  NO2        m432(.A(mai_mai_n208_), .B(mai_mai_n36_), .Y(mai_mai_n455_));
  AN2        m433(.A(mai_mai_n455_), .B(mai_mai_n454_), .Y(mai_mai_n456_));
  OA210      m434(.A0(mai_mai_n456_), .A1(mai_mai_n453_), .B0(mai_mai_n288_), .Y(mai_mai_n457_));
  NO2        m435(.A(mai_mai_n340_), .B(i_1_), .Y(mai_mai_n458_));
  AN3        m436(.A(mai_mai_n458_), .B(mai_mai_n337_), .C(i_2_), .Y(mai_mai_n459_));
  NO2        m437(.A(mai_mai_n459_), .B(mai_mai_n457_), .Y(mai_mai_n460_));
  NO2        m438(.A(mai_mai_n77_), .B(mai_mai_n25_), .Y(mai_mai_n461_));
  NA2        m439(.A(mai_mai_n238_), .B(i_10_), .Y(mai_mai_n462_));
  NO2        m440(.A(mai_mai_n462_), .B(mai_mai_n375_), .Y(mai_mai_n463_));
  NO2        m441(.A(mai_mai_n105_), .B(mai_mai_n23_), .Y(mai_mai_n464_));
  INV        m442(.A(mai_mai_n267_), .Y(mai_mai_n465_));
  AOI220     m443(.A0(mai_mai_n465_), .A1(mai_mai_n360_), .B0(mai_mai_n162_), .B1(mai_mai_n160_), .Y(mai_mai_n466_));
  NOi21      m444(.An(mai_mai_n135_), .B(mai_mai_n275_), .Y(mai_mai_n467_));
  NO3        m445(.A(mai_mai_n467_), .B(mai_mai_n466_), .C(mai_mai_n463_), .Y(mai_mai_n468_));
  NO2        m446(.A(mai_mai_n423_), .B(mai_mai_n310_), .Y(mai_mai_n469_));
  INV        m447(.A(mai_mai_n268_), .Y(mai_mai_n470_));
  NO2        m448(.A(i_12_), .B(mai_mai_n77_), .Y(mai_mai_n471_));
  NA2        m449(.A(mai_mai_n471_), .B(mai_mai_n238_), .Y(mai_mai_n472_));
  NA2        m450(.A(mai_mai_n318_), .B(mai_mai_n246_), .Y(mai_mai_n473_));
  AOI210     m451(.A0(mai_mai_n473_), .A1(mai_mai_n472_), .B0(mai_mai_n470_), .Y(mai_mai_n474_));
  NO3        m452(.A(i_4_), .B(i_8_), .C(mai_mai_n261_), .Y(mai_mai_n475_));
  OR2        m453(.A(i_2_), .B(i_5_), .Y(mai_mai_n476_));
  NO2        m454(.A(i_2_), .B(mai_mai_n410_), .Y(mai_mai_n477_));
  NO4        m455(.A(mai_mai_n477_), .B(mai_mai_n475_), .C(mai_mai_n474_), .D(mai_mai_n469_), .Y(mai_mai_n478_));
  NA4        m456(.A(mai_mai_n478_), .B(mai_mai_n468_), .C(mai_mai_n460_), .D(mai_mai_n452_), .Y(mai_mai_n479_));
  NO4        m457(.A(mai_mai_n479_), .B(mai_mai_n449_), .C(mai_mai_n432_), .D(mai_mai_n417_), .Y(mai_mai_n480_));
  NA4        m458(.A(mai_mai_n480_), .B(mai_mai_n367_), .C(mai_mai_n287_), .D(mai_mai_n265_), .Y(mai7));
  NO2        m459(.A(mai_mai_n99_), .B(mai_mai_n81_), .Y(mai_mai_n482_));
  NA2        m460(.A(mai_mai_n401_), .B(mai_mai_n76_), .Y(mai_mai_n483_));
  NA2        m461(.A(i_11_), .B(mai_mai_n172_), .Y(mai_mai_n484_));
  NA3        m462(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n485_));
  NO2        m463(.A(mai_mai_n210_), .B(i_4_), .Y(mai_mai_n486_));
  NA2        m464(.A(mai_mai_n486_), .B(i_8_), .Y(mai_mai_n487_));
  AOI210     m465(.A0(mai_mai_n487_), .A1(mai_mai_n96_), .B0(mai_mai_n485_), .Y(mai_mai_n488_));
  OAI210     m466(.A0(mai_mai_n80_), .A1(mai_mai_n181_), .B0(mai_mai_n182_), .Y(mai_mai_n489_));
  NA2        m467(.A(i_4_), .B(i_8_), .Y(mai_mai_n490_));
  NO2        m468(.A(mai_mai_n489_), .B(i_13_), .Y(mai_mai_n491_));
  NO3        m469(.A(mai_mai_n491_), .B(mai_mai_n488_), .C(mai_mai_n482_), .Y(mai_mai_n492_));
  AOI210     m470(.A0(mai_mai_n119_), .A1(mai_mai_n60_), .B0(i_10_), .Y(mai_mai_n493_));
  AOI210     m471(.A0(mai_mai_n493_), .A1(mai_mai_n210_), .B0(mai_mai_n146_), .Y(mai_mai_n494_));
  OR2        m472(.A(i_6_), .B(i_10_), .Y(mai_mai_n495_));
  NO2        m473(.A(mai_mai_n495_), .B(mai_mai_n23_), .Y(mai_mai_n496_));
  OR3        m474(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n497_));
  NO3        m475(.A(mai_mai_n497_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n498_));
  INV        m476(.A(mai_mai_n178_), .Y(mai_mai_n499_));
  NO2        m477(.A(mai_mai_n498_), .B(mai_mai_n496_), .Y(mai_mai_n500_));
  OA220      m478(.A0(mai_mai_n500_), .A1(mai_mai_n470_), .B0(mai_mai_n494_), .B1(mai_mai_n231_), .Y(mai_mai_n501_));
  AOI210     m479(.A0(mai_mai_n501_), .A1(mai_mai_n492_), .B0(mai_mai_n61_), .Y(mai_mai_n502_));
  NOi21      m480(.An(i_11_), .B(i_7_), .Y(mai_mai_n503_));
  AO210      m481(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n504_));
  NO2        m482(.A(mai_mai_n504_), .B(mai_mai_n503_), .Y(mai_mai_n505_));
  NA2        m483(.A(mai_mai_n505_), .B(mai_mai_n184_), .Y(mai_mai_n506_));
  NA3        m484(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n507_));
  NAi21      m485(.An(mai_mai_n507_), .B(i_11_), .Y(mai_mai_n508_));
  AOI210     m486(.A0(mai_mai_n508_), .A1(mai_mai_n506_), .B0(mai_mai_n61_), .Y(mai_mai_n509_));
  NA2        m487(.A(mai_mai_n79_), .B(mai_mai_n61_), .Y(mai_mai_n510_));
  AO210      m488(.A0(mai_mai_n510_), .A1(mai_mai_n310_), .B0(mai_mai_n40_), .Y(mai_mai_n511_));
  NO3        m489(.A(mai_mai_n222_), .B(mai_mai_n186_), .C(mai_mai_n484_), .Y(mai_mai_n512_));
  OAI210     m490(.A0(mai_mai_n512_), .A1(mai_mai_n201_), .B0(mai_mai_n61_), .Y(mai_mai_n513_));
  NA2        m491(.A(mai_mai_n335_), .B(mai_mai_n31_), .Y(mai_mai_n514_));
  OR2        m492(.A(mai_mai_n186_), .B(mai_mai_n99_), .Y(mai_mai_n515_));
  NA2        m493(.A(mai_mai_n515_), .B(mai_mai_n514_), .Y(mai_mai_n516_));
  NO2        m494(.A(mai_mai_n61_), .B(i_9_), .Y(mai_mai_n517_));
  NO2        m495(.A(mai_mai_n517_), .B(i_4_), .Y(mai_mai_n518_));
  NA2        m496(.A(mai_mai_n518_), .B(mai_mai_n516_), .Y(mai_mai_n519_));
  NO2        m497(.A(i_1_), .B(i_12_), .Y(mai_mai_n520_));
  NA3        m498(.A(mai_mai_n519_), .B(mai_mai_n513_), .C(mai_mai_n511_), .Y(mai_mai_n521_));
  OAI210     m499(.A0(mai_mai_n521_), .A1(mai_mai_n509_), .B0(i_6_), .Y(mai_mai_n522_));
  NO2        m500(.A(mai_mai_n507_), .B(mai_mai_n99_), .Y(mai_mai_n523_));
  NA2        m501(.A(mai_mai_n523_), .B(mai_mai_n471_), .Y(mai_mai_n524_));
  NO2        m502(.A(mai_mai_n210_), .B(mai_mai_n77_), .Y(mai_mai_n525_));
  NO2        m503(.A(mai_mai_n525_), .B(i_11_), .Y(mai_mai_n526_));
  INV        m504(.A(mai_mai_n524_), .Y(mai_mai_n527_));
  NO3        m505(.A(mai_mai_n191_), .B(i_13_), .C(mai_mai_n77_), .Y(mai_mai_n528_));
  NA2        m506(.A(mai_mai_n528_), .B(mai_mai_n517_), .Y(mai_mai_n529_));
  NO3        m507(.A(mai_mai_n495_), .B(mai_mai_n208_), .C(mai_mai_n23_), .Y(mai_mai_n530_));
  AOI210     m508(.A0(i_1_), .A1(mai_mai_n223_), .B0(mai_mai_n530_), .Y(mai_mai_n531_));
  OAI210     m509(.A0(mai_mai_n531_), .A1(mai_mai_n43_), .B0(mai_mai_n529_), .Y(mai_mai_n532_));
  NA3        m510(.A(mai_mai_n438_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n533_));
  INV        m511(.A(i_2_), .Y(mai_mai_n534_));
  NA2        m512(.A(mai_mai_n128_), .B(i_9_), .Y(mai_mai_n535_));
  NA3        m513(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n536_));
  NO2        m514(.A(mai_mai_n45_), .B(i_1_), .Y(mai_mai_n537_));
  NA3        m515(.A(mai_mai_n537_), .B(mai_mai_n230_), .C(mai_mai_n43_), .Y(mai_mai_n538_));
  OAI220     m516(.A0(mai_mai_n538_), .A1(mai_mai_n536_), .B0(mai_mai_n535_), .B1(mai_mai_n534_), .Y(mai_mai_n539_));
  NA3        m517(.A(mai_mai_n517_), .B(mai_mai_n268_), .C(i_6_), .Y(mai_mai_n540_));
  NO2        m518(.A(mai_mai_n540_), .B(mai_mai_n23_), .Y(mai_mai_n541_));
  NO2        m519(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n542_));
  OR2        m520(.A(mai_mai_n541_), .B(mai_mai_n539_), .Y(mai_mai_n543_));
  NO3        m521(.A(mai_mai_n543_), .B(mai_mai_n532_), .C(mai_mai_n527_), .Y(mai_mai_n544_));
  NO2        m522(.A(mai_mai_n210_), .B(mai_mai_n92_), .Y(mai_mai_n545_));
  NO2        m523(.A(mai_mai_n545_), .B(mai_mai_n503_), .Y(mai_mai_n546_));
  NA2        m524(.A(mai_mai_n546_), .B(i_1_), .Y(mai_mai_n547_));
  NO2        m525(.A(mai_mai_n547_), .B(mai_mai_n497_), .Y(mai_mai_n548_));
  NO2        m526(.A(mai_mai_n339_), .B(mai_mai_n77_), .Y(mai_mai_n549_));
  NA2        m527(.A(mai_mai_n548_), .B(mai_mai_n45_), .Y(mai_mai_n550_));
  NA2        m528(.A(i_3_), .B(mai_mai_n172_), .Y(mai_mai_n551_));
  NO2        m529(.A(mai_mai_n551_), .B(mai_mai_n105_), .Y(mai_mai_n552_));
  AN2        m530(.A(mai_mai_n552_), .B(mai_mai_n440_), .Y(mai_mai_n553_));
  NO2        m531(.A(mai_mai_n77_), .B(i_9_), .Y(mai_mai_n554_));
  NA2        m532(.A(i_1_), .B(i_3_), .Y(mai_mai_n555_));
  NO2        m533(.A(mai_mai_n378_), .B(mai_mai_n84_), .Y(mai_mai_n556_));
  INV        m534(.A(mai_mai_n556_), .Y(mai_mai_n557_));
  NO2        m535(.A(mai_mai_n557_), .B(mai_mai_n555_), .Y(mai_mai_n558_));
  NO2        m536(.A(mai_mai_n558_), .B(mai_mai_n553_), .Y(mai_mai_n559_));
  NA4        m537(.A(mai_mai_n559_), .B(mai_mai_n550_), .C(mai_mai_n544_), .D(mai_mai_n522_), .Y(mai_mai_n560_));
  NO3        m538(.A(i_11_), .B(i_3_), .C(i_7_), .Y(mai_mai_n561_));
  NOi21      m539(.An(mai_mai_n561_), .B(i_10_), .Y(mai_mai_n562_));
  OA210      m540(.A0(mai_mai_n562_), .A1(mai_mai_n215_), .B0(mai_mai_n77_), .Y(mai_mai_n563_));
  NA2        m541(.A(i_7_), .B(mai_mai_n302_), .Y(mai_mai_n564_));
  NA3        m542(.A(mai_mai_n401_), .B(mai_mai_n426_), .C(mai_mai_n45_), .Y(mai_mai_n565_));
  NO2        m543(.A(mai_mai_n490_), .B(mai_mai_n77_), .Y(mai_mai_n566_));
  NA2        m544(.A(mai_mai_n566_), .B(mai_mai_n25_), .Y(mai_mai_n567_));
  NA2        m545(.A(mai_mai_n567_), .B(mai_mai_n565_), .Y(mai_mai_n568_));
  OAI210     m546(.A0(mai_mai_n568_), .A1(mai_mai_n563_), .B0(i_1_), .Y(mai_mai_n569_));
  AOI210     m547(.A0(mai_mai_n230_), .A1(mai_mai_n88_), .B0(i_1_), .Y(mai_mai_n570_));
  NO2        m548(.A(mai_mai_n301_), .B(i_2_), .Y(mai_mai_n571_));
  NA2        m549(.A(mai_mai_n571_), .B(mai_mai_n570_), .Y(mai_mai_n572_));
  OAI210     m550(.A0(mai_mai_n540_), .A1(mai_mai_n371_), .B0(mai_mai_n572_), .Y(mai_mai_n573_));
  INV        m551(.A(mai_mai_n573_), .Y(mai_mai_n574_));
  AOI210     m552(.A0(mai_mai_n574_), .A1(mai_mai_n569_), .B0(i_13_), .Y(mai_mai_n575_));
  NA2        m553(.A(mai_mai_n97_), .B(mai_mai_n128_), .Y(mai_mai_n576_));
  AOI220     m554(.A0(mai_mai_n390_), .A1(mai_mai_n146_), .B0(i_2_), .B1(mai_mai_n128_), .Y(mai_mai_n577_));
  OAI210     m555(.A0(mai_mai_n577_), .A1(mai_mai_n43_), .B0(mai_mai_n576_), .Y(mai_mai_n578_));
  AOI220     m556(.A0(i_7_), .A1(mai_mai_n549_), .B0(mai_mai_n215_), .B1(mai_mai_n121_), .Y(mai_mai_n579_));
  NO2        m557(.A(mai_mai_n579_), .B(mai_mai_n40_), .Y(mai_mai_n580_));
  AOI210     m558(.A0(mai_mai_n578_), .A1(mai_mai_n276_), .B0(mai_mai_n580_), .Y(mai_mai_n581_));
  NA2        m559(.A(mai_mai_n318_), .B(mai_mai_n537_), .Y(mai_mai_n582_));
  NO2        m560(.A(mai_mai_n582_), .B(mai_mai_n213_), .Y(mai_mai_n583_));
  AOI210     m561(.A0(mai_mai_n371_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n584_));
  NOi31      m562(.An(mai_mai_n584_), .B(mai_mai_n483_), .C(mai_mai_n43_), .Y(mai_mai_n585_));
  NA2        m563(.A(mai_mai_n118_), .B(i_13_), .Y(mai_mai_n586_));
  NO2        m564(.A(mai_mai_n536_), .B(mai_mai_n105_), .Y(mai_mai_n587_));
  INV        m565(.A(mai_mai_n587_), .Y(mai_mai_n588_));
  OAI220     m566(.A0(mai_mai_n588_), .A1(mai_mai_n65_), .B0(mai_mai_n586_), .B1(mai_mai_n570_), .Y(mai_mai_n589_));
  NA2        m567(.A(i_3_), .B(i_7_), .Y(mai_mai_n590_));
  NO3        m568(.A(mai_mai_n395_), .B(mai_mai_n210_), .C(mai_mai_n77_), .Y(mai_mai_n591_));
  NA2        m569(.A(mai_mai_n591_), .B(mai_mai_n590_), .Y(mai_mai_n592_));
  AOI220     m570(.A0(mai_mai_n318_), .A1(mai_mai_n537_), .B0(mai_mai_n83_), .B1(mai_mai_n93_), .Y(mai_mai_n593_));
  OAI220     m571(.A0(mai_mai_n593_), .A1(mai_mai_n487_), .B0(mai_mai_n592_), .B1(mai_mai_n499_), .Y(mai_mai_n594_));
  NO4        m572(.A(mai_mai_n594_), .B(mai_mai_n589_), .C(mai_mai_n585_), .D(mai_mai_n583_), .Y(mai_mai_n595_));
  OR2        m573(.A(i_11_), .B(i_6_), .Y(mai_mai_n596_));
  NA2        m574(.A(mai_mai_n486_), .B(i_7_), .Y(mai_mai_n597_));
  AOI210     m575(.A0(mai_mai_n597_), .A1(mai_mai_n588_), .B0(mai_mai_n596_), .Y(mai_mai_n598_));
  NA3        m576(.A(mai_mai_n335_), .B(i_10_), .C(mai_mai_n88_), .Y(mai_mai_n599_));
  NA2        m577(.A(mai_mai_n526_), .B(i_13_), .Y(mai_mai_n600_));
  NAi21      m578(.An(i_11_), .B(i_12_), .Y(mai_mai_n601_));
  NOi41      m579(.An(mai_mai_n101_), .B(mai_mai_n601_), .C(i_13_), .D(mai_mai_n77_), .Y(mai_mai_n602_));
  NO2        m580(.A(mai_mai_n471_), .B(mai_mai_n490_), .Y(mai_mai_n603_));
  AOI210     m581(.A0(mai_mai_n603_), .A1(mai_mai_n266_), .B0(mai_mai_n602_), .Y(mai_mai_n604_));
  NA3        m582(.A(mai_mai_n604_), .B(mai_mai_n600_), .C(mai_mai_n599_), .Y(mai_mai_n605_));
  OAI210     m583(.A0(mai_mai_n605_), .A1(mai_mai_n598_), .B0(mai_mai_n61_), .Y(mai_mai_n606_));
  NO2        m584(.A(i_2_), .B(i_12_), .Y(mai_mai_n607_));
  NA2        m585(.A(mai_mai_n300_), .B(mai_mai_n607_), .Y(mai_mai_n608_));
  NO3        m586(.A(i_9_), .B(mai_mai_n316_), .C(mai_mai_n486_), .Y(mai_mai_n609_));
  NA2        m587(.A(mai_mai_n609_), .B(mai_mai_n300_), .Y(mai_mai_n610_));
  NO2        m588(.A(mai_mai_n119_), .B(i_2_), .Y(mai_mai_n611_));
  NA2        m589(.A(mai_mai_n611_), .B(mai_mai_n520_), .Y(mai_mai_n612_));
  NA3        m590(.A(mai_mai_n612_), .B(mai_mai_n610_), .C(mai_mai_n608_), .Y(mai_mai_n613_));
  NA3        m591(.A(mai_mai_n613_), .B(mai_mai_n44_), .C(mai_mai_n200_), .Y(mai_mai_n614_));
  NA4        m592(.A(mai_mai_n614_), .B(mai_mai_n606_), .C(mai_mai_n595_), .D(mai_mai_n581_), .Y(mai_mai_n615_));
  OR4        m593(.A(mai_mai_n615_), .B(mai_mai_n575_), .C(mai_mai_n560_), .D(mai_mai_n502_), .Y(mai5));
  AOI210     m594(.A0(mai_mai_n546_), .A1(mai_mai_n233_), .B0(mai_mai_n341_), .Y(mai_mai_n617_));
  AO210      m595(.A0(mai_mai_n24_), .A1(i_10_), .B0(mai_mai_n216_), .Y(mai_mai_n618_));
  NA3        m596(.A(mai_mai_n618_), .B(mai_mai_n607_), .C(mai_mai_n99_), .Y(mai_mai_n619_));
  NO2        m597(.A(mai_mai_n487_), .B(i_11_), .Y(mai_mai_n620_));
  NA2        m598(.A(mai_mai_n80_), .B(mai_mai_n620_), .Y(mai_mai_n621_));
  NA3        m599(.A(mai_mai_n621_), .B(mai_mai_n619_), .C(mai_mai_n617_), .Y(mai_mai_n622_));
  NO3        m600(.A(i_11_), .B(mai_mai_n210_), .C(i_13_), .Y(mai_mai_n623_));
  NO2        m601(.A(mai_mai_n115_), .B(mai_mai_n23_), .Y(mai_mai_n624_));
  NA2        m602(.A(i_12_), .B(i_8_), .Y(mai_mai_n625_));
  OAI210     m603(.A0(mai_mai_n45_), .A1(i_3_), .B0(mai_mai_n625_), .Y(mai_mai_n626_));
  INV        m604(.A(mai_mai_n370_), .Y(mai_mai_n627_));
  AOI220     m605(.A0(mai_mai_n268_), .A1(mai_mai_n464_), .B0(mai_mai_n626_), .B1(mai_mai_n624_), .Y(mai_mai_n628_));
  INV        m606(.A(mai_mai_n628_), .Y(mai_mai_n629_));
  NO2        m607(.A(mai_mai_n629_), .B(mai_mai_n622_), .Y(mai_mai_n630_));
  INV        m608(.A(mai_mai_n154_), .Y(mai_mai_n631_));
  INV        m609(.A(mai_mai_n215_), .Y(mai_mai_n632_));
  OAI210     m610(.A0(mai_mai_n571_), .A1(mai_mai_n372_), .B0(mai_mai_n101_), .Y(mai_mai_n633_));
  AOI210     m611(.A0(mai_mai_n633_), .A1(mai_mai_n632_), .B0(mai_mai_n631_), .Y(mai_mai_n634_));
  NO2        m612(.A(mai_mai_n378_), .B(mai_mai_n26_), .Y(mai_mai_n635_));
  NO2        m613(.A(mai_mai_n635_), .B(mai_mai_n343_), .Y(mai_mai_n636_));
  NA2        m614(.A(mai_mai_n636_), .B(i_2_), .Y(mai_mai_n637_));
  INV        m615(.A(mai_mai_n637_), .Y(mai_mai_n638_));
  AOI210     m616(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n340_), .Y(mai_mai_n639_));
  AOI210     m617(.A0(mai_mai_n639_), .A1(mai_mai_n638_), .B0(mai_mai_n634_), .Y(mai_mai_n640_));
  NO2        m618(.A(mai_mai_n169_), .B(mai_mai_n116_), .Y(mai_mai_n641_));
  NA2        m619(.A(mai_mai_n641_), .B(i_2_), .Y(mai_mai_n642_));
  INV        m620(.A(mai_mai_n155_), .Y(mai_mai_n643_));
  NO3        m621(.A(mai_mai_n504_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n644_));
  AOI210     m622(.A0(mai_mai_n643_), .A1(mai_mai_n80_), .B0(mai_mai_n644_), .Y(mai_mai_n645_));
  AOI210     m623(.A0(mai_mai_n645_), .A1(mai_mai_n642_), .B0(mai_mai_n172_), .Y(mai_mai_n646_));
  OA210      m624(.A0(mai_mai_n505_), .A1(mai_mai_n117_), .B0(i_13_), .Y(mai_mai_n647_));
  NA2        m625(.A(mai_mai_n178_), .B(mai_mai_n181_), .Y(mai_mai_n648_));
  INV        m626(.A(mai_mai_n137_), .Y(mai_mai_n649_));
  AOI210     m627(.A0(mai_mai_n649_), .A1(mai_mai_n648_), .B0(mai_mai_n304_), .Y(mai_mai_n650_));
  NA3        m628(.A(i_2_), .B(mai_mai_n262_), .C(mai_mai_n115_), .Y(mai_mai_n651_));
  INV        m629(.A(mai_mai_n651_), .Y(mai_mai_n652_));
  NO4        m630(.A(mai_mai_n652_), .B(mai_mai_n650_), .C(mai_mai_n647_), .D(mai_mai_n646_), .Y(mai_mai_n653_));
  NA2        m631(.A(mai_mai_n464_), .B(mai_mai_n28_), .Y(mai_mai_n654_));
  NA2        m632(.A(mai_mai_n623_), .B(mai_mai_n239_), .Y(mai_mai_n655_));
  NA2        m633(.A(mai_mai_n655_), .B(mai_mai_n654_), .Y(mai_mai_n656_));
  NO2        m634(.A(mai_mai_n60_), .B(i_12_), .Y(mai_mai_n657_));
  NO2        m635(.A(mai_mai_n657_), .B(mai_mai_n117_), .Y(mai_mai_n658_));
  NO2        m636(.A(mai_mai_n658_), .B(mai_mai_n484_), .Y(mai_mai_n659_));
  AOI220     m637(.A0(mai_mai_n659_), .A1(mai_mai_n36_), .B0(mai_mai_n656_), .B1(mai_mai_n45_), .Y(mai_mai_n660_));
  NA4        m638(.A(mai_mai_n660_), .B(mai_mai_n653_), .C(mai_mai_n640_), .D(mai_mai_n630_), .Y(mai6));
  NO2        m639(.A(i_9_), .B(mai_mai_n871_), .Y(mai_mai_n662_));
  OAI210     m640(.A0(mai_mai_n67_), .A1(mai_mai_n662_), .B0(mai_mai_n611_), .Y(mai_mai_n663_));
  NA4        m641(.A(mai_mai_n322_), .B(mai_mai_n400_), .C(mai_mai_n65_), .D(mai_mai_n92_), .Y(mai_mai_n664_));
  INV        m642(.A(mai_mai_n664_), .Y(mai_mai_n665_));
  NO2        m643(.A(mai_mai_n196_), .B(mai_mai_n403_), .Y(mai_mai_n666_));
  NO2        m644(.A(i_11_), .B(i_9_), .Y(mai_mai_n667_));
  NO2        m645(.A(mai_mai_n665_), .B(mai_mai_n274_), .Y(mai_mai_n668_));
  AO210      m646(.A0(mai_mai_n668_), .A1(mai_mai_n663_), .B0(i_12_), .Y(mai_mai_n669_));
  NA2        m647(.A(mai_mai_n305_), .B(mai_mai_n278_), .Y(mai_mai_n670_));
  NA2        m648(.A(mai_mai_n471_), .B(mai_mai_n61_), .Y(mai_mai_n671_));
  NA2        m649(.A(mai_mai_n562_), .B(mai_mai_n65_), .Y(mai_mai_n672_));
  NA4        m650(.A(mai_mai_n510_), .B(mai_mai_n672_), .C(mai_mai_n671_), .D(mai_mai_n670_), .Y(mai_mai_n673_));
  INV        m651(.A(mai_mai_n175_), .Y(mai_mai_n674_));
  AOI220     m652(.A0(mai_mai_n674_), .A1(mai_mai_n667_), .B0(mai_mai_n673_), .B1(mai_mai_n67_), .Y(mai_mai_n675_));
  NA2        m653(.A(mai_mai_n864_), .B(mai_mai_n657_), .Y(mai_mai_n676_));
  AOI210     m654(.A0(mai_mai_n676_), .A1(mai_mai_n424_), .B0(mai_mai_n164_), .Y(mai_mai_n677_));
  NO2        m655(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n678_));
  NA3        m656(.A(mai_mai_n678_), .B(mai_mai_n394_), .C(mai_mai_n322_), .Y(mai_mai_n679_));
  NA2        m657(.A(mai_mai_n455_), .B(mai_mai_n454_), .Y(mai_mai_n680_));
  NA2        m658(.A(mai_mai_n680_), .B(mai_mai_n679_), .Y(mai_mai_n681_));
  OR2        m659(.A(mai_mai_n681_), .B(mai_mai_n677_), .Y(mai_mai_n682_));
  NO2        m660(.A(i_11_), .B(i_2_), .Y(mai_mai_n683_));
  NA2        m661(.A(mai_mai_n47_), .B(mai_mai_n37_), .Y(mai_mai_n684_));
  NA2        m662(.A(mai_mai_n867_), .B(mai_mai_n683_), .Y(mai_mai_n685_));
  NA3        m663(.A(mai_mai_n284_), .B(mai_mai_n220_), .C(i_7_), .Y(mai_mai_n686_));
  OR2        m664(.A(mai_mai_n627_), .B(mai_mai_n36_), .Y(mai_mai_n687_));
  NA3        m665(.A(mai_mai_n687_), .B(mai_mai_n686_), .C(mai_mai_n685_), .Y(mai_mai_n688_));
  AOI220     m666(.A0(mai_mai_n866_), .A1(mai_mai_n454_), .B0(mai_mai_n666_), .B1(mai_mai_n590_), .Y(mai_mai_n689_));
  NA3        m667(.A(mai_mai_n304_), .B(mai_mai_n211_), .C(mai_mai_n136_), .Y(mai_mai_n690_));
  NA3        m668(.A(mai_mai_n690_), .B(mai_mai_n689_), .C(mai_mai_n489_), .Y(mai_mai_n691_));
  NA3        m669(.A(mai_mai_n426_), .B(mai_mai_n401_), .C(mai_mai_n194_), .Y(mai_mai_n692_));
  AOI210     m670(.A0(mai_mai_n372_), .A1(mai_mai_n370_), .B0(mai_mai_n453_), .Y(mai_mai_n693_));
  OAI210     m671(.A0(mai_mai_n870_), .A1(mai_mai_n102_), .B0(mai_mai_n334_), .Y(mai_mai_n694_));
  INV        m672(.A(mai_mai_n476_), .Y(mai_mai_n695_));
  NA3        m673(.A(mai_mai_n695_), .B(mai_mai_n273_), .C(i_7_), .Y(mai_mai_n696_));
  NA4        m674(.A(mai_mai_n696_), .B(mai_mai_n694_), .C(mai_mai_n693_), .D(mai_mai_n692_), .Y(mai_mai_n697_));
  NO4        m675(.A(mai_mai_n697_), .B(mai_mai_n691_), .C(mai_mai_n688_), .D(mai_mai_n682_), .Y(mai_mai_n698_));
  NA4        m676(.A(mai_mai_n698_), .B(mai_mai_n675_), .C(mai_mai_n669_), .D(mai_mai_n312_), .Y(mai3));
  NO2        m677(.A(i_11_), .B(mai_mai_n210_), .Y(mai_mai_n700_));
  NA2        m678(.A(mai_mai_n250_), .B(mai_mai_n700_), .Y(mai_mai_n701_));
  NO2        m679(.A(mai_mai_n701_), .B(mai_mai_n172_), .Y(mai_mai_n702_));
  AN2        m680(.A(mai_mai_n702_), .B(mai_mai_n156_), .Y(mai_mai_n703_));
  NA3        m681(.A(mai_mai_n690_), .B(mai_mai_n489_), .C(mai_mai_n303_), .Y(mai_mai_n704_));
  NA2        m682(.A(mai_mai_n704_), .B(mai_mai_n39_), .Y(mai_mai_n705_));
  NO3        m683(.A(mai_mai_n515_), .B(mai_mai_n378_), .C(mai_mai_n121_), .Y(mai_mai_n706_));
  NA2        m684(.A(mai_mai_n335_), .B(mai_mai_n44_), .Y(mai_mai_n707_));
  AN2        m685(.A(mai_mai_n377_), .B(mai_mai_n53_), .Y(mai_mai_n708_));
  NO2        m686(.A(mai_mai_n708_), .B(mai_mai_n706_), .Y(mai_mai_n709_));
  AOI210     m687(.A0(mai_mai_n709_), .A1(mai_mai_n705_), .B0(mai_mai_n47_), .Y(mai_mai_n710_));
  NOi21      m688(.An(i_5_), .B(i_9_), .Y(mai_mai_n711_));
  NA2        m689(.A(mai_mai_n711_), .B(mai_mai_n368_), .Y(mai_mai_n712_));
  NO3        m690(.A(mai_mai_n336_), .B(mai_mai_n230_), .C(mai_mai_n67_), .Y(mai_mai_n713_));
  INV        m691(.A(mai_mai_n713_), .Y(mai_mai_n714_));
  NO2        m692(.A(mai_mai_n714_), .B(i_4_), .Y(mai_mai_n715_));
  NO3        m693(.A(mai_mai_n715_), .B(mai_mai_n710_), .C(mai_mai_n703_), .Y(mai_mai_n716_));
  NA2        m694(.A(mai_mai_n266_), .B(mai_mai_n120_), .Y(mai_mai_n717_));
  NAi21      m695(.An(mai_mai_n147_), .B(i_5_), .Y(mai_mai_n718_));
  NO2        m696(.A(mai_mai_n717_), .B(mai_mai_n329_), .Y(mai_mai_n719_));
  INV        m697(.A(mai_mai_n719_), .Y(mai_mai_n720_));
  NA2        m698(.A(mai_mai_n461_), .B(i_0_), .Y(mai_mai_n721_));
  NO3        m699(.A(mai_mai_n721_), .B(mai_mai_n317_), .C(mai_mai_n80_), .Y(mai_mai_n722_));
  NO3        m700(.A(mai_mai_n476_), .B(mai_mai_n191_), .C(mai_mai_n340_), .Y(mai_mai_n723_));
  AOI210     m701(.A0(mai_mai_n723_), .A1(i_11_), .B0(mai_mai_n722_), .Y(mai_mai_n724_));
  NA2        m702(.A(mai_mai_n623_), .B(mai_mai_n274_), .Y(mai_mai_n725_));
  NO2        m703(.A(mai_mai_n401_), .B(mai_mai_n56_), .Y(mai_mai_n726_));
  NO2        m704(.A(mai_mai_n726_), .B(mai_mai_n725_), .Y(mai_mai_n727_));
  NO2        m705(.A(mai_mai_n218_), .B(mai_mai_n138_), .Y(mai_mai_n728_));
  INV        m706(.A(mai_mai_n439_), .Y(mai_mai_n729_));
  NO4        m707(.A(mai_mai_n105_), .B(mai_mai_n56_), .C(mai_mai_n551_), .D(i_5_), .Y(mai_mai_n730_));
  AO220      m708(.A0(mai_mai_n730_), .A1(mai_mai_n729_), .B0(mai_mai_n728_), .B1(i_6_), .Y(mai_mai_n731_));
  NA2        m709(.A(mai_mai_n167_), .B(mai_mai_n181_), .Y(mai_mai_n732_));
  NO2        m710(.A(mai_mai_n732_), .B(mai_mai_n725_), .Y(mai_mai_n733_));
  NO3        m711(.A(mai_mai_n733_), .B(mai_mai_n731_), .C(mai_mai_n727_), .Y(mai_mai_n734_));
  NA3        m712(.A(mai_mai_n734_), .B(mai_mai_n724_), .C(mai_mai_n720_), .Y(mai_mai_n735_));
  NA2        m713(.A(i_11_), .B(i_9_), .Y(mai_mai_n736_));
  NO2        m714(.A(mai_mai_n47_), .B(i_7_), .Y(mai_mai_n737_));
  NA2        m715(.A(mai_mai_n326_), .B(mai_mai_n159_), .Y(mai_mai_n738_));
  NAi31      m716(.An(mai_mai_n227_), .B(mai_mai_n738_), .C(mai_mai_n145_), .Y(mai_mai_n739_));
  NO2        m717(.A(mai_mai_n157_), .B(i_0_), .Y(mai_mai_n740_));
  NA2        m718(.A(mai_mai_n394_), .B(mai_mai_n206_), .Y(mai_mai_n741_));
  OAI220     m719(.A0(i_12_), .A1(mai_mai_n712_), .B0(mai_mai_n741_), .B1(mai_mai_n157_), .Y(mai_mai_n742_));
  NO2        m720(.A(mai_mai_n742_), .B(mai_mai_n739_), .Y(mai_mai_n743_));
  NA2        m721(.A(mai_mai_n542_), .B(mai_mai_n112_), .Y(mai_mai_n744_));
  NO2        m722(.A(i_6_), .B(mai_mai_n744_), .Y(mai_mai_n745_));
  AOI210     m723(.A0(mai_mai_n371_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n746_));
  NA2        m724(.A(mai_mai_n154_), .B(mai_mai_n94_), .Y(mai_mai_n747_));
  NOi32      m725(.An(mai_mai_n746_), .Bn(mai_mai_n167_), .C(mai_mai_n747_), .Y(mai_mai_n748_));
  NO2        m726(.A(mai_mai_n869_), .B(mai_mai_n707_), .Y(mai_mai_n749_));
  NO3        m727(.A(mai_mai_n749_), .B(mai_mai_n748_), .C(mai_mai_n745_), .Y(mai_mai_n750_));
  NOi21      m728(.An(i_7_), .B(i_5_), .Y(mai_mai_n751_));
  NOi31      m729(.An(mai_mai_n751_), .B(i_0_), .C(mai_mai_n601_), .Y(mai_mai_n752_));
  NA3        m730(.A(mai_mai_n752_), .B(mai_mai_n316_), .C(i_6_), .Y(mai_mai_n753_));
  BUFFER     m731(.A(mai_mai_n753_), .Y(mai_mai_n754_));
  NA3        m732(.A(mai_mai_n754_), .B(mai_mai_n750_), .C(mai_mai_n743_), .Y(mai_mai_n755_));
  OA210      m733(.A0(mai_mai_n394_), .A1(mai_mai_n198_), .B0(mai_mai_n393_), .Y(mai_mai_n756_));
  NA3        m734(.A(mai_mai_n393_), .B(mai_mai_n335_), .C(mai_mai_n44_), .Y(mai_mai_n757_));
  OAI210     m735(.A0(mai_mai_n718_), .A1(i_6_), .B0(mai_mai_n757_), .Y(mai_mai_n758_));
  INV        m736(.A(mai_mai_n166_), .Y(mai_mai_n759_));
  AOI220     m737(.A0(mai_mai_n759_), .A1(mai_mai_n394_), .B0(mai_mai_n758_), .B1(mai_mai_n67_), .Y(mai_mai_n760_));
  NA2        m738(.A(mai_mai_n314_), .B(mai_mai_n525_), .Y(mai_mai_n761_));
  NA2        m739(.A(mai_mai_n84_), .B(mai_mai_n43_), .Y(mai_mai_n762_));
  NO2        m740(.A(mai_mai_n69_), .B(mai_mai_n625_), .Y(mai_mai_n763_));
  NA2        m741(.A(mai_mai_n763_), .B(mai_mai_n762_), .Y(mai_mai_n764_));
  AOI210     m742(.A0(mai_mai_n764_), .A1(mai_mai_n761_), .B0(mai_mai_n46_), .Y(mai_mai_n765_));
  NO3        m743(.A(mai_mai_n476_), .B(i_0_), .C(mai_mai_n24_), .Y(mai_mai_n766_));
  NO2        m744(.A(mai_mai_n445_), .B(mai_mai_n766_), .Y(mai_mai_n767_));
  NAi21      m745(.An(i_9_), .B(i_5_), .Y(mai_mai_n768_));
  NO2        m746(.A(mai_mai_n485_), .B(mai_mai_n96_), .Y(mai_mai_n769_));
  NA2        m747(.A(mai_mai_n769_), .B(i_0_), .Y(mai_mai_n770_));
  OAI220     m748(.A0(mai_mai_n770_), .A1(mai_mai_n77_), .B0(mai_mai_n767_), .B1(mai_mai_n155_), .Y(mai_mai_n771_));
  NO3        m749(.A(mai_mai_n771_), .B(mai_mai_n765_), .C(mai_mai_n427_), .Y(mai_mai_n772_));
  NA2        m750(.A(mai_mai_n772_), .B(mai_mai_n760_), .Y(mai_mai_n773_));
  NO3        m751(.A(mai_mai_n773_), .B(mai_mai_n755_), .C(mai_mai_n735_), .Y(mai_mai_n774_));
  NO2        m752(.A(i_0_), .B(mai_mai_n601_), .Y(mai_mai_n775_));
  NA2        m753(.A(mai_mai_n67_), .B(mai_mai_n43_), .Y(mai_mai_n776_));
  NO3        m754(.A(mai_mai_n96_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n777_));
  AO220      m755(.A0(mai_mai_n777_), .A1(mai_mai_n43_), .B0(mai_mai_n775_), .B1(mai_mai_n156_), .Y(mai_mai_n778_));
  AOI210     m756(.A0(mai_mai_n671_), .A1(mai_mai_n564_), .B0(mai_mai_n747_), .Y(mai_mai_n779_));
  AOI210     m757(.A0(mai_mai_n778_), .A1(mai_mai_n283_), .B0(mai_mai_n779_), .Y(mai_mai_n780_));
  NA3        m758(.A(mai_mai_n135_), .B(mai_mai_n554_), .C(mai_mai_n67_), .Y(mai_mai_n781_));
  NA3        m759(.A(i_6_), .B(i_2_), .C(mai_mai_n47_), .Y(mai_mai_n782_));
  NA2        m760(.A(mai_mai_n700_), .B(i_9_), .Y(mai_mai_n783_));
  AOI210     m761(.A0(mai_mai_n782_), .A1(mai_mai_n412_), .B0(mai_mai_n783_), .Y(mai_mai_n784_));
  NA2        m762(.A(mai_mai_n214_), .B(mai_mai_n205_), .Y(mai_mai_n785_));
  AOI210     m763(.A0(mai_mai_n785_), .A1(mai_mai_n721_), .B0(mai_mai_n138_), .Y(mai_mai_n786_));
  NO2        m764(.A(mai_mai_n786_), .B(mai_mai_n784_), .Y(mai_mai_n787_));
  NA3        m765(.A(mai_mai_n787_), .B(mai_mai_n781_), .C(mai_mai_n780_), .Y(mai_mai_n788_));
  NA3        m766(.A(mai_mai_n39_), .B(mai_mai_n28_), .C(mai_mai_n43_), .Y(mai_mai_n789_));
  NA2        m767(.A(mai_mai_n737_), .B(mai_mai_n404_), .Y(mai_mai_n790_));
  AOI210     m768(.A0(mai_mai_n789_), .A1(mai_mai_n147_), .B0(mai_mai_n790_), .Y(mai_mai_n791_));
  INV        m769(.A(mai_mai_n791_), .Y(mai_mai_n792_));
  NO3        m770(.A(mai_mai_n187_), .B(mai_mai_n315_), .C(i_0_), .Y(mai_mai_n793_));
  OAI210     m771(.A0(mai_mai_n793_), .A1(mai_mai_n70_), .B0(i_13_), .Y(mai_mai_n794_));
  NA2        m772(.A(mai_mai_n794_), .B(mai_mai_n792_), .Y(mai_mai_n795_));
  NO2        m773(.A(mai_mai_n213_), .B(mai_mai_n84_), .Y(mai_mai_n796_));
  NA2        m774(.A(mai_mai_n796_), .B(mai_mai_n775_), .Y(mai_mai_n797_));
  NA2        m775(.A(mai_mai_n751_), .B(mai_mai_n404_), .Y(mai_mai_n798_));
  INV        m776(.A(mai_mai_n158_), .Y(mai_mai_n799_));
  OA220      m777(.A0(mai_mai_n799_), .A1(mai_mai_n798_), .B0(mai_mai_n797_), .B1(i_5_), .Y(mai_mai_n800_));
  AOI210     m778(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n157_), .Y(mai_mai_n801_));
  NA2        m779(.A(mai_mai_n801_), .B(mai_mai_n756_), .Y(mai_mai_n802_));
  NA2        m780(.A(mai_mai_n402_), .B(mai_mai_n391_), .Y(mai_mai_n803_));
  INV        m781(.A(mai_mai_n803_), .Y(mai_mai_n804_));
  NA3        m782(.A(mai_mai_n322_), .B(mai_mai_n277_), .C(mai_mai_n197_), .Y(mai_mai_n805_));
  INV        m783(.A(mai_mai_n805_), .Y(mai_mai_n806_));
  NOi31      m784(.An(mai_mai_n321_), .B(mai_mai_n776_), .C(mai_mai_n212_), .Y(mai_mai_n807_));
  NO3        m785(.A(mai_mai_n736_), .B(mai_mai_n194_), .C(mai_mai_n169_), .Y(mai_mai_n808_));
  NO3        m786(.A(mai_mai_n808_), .B(mai_mai_n807_), .C(mai_mai_n806_), .Y(mai_mai_n809_));
  NA4        m787(.A(mai_mai_n809_), .B(mai_mai_n804_), .C(mai_mai_n802_), .D(mai_mai_n800_), .Y(mai_mai_n810_));
  NO2        m788(.A(mai_mai_n77_), .B(i_5_), .Y(mai_mai_n811_));
  NA3        m789(.A(mai_mai_n700_), .B(mai_mai_n100_), .C(mai_mai_n115_), .Y(mai_mai_n812_));
  INV        m790(.A(mai_mai_n812_), .Y(mai_mai_n813_));
  NA2        m791(.A(mai_mai_n813_), .B(mai_mai_n811_), .Y(mai_mai_n814_));
  NA2        m792(.A(mai_mai_n262_), .B(i_5_), .Y(mai_mai_n815_));
  NO4        m793(.A(mai_mai_n212_), .B(mai_mai_n187_), .C(i_0_), .D(i_12_), .Y(mai_mai_n816_));
  AOI220     m794(.A0(mai_mai_n816_), .A1(mai_mai_n863_), .B0(mai_mai_n665_), .B1(mai_mai_n158_), .Y(mai_mai_n817_));
  BUFFER     m795(.A(mai_mai_n138_), .Y(mai_mai_n818_));
  NO4        m796(.A(mai_mai_n818_), .B(i_12_), .C(mai_mai_n533_), .D(mai_mai_n121_), .Y(mai_mai_n819_));
  NA2        m797(.A(mai_mai_n819_), .B(mai_mai_n194_), .Y(mai_mai_n820_));
  NA2        m798(.A(mai_mai_n751_), .B(mai_mai_n390_), .Y(mai_mai_n821_));
  OAI220     m799(.A0(i_6_), .A1(mai_mai_n815_), .B0(mai_mai_n821_), .B1(i_1_), .Y(mai_mai_n822_));
  NA2        m800(.A(mai_mai_n822_), .B(mai_mai_n740_), .Y(mai_mai_n823_));
  NA4        m801(.A(mai_mai_n823_), .B(mai_mai_n820_), .C(mai_mai_n817_), .D(mai_mai_n814_), .Y(mai_mai_n824_));
  NO4        m802(.A(mai_mai_n824_), .B(mai_mai_n810_), .C(mai_mai_n795_), .D(mai_mai_n788_), .Y(mai_mai_n825_));
  OAI210     m803(.A0(mai_mai_n683_), .A1(mai_mai_n678_), .B0(mai_mai_n37_), .Y(mai_mai_n826_));
  NA2        m804(.A(mai_mai_n826_), .B(mai_mai_n494_), .Y(mai_mai_n827_));
  NA2        m805(.A(mai_mai_n827_), .B(mai_mai_n184_), .Y(mai_mai_n828_));
  NA2        m806(.A(mai_mai_n165_), .B(mai_mai_n167_), .Y(mai_mai_n829_));
  OAI210     m807(.A0(mai_mai_n498_), .A1(mai_mai_n496_), .B0(mai_mai_n268_), .Y(mai_mai_n830_));
  NA2        m808(.A(mai_mai_n830_), .B(mai_mai_n829_), .Y(mai_mai_n831_));
  NO2        m809(.A(mai_mai_n382_), .B(mai_mai_n230_), .Y(mai_mai_n832_));
  NO2        m810(.A(mai_mai_n832_), .B(mai_mai_n723_), .Y(mai_mai_n833_));
  INV        m811(.A(mai_mai_n833_), .Y(mai_mai_n834_));
  AOI210     m812(.A0(mai_mai_n831_), .A1(mai_mai_n47_), .B0(mai_mai_n834_), .Y(mai_mai_n835_));
  AOI210     m813(.A0(mai_mai_n835_), .A1(mai_mai_n828_), .B0(mai_mai_n67_), .Y(mai_mai_n836_));
  NO2        m814(.A(mai_mai_n456_), .B(mai_mai_n311_), .Y(mai_mai_n837_));
  NO2        m815(.A(mai_mai_n837_), .B(mai_mai_n631_), .Y(mai_mai_n838_));
  AOI210     m816(.A0(mai_mai_n801_), .A1(mai_mai_n737_), .B0(mai_mai_n752_), .Y(mai_mai_n839_));
  NO2        m817(.A(mai_mai_n839_), .B(mai_mai_n555_), .Y(mai_mai_n840_));
  INV        m818(.A(mai_mai_n55_), .Y(mai_mai_n841_));
  NA2        m819(.A(mai_mai_n841_), .B(mai_mai_n70_), .Y(mai_mai_n842_));
  NO2        m820(.A(mai_mai_n842_), .B(mai_mai_n210_), .Y(mai_mai_n843_));
  NO2        m821(.A(mai_mai_n843_), .B(mai_mai_n840_), .Y(mai_mai_n844_));
  OAI210     m822(.A0(mai_mai_n232_), .A1(mai_mai_n143_), .B0(mai_mai_n80_), .Y(mai_mai_n845_));
  NO2        m823(.A(mai_mai_n845_), .B(i_11_), .Y(mai_mai_n846_));
  NA2        m824(.A(mai_mai_n746_), .B(mai_mai_n184_), .Y(mai_mai_n847_));
  NA2        m825(.A(i_0_), .B(i_5_), .Y(mai_mai_n848_));
  AOI210     m826(.A0(mai_mai_n847_), .A1(mai_mai_n648_), .B0(mai_mai_n848_), .Y(mai_mai_n849_));
  NO3        m827(.A(mai_mai_n57_), .B(mai_mai_n56_), .C(i_4_), .Y(mai_mai_n850_));
  NA2        m828(.A(mai_mai_n871_), .B(mai_mai_n850_), .Y(mai_mai_n851_));
  NO2        m829(.A(mai_mai_n851_), .B(mai_mai_n601_), .Y(mai_mai_n852_));
  NO3        m830(.A(mai_mai_n768_), .B(i_11_), .C(mai_mai_n217_), .Y(mai_mai_n853_));
  NO2        m831(.A(mai_mai_n853_), .B(mai_mai_n453_), .Y(mai_mai_n854_));
  INV        m832(.A(mai_mai_n294_), .Y(mai_mai_n855_));
  AOI210     m833(.A0(mai_mai_n855_), .A1(mai_mai_n854_), .B0(mai_mai_n40_), .Y(mai_mai_n856_));
  NO4        m834(.A(mai_mai_n856_), .B(mai_mai_n852_), .C(mai_mai_n849_), .D(mai_mai_n846_), .Y(mai_mai_n857_));
  OAI210     m835(.A0(mai_mai_n844_), .A1(i_4_), .B0(mai_mai_n857_), .Y(mai_mai_n858_));
  NO3        m836(.A(mai_mai_n858_), .B(mai_mai_n838_), .C(mai_mai_n836_), .Y(mai_mai_n859_));
  NA4        m837(.A(mai_mai_n859_), .B(mai_mai_n825_), .C(mai_mai_n774_), .D(mai_mai_n716_), .Y(mai4));
  INV        m838(.A(mai_mai_n213_), .Y(mai_mai_n863_));
  INV        m839(.A(i_9_), .Y(mai_mai_n864_));
  INV        m840(.A(mai_mai_n213_), .Y(mai_mai_n865_));
  INV        m841(.A(i_11_), .Y(mai_mai_n866_));
  INV        m842(.A(mai_mai_n684_), .Y(mai_mai_n867_));
  INV        m843(.A(i_6_), .Y(mai_mai_n868_));
  INV        m844(.A(mai_mai_n274_), .Y(mai_mai_n869_));
  INV        m845(.A(mai_mai_n495_), .Y(mai_mai_n870_));
  INV        m846(.A(i_5_), .Y(mai_mai_n871_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NOi21      u0016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u0017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u0018(.A(men_men_n36_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n35_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NO2        u0026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u0027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  OAI210     u0028(.A0(men_men_n50_), .A1(i_3_), .B0(men_men_n48_), .Y(men_men_n51_));
  AOI210     u0029(.A0(men_men_n51_), .A1(men_men_n47_), .B0(men_men_n46_), .Y(men_men_n52_));
  NA2        u0030(.A(i_0_), .B(i_2_), .Y(men_men_n53_));
  NA2        u0031(.A(i_7_), .B(i_9_), .Y(men_men_n54_));
  NO2        u0032(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n52_), .B(men_men_n45_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_10_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(i_6_), .Y(men_men_n67_));
  NAi31      u0045(.An(men_men_n67_), .B(men_men_n65_), .C(men_men_n61_), .Y(men_men_n68_));
  NA2        u0046(.A(men_men_n50_), .B(i_2_), .Y(men_men_n69_));
  AOI210     u0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n70_));
  NA2        u0048(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n25_), .Y(men_men_n72_));
  INV        u0050(.A(i_0_), .Y(men_men_n73_));
  NAi21      u0051(.An(i_5_), .B(i_10_), .Y(men_men_n74_));
  NA2        u0052(.A(i_5_), .B(i_9_), .Y(men_men_n75_));
  AOI210     u0053(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n72_), .Y(men_men_n77_));
  OAI210     u0055(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n77_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n78_), .A1(men_men_n68_), .B0(i_0_), .Y(men_men_n79_));
  NA2        u0057(.A(i_12_), .B(i_5_), .Y(men_men_n80_));
  NA2        u0058(.A(i_2_), .B(i_8_), .Y(men_men_n81_));
  NO2        u0059(.A(men_men_n81_), .B(men_men_n58_), .Y(men_men_n82_));
  NO2        u0060(.A(i_3_), .B(i_9_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_7_), .Y(men_men_n84_));
  NO3        u0062(.A(men_men_n84_), .B(men_men_n83_), .C(men_men_n63_), .Y(men_men_n85_));
  INV        u0063(.A(i_6_), .Y(men_men_n86_));
  OR4        u0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n87_));
  INV        u0065(.A(men_men_n87_), .Y(men_men_n88_));
  NO2        u0066(.A(i_2_), .B(i_7_), .Y(men_men_n89_));
  AOI210     u0067(.A0(men_men_n88_), .A1(men_men_n86_), .B0(men_men_n89_), .Y(men_men_n90_));
  OAI210     u0068(.A0(men_men_n85_), .A1(men_men_n82_), .B0(men_men_n90_), .Y(men_men_n91_));
  NAi21      u0069(.An(i_6_), .B(i_10_), .Y(men_men_n92_));
  NA2        u0070(.A(i_6_), .B(i_9_), .Y(men_men_n93_));
  AOI210     u0071(.A0(men_men_n93_), .A1(men_men_n92_), .B0(men_men_n63_), .Y(men_men_n94_));
  NA2        u0072(.A(i_2_), .B(i_6_), .Y(men_men_n95_));
  NO3        u0073(.A(men_men_n95_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n96_));
  NO2        u0074(.A(men_men_n96_), .B(men_men_n94_), .Y(men_men_n97_));
  AOI210     u0075(.A0(men_men_n97_), .A1(men_men_n91_), .B0(men_men_n80_), .Y(men_men_n98_));
  AN3        u0076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n99_));
  NAi21      u0077(.An(i_6_), .B(i_11_), .Y(men_men_n100_));
  NO2        u0078(.A(i_5_), .B(i_8_), .Y(men_men_n101_));
  NOi21      u0079(.An(men_men_n101_), .B(men_men_n100_), .Y(men_men_n102_));
  NA2        u0080(.A(men_men_n102_), .B(men_men_n62_), .Y(men_men_n103_));
  INV        u0081(.A(i_7_), .Y(men_men_n104_));
  NA2        u0082(.A(men_men_n46_), .B(men_men_n104_), .Y(men_men_n105_));
  NO2        u0083(.A(i_0_), .B(i_5_), .Y(men_men_n106_));
  NO2        u0084(.A(men_men_n106_), .B(men_men_n86_), .Y(men_men_n107_));
  NA2        u0085(.A(i_12_), .B(i_3_), .Y(men_men_n108_));
  NAi21      u0086(.An(i_7_), .B(i_11_), .Y(men_men_n109_));
  NO3        u0087(.A(men_men_n109_), .B(men_men_n92_), .C(men_men_n53_), .Y(men_men_n110_));
  AN2        u0088(.A(i_2_), .B(i_10_), .Y(men_men_n111_));
  OR2        u0089(.A(men_men_n80_), .B(men_men_n58_), .Y(men_men_n112_));
  NO2        u0090(.A(i_8_), .B(men_men_n104_), .Y(men_men_n113_));
  NA2        u0091(.A(i_12_), .B(i_7_), .Y(men_men_n114_));
  NO2        u0092(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n115_));
  NA2        u0093(.A(men_men_n115_), .B(i_0_), .Y(men_men_n116_));
  NA2        u0094(.A(i_11_), .B(i_12_), .Y(men_men_n117_));
  OAI210     u0095(.A0(men_men_n116_), .A1(men_men_n114_), .B0(men_men_n117_), .Y(men_men_n118_));
  INV        u0096(.A(men_men_n118_), .Y(men_men_n119_));
  NAi31      u0097(.An(men_men_n110_), .B(men_men_n119_), .C(men_men_n103_), .Y(men_men_n120_));
  NOi21      u0098(.An(i_1_), .B(i_5_), .Y(men_men_n121_));
  NA2        u0099(.A(men_men_n121_), .B(i_11_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n104_), .B(men_men_n37_), .Y(men_men_n123_));
  NA2        u0101(.A(i_7_), .B(men_men_n25_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NO2        u0103(.A(men_men_n125_), .B(men_men_n46_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n127_));
  NAi21      u0105(.An(i_3_), .B(i_8_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n128_), .B(men_men_n62_), .Y(men_men_n129_));
  NO2        u0107(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n130_));
  NO2        u0108(.A(i_1_), .B(men_men_n86_), .Y(men_men_n131_));
  NO2        u0109(.A(i_6_), .B(i_5_), .Y(men_men_n132_));
  NA2        u0110(.A(men_men_n132_), .B(i_3_), .Y(men_men_n133_));
  AO210      u0111(.A0(men_men_n133_), .A1(men_men_n47_), .B0(men_men_n131_), .Y(men_men_n134_));
  OAI220     u0112(.A0(men_men_n134_), .A1(men_men_n109_), .B0(men_men_n130_), .B1(men_men_n122_), .Y(men_men_n135_));
  NO3        u0113(.A(men_men_n135_), .B(men_men_n120_), .C(men_men_n98_), .Y(men_men_n136_));
  NA3        u0114(.A(men_men_n136_), .B(men_men_n79_), .C(men_men_n56_), .Y(men2));
  NO2        u0115(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n138_));
  NA2        u0116(.A(i_6_), .B(men_men_n25_), .Y(men_men_n139_));
  NA2        u0117(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  NA4        u0118(.A(men_men_n140_), .B(men_men_n77_), .C(men_men_n69_), .D(men_men_n30_), .Y(men0));
  AN2        u0119(.A(i_8_), .B(i_7_), .Y(men_men_n142_));
  NA2        u0120(.A(men_men_n142_), .B(i_6_), .Y(men_men_n143_));
  NO2        u0121(.A(i_12_), .B(i_13_), .Y(men_men_n144_));
  NAi21      u0122(.An(i_5_), .B(i_11_), .Y(men_men_n145_));
  NOi21      u0123(.An(men_men_n144_), .B(men_men_n145_), .Y(men_men_n146_));
  NO2        u0124(.A(i_0_), .B(i_1_), .Y(men_men_n147_));
  NA2        u0125(.A(i_2_), .B(i_3_), .Y(men_men_n148_));
  NO2        u0126(.A(men_men_n148_), .B(i_4_), .Y(men_men_n149_));
  NA3        u0127(.A(men_men_n149_), .B(men_men_n147_), .C(men_men_n146_), .Y(men_men_n150_));
  OR2        u0128(.A(men_men_n150_), .B(men_men_n25_), .Y(men_men_n151_));
  AN2        u0129(.A(men_men_n144_), .B(men_men_n83_), .Y(men_men_n152_));
  NO2        u0130(.A(men_men_n152_), .B(men_men_n27_), .Y(men_men_n153_));
  NA2        u0131(.A(i_1_), .B(i_5_), .Y(men_men_n154_));
  NO2        u0132(.A(men_men_n73_), .B(men_men_n46_), .Y(men_men_n155_));
  NA2        u0133(.A(men_men_n155_), .B(men_men_n36_), .Y(men_men_n156_));
  NO3        u0134(.A(men_men_n156_), .B(men_men_n154_), .C(men_men_n153_), .Y(men_men_n157_));
  OR2        u0135(.A(i_0_), .B(i_1_), .Y(men_men_n158_));
  NO3        u0136(.A(men_men_n158_), .B(men_men_n80_), .C(i_13_), .Y(men_men_n159_));
  NAi32      u0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n160_));
  NAi21      u0138(.An(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  NOi21      u0139(.An(i_4_), .B(i_10_), .Y(men_men_n162_));
  NA2        u0140(.A(men_men_n162_), .B(men_men_n39_), .Y(men_men_n163_));
  NO2        u0141(.A(i_3_), .B(i_5_), .Y(men_men_n164_));
  NO3        u0142(.A(men_men_n73_), .B(i_2_), .C(i_1_), .Y(men_men_n165_));
  NA2        u0143(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  OAI210     u0144(.A0(men_men_n166_), .A1(men_men_n163_), .B0(men_men_n161_), .Y(men_men_n167_));
  NO2        u0145(.A(men_men_n167_), .B(men_men_n157_), .Y(men_men_n168_));
  AOI210     u0146(.A0(men_men_n168_), .A1(men_men_n151_), .B0(men_men_n143_), .Y(men_men_n169_));
  NA3        u0147(.A(men_men_n73_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n170_));
  NA2        u0148(.A(i_3_), .B(men_men_n48_), .Y(men_men_n171_));
  NOi21      u0149(.An(i_4_), .B(i_9_), .Y(men_men_n172_));
  NOi21      u0150(.An(i_11_), .B(i_13_), .Y(men_men_n173_));
  NA2        u0151(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  OR2        u0152(.A(men_men_n174_), .B(men_men_n171_), .Y(men_men_n175_));
  NO2        u0153(.A(i_4_), .B(i_5_), .Y(men_men_n176_));
  NAi21      u0154(.An(i_12_), .B(i_11_), .Y(men_men_n177_));
  NO2        u0155(.A(men_men_n177_), .B(i_13_), .Y(men_men_n178_));
  NA3        u0156(.A(men_men_n178_), .B(men_men_n176_), .C(men_men_n83_), .Y(men_men_n179_));
  AOI210     u0157(.A0(men_men_n179_), .A1(men_men_n175_), .B0(men_men_n170_), .Y(men_men_n180_));
  NO2        u0158(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n181_));
  NA2        u0159(.A(men_men_n181_), .B(men_men_n46_), .Y(men_men_n182_));
  NA2        u0160(.A(men_men_n36_), .B(i_5_), .Y(men_men_n183_));
  NAi31      u0161(.An(men_men_n183_), .B(men_men_n152_), .C(i_11_), .Y(men_men_n184_));
  NA2        u0162(.A(i_3_), .B(i_5_), .Y(men_men_n185_));
  OR2        u0163(.A(men_men_n185_), .B(men_men_n174_), .Y(men_men_n186_));
  AOI210     u0164(.A0(men_men_n186_), .A1(men_men_n184_), .B0(men_men_n182_), .Y(men_men_n187_));
  NO2        u0165(.A(men_men_n73_), .B(i_5_), .Y(men_men_n188_));
  NO2        u0166(.A(i_13_), .B(i_10_), .Y(men_men_n189_));
  NA3        u0167(.A(men_men_n189_), .B(men_men_n188_), .C(men_men_n44_), .Y(men_men_n190_));
  NO2        u0168(.A(i_2_), .B(i_1_), .Y(men_men_n191_));
  NAi21      u0169(.An(i_4_), .B(i_12_), .Y(men_men_n192_));
  NO4        u0170(.A(men_men_n192_), .B(i_1_), .C(men_men_n190_), .D(men_men_n25_), .Y(men_men_n193_));
  NO3        u0171(.A(men_men_n193_), .B(men_men_n187_), .C(men_men_n180_), .Y(men_men_n194_));
  INV        u0172(.A(i_8_), .Y(men_men_n195_));
  NO2        u0173(.A(men_men_n195_), .B(i_7_), .Y(men_men_n196_));
  NA2        u0174(.A(men_men_n196_), .B(i_6_), .Y(men_men_n197_));
  NO3        u0175(.A(i_3_), .B(men_men_n86_), .C(men_men_n48_), .Y(men_men_n198_));
  NA2        u0176(.A(men_men_n198_), .B(men_men_n113_), .Y(men_men_n199_));
  NO3        u0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n200_));
  NA3        u0178(.A(men_men_n200_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n201_));
  NO3        u0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n202_));
  OAI210     u0180(.A0(men_men_n99_), .A1(i_12_), .B0(men_men_n202_), .Y(men_men_n203_));
  AOI210     u0181(.A0(men_men_n203_), .A1(men_men_n201_), .B0(men_men_n199_), .Y(men_men_n204_));
  NO2        u0182(.A(i_3_), .B(i_8_), .Y(men_men_n205_));
  NO3        u0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n206_));
  NA3        u0184(.A(men_men_n206_), .B(men_men_n205_), .C(men_men_n39_), .Y(men_men_n207_));
  NO2        u0185(.A(men_men_n106_), .B(men_men_n58_), .Y(men_men_n208_));
  INV        u0186(.A(men_men_n208_), .Y(men_men_n209_));
  NO2        u0187(.A(i_13_), .B(i_9_), .Y(men_men_n210_));
  NA3        u0188(.A(men_men_n210_), .B(i_6_), .C(men_men_n195_), .Y(men_men_n211_));
  NAi21      u0189(.An(i_12_), .B(i_3_), .Y(men_men_n212_));
  NO2        u0190(.A(men_men_n44_), .B(i_5_), .Y(men_men_n213_));
  NO3        u0191(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n214_));
  NA3        u0192(.A(men_men_n214_), .B(men_men_n213_), .C(i_10_), .Y(men_men_n215_));
  OAI220     u0193(.A0(men_men_n215_), .A1(men_men_n211_), .B0(men_men_n209_), .B1(men_men_n207_), .Y(men_men_n216_));
  AOI210     u0194(.A0(men_men_n216_), .A1(i_7_), .B0(men_men_n204_), .Y(men_men_n217_));
  OAI220     u0195(.A0(men_men_n217_), .A1(i_4_), .B0(men_men_n197_), .B1(men_men_n194_), .Y(men_men_n218_));
  NAi21      u0196(.An(i_12_), .B(i_7_), .Y(men_men_n219_));
  NA3        u0197(.A(i_13_), .B(men_men_n195_), .C(i_10_), .Y(men_men_n220_));
  NO2        u0198(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n221_));
  NA2        u0199(.A(i_0_), .B(i_5_), .Y(men_men_n222_));
  NA2        u0200(.A(men_men_n222_), .B(men_men_n107_), .Y(men_men_n223_));
  OAI220     u0201(.A0(men_men_n223_), .A1(i_1_), .B0(men_men_n182_), .B1(men_men_n133_), .Y(men_men_n224_));
  NAi31      u0202(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n225_));
  NO2        u0203(.A(men_men_n36_), .B(i_13_), .Y(men_men_n226_));
  NO2        u0204(.A(men_men_n73_), .B(men_men_n26_), .Y(men_men_n227_));
  NO2        u0205(.A(men_men_n46_), .B(men_men_n63_), .Y(men_men_n228_));
  NA3        u0206(.A(men_men_n228_), .B(men_men_n227_), .C(men_men_n226_), .Y(men_men_n229_));
  INV        u0207(.A(i_13_), .Y(men_men_n230_));
  NO2        u0208(.A(i_12_), .B(men_men_n230_), .Y(men_men_n231_));
  NA3        u0209(.A(men_men_n231_), .B(men_men_n200_), .C(men_men_n198_), .Y(men_men_n232_));
  OAI210     u0210(.A0(men_men_n229_), .A1(men_men_n225_), .B0(men_men_n232_), .Y(men_men_n233_));
  AOI220     u0211(.A0(men_men_n233_), .A1(men_men_n142_), .B0(men_men_n224_), .B1(men_men_n221_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n185_), .B(i_4_), .Y(men_men_n235_));
  INV        u0213(.A(men_men_n235_), .Y(men_men_n236_));
  OR2        u0214(.A(i_8_), .B(i_7_), .Y(men_men_n237_));
  NO2        u0215(.A(men_men_n237_), .B(men_men_n86_), .Y(men_men_n238_));
  NO2        u0216(.A(men_men_n53_), .B(i_1_), .Y(men_men_n239_));
  NA2        u0217(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n240_));
  INV        u0218(.A(i_12_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n44_), .B(men_men_n241_), .Y(men_men_n242_));
  NO3        u0220(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n243_));
  NA2        u0221(.A(i_2_), .B(i_1_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n240_), .B(men_men_n236_), .Y(men_men_n245_));
  NO3        u0223(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n246_));
  NAi21      u0224(.An(i_4_), .B(i_3_), .Y(men_men_n247_));
  NO2        u0225(.A(men_men_n247_), .B(men_men_n75_), .Y(men_men_n248_));
  NO2        u0226(.A(i_0_), .B(i_6_), .Y(men_men_n249_));
  NOi41      u0227(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n250_));
  NA2        u0228(.A(men_men_n250_), .B(men_men_n249_), .Y(men_men_n251_));
  NO2        u0229(.A(men_men_n244_), .B(men_men_n185_), .Y(men_men_n252_));
  NAi21      u0230(.An(men_men_n251_), .B(men_men_n252_), .Y(men_men_n253_));
  INV        u0231(.A(men_men_n253_), .Y(men_men_n254_));
  AOI220     u0232(.A0(men_men_n254_), .A1(men_men_n39_), .B0(men_men_n245_), .B1(men_men_n210_), .Y(men_men_n255_));
  NO2        u0233(.A(i_11_), .B(men_men_n230_), .Y(men_men_n256_));
  NOi21      u0234(.An(i_1_), .B(i_6_), .Y(men_men_n257_));
  NAi21      u0235(.An(i_3_), .B(i_7_), .Y(men_men_n258_));
  NA2        u0236(.A(men_men_n241_), .B(i_9_), .Y(men_men_n259_));
  OR4        u0237(.A(men_men_n259_), .B(men_men_n258_), .C(men_men_n257_), .D(men_men_n188_), .Y(men_men_n260_));
  NO2        u0238(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n261_));
  NO2        u0239(.A(i_12_), .B(i_3_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n73_), .B(i_5_), .Y(men_men_n263_));
  NA2        u0241(.A(i_3_), .B(i_9_), .Y(men_men_n264_));
  NAi21      u0242(.An(i_7_), .B(i_10_), .Y(men_men_n265_));
  NO2        u0243(.A(men_men_n265_), .B(men_men_n264_), .Y(men_men_n266_));
  NA3        u0244(.A(men_men_n266_), .B(men_men_n263_), .C(men_men_n64_), .Y(men_men_n267_));
  NA2        u0245(.A(men_men_n267_), .B(men_men_n260_), .Y(men_men_n268_));
  NA3        u0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n269_));
  INV        u0247(.A(men_men_n143_), .Y(men_men_n270_));
  NA2        u0248(.A(men_men_n241_), .B(i_13_), .Y(men_men_n271_));
  NO2        u0249(.A(men_men_n271_), .B(men_men_n75_), .Y(men_men_n272_));
  AOI220     u0250(.A0(men_men_n272_), .A1(men_men_n270_), .B0(men_men_n268_), .B1(men_men_n256_), .Y(men_men_n273_));
  NO2        u0251(.A(men_men_n237_), .B(men_men_n37_), .Y(men_men_n274_));
  NA2        u0252(.A(i_12_), .B(i_6_), .Y(men_men_n275_));
  OR2        u0253(.A(i_13_), .B(i_9_), .Y(men_men_n276_));
  NO3        u0254(.A(men_men_n276_), .B(men_men_n275_), .C(men_men_n48_), .Y(men_men_n277_));
  NO2        u0255(.A(men_men_n247_), .B(i_2_), .Y(men_men_n278_));
  NA3        u0256(.A(men_men_n278_), .B(men_men_n277_), .C(men_men_n44_), .Y(men_men_n279_));
  NA2        u0257(.A(men_men_n256_), .B(i_9_), .Y(men_men_n280_));
  NA2        u0258(.A(men_men_n263_), .B(men_men_n64_), .Y(men_men_n281_));
  OAI210     u0259(.A0(men_men_n281_), .A1(men_men_n280_), .B0(men_men_n279_), .Y(men_men_n282_));
  NO3        u0260(.A(i_11_), .B(men_men_n230_), .C(men_men_n25_), .Y(men_men_n283_));
  NO2        u0261(.A(men_men_n258_), .B(i_8_), .Y(men_men_n284_));
  NO2        u0262(.A(i_6_), .B(men_men_n48_), .Y(men_men_n285_));
  NA3        u0263(.A(men_men_n285_), .B(men_men_n284_), .C(men_men_n283_), .Y(men_men_n286_));
  NO3        u0264(.A(men_men_n26_), .B(men_men_n86_), .C(i_5_), .Y(men_men_n287_));
  NA3        u0265(.A(men_men_n287_), .B(men_men_n274_), .C(men_men_n231_), .Y(men_men_n288_));
  AOI210     u0266(.A0(men_men_n288_), .A1(men_men_n286_), .B0(i_1_), .Y(men_men_n289_));
  AOI210     u0267(.A0(men_men_n282_), .A1(men_men_n274_), .B0(men_men_n289_), .Y(men_men_n290_));
  NA4        u0268(.A(men_men_n290_), .B(men_men_n273_), .C(men_men_n255_), .D(men_men_n234_), .Y(men_men_n291_));
  NO3        u0269(.A(i_12_), .B(men_men_n230_), .C(men_men_n37_), .Y(men_men_n292_));
  INV        u0270(.A(men_men_n292_), .Y(men_men_n293_));
  NOi21      u0271(.An(men_men_n164_), .B(men_men_n86_), .Y(men_men_n294_));
  NO3        u0272(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n295_));
  AOI220     u0273(.A0(men_men_n295_), .A1(men_men_n198_), .B0(men_men_n294_), .B1(men_men_n239_), .Y(men_men_n296_));
  NO2        u0274(.A(men_men_n296_), .B(i_7_), .Y(men_men_n297_));
  NO3        u0275(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n298_));
  NO2        u0276(.A(men_men_n244_), .B(i_0_), .Y(men_men_n299_));
  AOI220     u0277(.A0(men_men_n299_), .A1(men_men_n196_), .B0(men_men_n298_), .B1(men_men_n142_), .Y(men_men_n300_));
  NA2        u0278(.A(men_men_n285_), .B(men_men_n26_), .Y(men_men_n301_));
  NO2        u0279(.A(men_men_n301_), .B(men_men_n300_), .Y(men_men_n302_));
  NA2        u0280(.A(i_0_), .B(i_1_), .Y(men_men_n303_));
  NO2        u0281(.A(men_men_n303_), .B(i_2_), .Y(men_men_n304_));
  NO2        u0282(.A(men_men_n59_), .B(i_6_), .Y(men_men_n305_));
  NA3        u0283(.A(men_men_n305_), .B(men_men_n304_), .C(men_men_n164_), .Y(men_men_n306_));
  OAI210     u0284(.A0(men_men_n166_), .A1(men_men_n143_), .B0(men_men_n306_), .Y(men_men_n307_));
  NO3        u0285(.A(men_men_n307_), .B(men_men_n302_), .C(men_men_n297_), .Y(men_men_n308_));
  NO2        u0286(.A(i_3_), .B(i_10_), .Y(men_men_n309_));
  NA3        u0287(.A(men_men_n309_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n310_));
  NO2        u0288(.A(i_2_), .B(men_men_n104_), .Y(men_men_n311_));
  NA2        u0289(.A(i_1_), .B(men_men_n36_), .Y(men_men_n312_));
  NOi21      u0290(.An(men_men_n222_), .B(men_men_n106_), .Y(men_men_n313_));
  NA3        u0291(.A(men_men_n313_), .B(i_1_), .C(men_men_n311_), .Y(men_men_n314_));
  AN2        u0292(.A(i_3_), .B(i_10_), .Y(men_men_n315_));
  NA4        u0293(.A(men_men_n315_), .B(men_men_n200_), .C(men_men_n178_), .D(men_men_n176_), .Y(men_men_n316_));
  NO2        u0294(.A(i_5_), .B(men_men_n37_), .Y(men_men_n317_));
  NO2        u0295(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n318_));
  OR2        u0296(.A(men_men_n314_), .B(men_men_n310_), .Y(men_men_n319_));
  OAI220     u0297(.A0(men_men_n319_), .A1(i_6_), .B0(men_men_n308_), .B1(men_men_n293_), .Y(men_men_n320_));
  NO4        u0298(.A(men_men_n320_), .B(men_men_n291_), .C(men_men_n218_), .D(men_men_n169_), .Y(men_men_n321_));
  NO3        u0299(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n322_));
  NO2        u0300(.A(men_men_n59_), .B(men_men_n86_), .Y(men_men_n323_));
  NA2        u0301(.A(men_men_n299_), .B(men_men_n323_), .Y(men_men_n324_));
  NO3        u0302(.A(i_6_), .B(men_men_n195_), .C(i_7_), .Y(men_men_n325_));
  NA2        u0303(.A(men_men_n325_), .B(men_men_n200_), .Y(men_men_n326_));
  AOI210     u0304(.A0(men_men_n326_), .A1(men_men_n324_), .B0(men_men_n171_), .Y(men_men_n327_));
  NO2        u0305(.A(i_2_), .B(i_3_), .Y(men_men_n328_));
  OR2        u0306(.A(i_0_), .B(i_5_), .Y(men_men_n329_));
  NA2        u0307(.A(men_men_n222_), .B(men_men_n329_), .Y(men_men_n330_));
  NA4        u0308(.A(men_men_n330_), .B(men_men_n238_), .C(men_men_n328_), .D(i_1_), .Y(men_men_n331_));
  NA3        u0309(.A(men_men_n299_), .B(men_men_n294_), .C(men_men_n113_), .Y(men_men_n332_));
  NAi21      u0310(.An(i_8_), .B(i_7_), .Y(men_men_n333_));
  NO2        u0311(.A(men_men_n333_), .B(i_6_), .Y(men_men_n334_));
  NO2        u0312(.A(men_men_n158_), .B(men_men_n46_), .Y(men_men_n335_));
  NA3        u0313(.A(men_men_n335_), .B(men_men_n334_), .C(men_men_n164_), .Y(men_men_n336_));
  NA3        u0314(.A(men_men_n336_), .B(men_men_n332_), .C(men_men_n331_), .Y(men_men_n337_));
  OAI210     u0315(.A0(men_men_n337_), .A1(men_men_n327_), .B0(i_4_), .Y(men_men_n338_));
  NO2        u0316(.A(i_12_), .B(i_10_), .Y(men_men_n339_));
  NOi21      u0317(.An(i_5_), .B(i_0_), .Y(men_men_n340_));
  AOI210     u0318(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n104_), .Y(men_men_n341_));
  NO4        u0319(.A(men_men_n341_), .B(men_men_n312_), .C(men_men_n340_), .D(men_men_n128_), .Y(men_men_n342_));
  NA4        u0320(.A(men_men_n84_), .B(men_men_n36_), .C(men_men_n86_), .D(i_8_), .Y(men_men_n343_));
  NA2        u0321(.A(men_men_n342_), .B(men_men_n339_), .Y(men_men_n344_));
  NO2        u0322(.A(i_6_), .B(i_8_), .Y(men_men_n345_));
  NOi21      u0323(.An(i_0_), .B(i_2_), .Y(men_men_n346_));
  AN2        u0324(.A(men_men_n346_), .B(men_men_n345_), .Y(men_men_n347_));
  NO2        u0325(.A(i_1_), .B(i_7_), .Y(men_men_n348_));
  AO220      u0326(.A0(men_men_n348_), .A1(men_men_n347_), .B0(men_men_n334_), .B1(men_men_n239_), .Y(men_men_n349_));
  NA3        u0327(.A(men_men_n349_), .B(men_men_n41_), .C(i_5_), .Y(men_men_n350_));
  NA3        u0328(.A(men_men_n350_), .B(men_men_n344_), .C(men_men_n338_), .Y(men_men_n351_));
  NO3        u0329(.A(men_men_n237_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n352_));
  NO3        u0330(.A(men_men_n333_), .B(i_2_), .C(i_1_), .Y(men_men_n353_));
  OAI210     u0331(.A0(men_men_n353_), .A1(men_men_n352_), .B0(i_6_), .Y(men_men_n354_));
  NA3        u0332(.A(men_men_n257_), .B(men_men_n311_), .C(men_men_n195_), .Y(men_men_n355_));
  AOI210     u0333(.A0(men_men_n355_), .A1(men_men_n354_), .B0(men_men_n330_), .Y(men_men_n356_));
  NOi21      u0334(.An(men_men_n154_), .B(men_men_n107_), .Y(men_men_n357_));
  NO2        u0335(.A(men_men_n357_), .B(men_men_n124_), .Y(men_men_n358_));
  OAI210     u0336(.A0(men_men_n358_), .A1(men_men_n356_), .B0(i_3_), .Y(men_men_n359_));
  INV        u0337(.A(men_men_n84_), .Y(men_men_n360_));
  NO2        u0338(.A(men_men_n303_), .B(men_men_n81_), .Y(men_men_n361_));
  NA2        u0339(.A(men_men_n361_), .B(men_men_n132_), .Y(men_men_n362_));
  NO2        u0340(.A(men_men_n95_), .B(men_men_n195_), .Y(men_men_n363_));
  NA3        u0341(.A(men_men_n313_), .B(men_men_n363_), .C(men_men_n63_), .Y(men_men_n364_));
  AOI210     u0342(.A0(men_men_n364_), .A1(men_men_n362_), .B0(men_men_n360_), .Y(men_men_n365_));
  NO2        u0343(.A(men_men_n195_), .B(i_9_), .Y(men_men_n366_));
  NA2        u0344(.A(men_men_n366_), .B(men_men_n208_), .Y(men_men_n367_));
  NO2        u0345(.A(men_men_n367_), .B(men_men_n46_), .Y(men_men_n368_));
  NO3        u0346(.A(men_men_n368_), .B(men_men_n365_), .C(men_men_n302_), .Y(men_men_n369_));
  AOI210     u0347(.A0(men_men_n369_), .A1(men_men_n359_), .B0(men_men_n163_), .Y(men_men_n370_));
  AOI210     u0348(.A0(men_men_n351_), .A1(men_men_n322_), .B0(men_men_n370_), .Y(men_men_n371_));
  NOi32      u0349(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n372_));
  INV        u0350(.A(men_men_n372_), .Y(men_men_n373_));
  NAi21      u0351(.An(i_0_), .B(i_6_), .Y(men_men_n374_));
  NAi21      u0352(.An(i_1_), .B(i_5_), .Y(men_men_n375_));
  NA2        u0353(.A(men_men_n375_), .B(men_men_n374_), .Y(men_men_n376_));
  NA2        u0354(.A(men_men_n376_), .B(men_men_n25_), .Y(men_men_n377_));
  OAI210     u0355(.A0(men_men_n377_), .A1(men_men_n160_), .B0(men_men_n251_), .Y(men_men_n378_));
  NAi41      u0356(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n379_));
  OAI220     u0357(.A0(men_men_n379_), .A1(men_men_n375_), .B0(men_men_n225_), .B1(men_men_n160_), .Y(men_men_n380_));
  AOI210     u0358(.A0(men_men_n379_), .A1(men_men_n160_), .B0(men_men_n158_), .Y(men_men_n381_));
  NOi32      u0359(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n382_));
  NAi21      u0360(.An(i_6_), .B(i_1_), .Y(men_men_n383_));
  NA3        u0361(.A(men_men_n383_), .B(men_men_n382_), .C(men_men_n46_), .Y(men_men_n384_));
  NO2        u0362(.A(men_men_n384_), .B(i_0_), .Y(men_men_n385_));
  OR3        u0363(.A(men_men_n385_), .B(men_men_n381_), .C(men_men_n380_), .Y(men_men_n386_));
  NO2        u0364(.A(i_1_), .B(men_men_n104_), .Y(men_men_n387_));
  NAi21      u0365(.An(i_3_), .B(i_4_), .Y(men_men_n388_));
  NO2        u0366(.A(men_men_n388_), .B(i_9_), .Y(men_men_n389_));
  AN2        u0367(.A(i_6_), .B(i_7_), .Y(men_men_n390_));
  OAI210     u0368(.A0(men_men_n390_), .A1(men_men_n387_), .B0(men_men_n389_), .Y(men_men_n391_));
  NA2        u0369(.A(i_2_), .B(i_7_), .Y(men_men_n392_));
  NO2        u0370(.A(men_men_n388_), .B(i_10_), .Y(men_men_n393_));
  NA3        u0371(.A(men_men_n393_), .B(men_men_n392_), .C(men_men_n249_), .Y(men_men_n394_));
  AOI210     u0372(.A0(men_men_n394_), .A1(men_men_n391_), .B0(men_men_n188_), .Y(men_men_n395_));
  AOI210     u0373(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n396_));
  OAI210     u0374(.A0(men_men_n396_), .A1(men_men_n191_), .B0(men_men_n393_), .Y(men_men_n397_));
  AOI220     u0375(.A0(men_men_n393_), .A1(men_men_n348_), .B0(men_men_n243_), .B1(men_men_n191_), .Y(men_men_n398_));
  AOI210     u0376(.A0(men_men_n398_), .A1(men_men_n397_), .B0(i_5_), .Y(men_men_n399_));
  NO4        u0377(.A(men_men_n399_), .B(men_men_n395_), .C(men_men_n386_), .D(men_men_n378_), .Y(men_men_n400_));
  NO2        u0378(.A(men_men_n400_), .B(men_men_n373_), .Y(men_men_n401_));
  NO2        u0379(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n402_));
  AN2        u0380(.A(i_12_), .B(i_5_), .Y(men_men_n403_));
  NO2        u0381(.A(i_4_), .B(men_men_n26_), .Y(men_men_n404_));
  NA2        u0382(.A(men_men_n404_), .B(men_men_n403_), .Y(men_men_n405_));
  NO2        u0383(.A(i_11_), .B(i_6_), .Y(men_men_n406_));
  NA3        u0384(.A(men_men_n406_), .B(men_men_n335_), .C(men_men_n230_), .Y(men_men_n407_));
  NO2        u0385(.A(men_men_n407_), .B(men_men_n405_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n247_), .B(i_5_), .Y(men_men_n409_));
  NO2        u0387(.A(i_5_), .B(i_10_), .Y(men_men_n410_));
  AOI220     u0388(.A0(men_men_n410_), .A1(men_men_n278_), .B0(men_men_n409_), .B1(men_men_n200_), .Y(men_men_n411_));
  NA2        u0389(.A(men_men_n144_), .B(men_men_n45_), .Y(men_men_n412_));
  NO2        u0390(.A(men_men_n412_), .B(men_men_n411_), .Y(men_men_n413_));
  OAI210     u0391(.A0(men_men_n413_), .A1(men_men_n408_), .B0(men_men_n402_), .Y(men_men_n414_));
  NO2        u0392(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n415_));
  NO2        u0393(.A(men_men_n150_), .B(men_men_n86_), .Y(men_men_n416_));
  OAI210     u0394(.A0(men_men_n416_), .A1(men_men_n408_), .B0(men_men_n415_), .Y(men_men_n417_));
  NO3        u0395(.A(men_men_n86_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n418_));
  NO2        u0396(.A(i_3_), .B(men_men_n104_), .Y(men_men_n419_));
  NA2        u0397(.A(men_men_n309_), .B(men_men_n75_), .Y(men_men_n420_));
  NO2        u0398(.A(i_11_), .B(i_12_), .Y(men_men_n421_));
  NA2        u0399(.A(men_men_n421_), .B(men_men_n36_), .Y(men_men_n422_));
  NO2        u0400(.A(men_men_n420_), .B(men_men_n422_), .Y(men_men_n423_));
  NA2        u0401(.A(men_men_n410_), .B(men_men_n241_), .Y(men_men_n424_));
  NA3        u0402(.A(men_men_n113_), .B(men_men_n41_), .C(i_11_), .Y(men_men_n425_));
  NO2        u0403(.A(men_men_n425_), .B(men_men_n225_), .Y(men_men_n426_));
  NAi21      u0404(.An(i_13_), .B(i_0_), .Y(men_men_n427_));
  NO2        u0405(.A(men_men_n427_), .B(men_men_n244_), .Y(men_men_n428_));
  OAI210     u0406(.A0(men_men_n426_), .A1(men_men_n423_), .B0(men_men_n428_), .Y(men_men_n429_));
  NA3        u0407(.A(men_men_n429_), .B(men_men_n417_), .C(men_men_n414_), .Y(men_men_n430_));
  NA2        u0408(.A(men_men_n44_), .B(men_men_n230_), .Y(men_men_n431_));
  NO3        u0409(.A(i_1_), .B(i_12_), .C(men_men_n86_), .Y(men_men_n432_));
  NO2        u0410(.A(i_0_), .B(i_11_), .Y(men_men_n433_));
  AN2        u0411(.A(i_1_), .B(i_6_), .Y(men_men_n434_));
  NOi21      u0412(.An(i_2_), .B(i_12_), .Y(men_men_n435_));
  NA2        u0413(.A(men_men_n435_), .B(men_men_n434_), .Y(men_men_n436_));
  NO2        u0414(.A(men_men_n436_), .B(men_men_n1109_), .Y(men_men_n437_));
  NO2        u0415(.A(men_men_n1113_), .B(i_4_), .Y(men_men_n438_));
  NA2        u0416(.A(men_men_n437_), .B(men_men_n438_), .Y(men_men_n439_));
  NAi21      u0417(.An(i_9_), .B(i_4_), .Y(men_men_n440_));
  OR2        u0418(.A(i_13_), .B(i_10_), .Y(men_men_n441_));
  NO3        u0419(.A(men_men_n441_), .B(men_men_n117_), .C(men_men_n440_), .Y(men_men_n442_));
  NO2        u0420(.A(men_men_n174_), .B(men_men_n123_), .Y(men_men_n443_));
  OR2        u0421(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n444_));
  NO2        u0422(.A(men_men_n104_), .B(men_men_n25_), .Y(men_men_n445_));
  NA2        u0423(.A(men_men_n292_), .B(men_men_n445_), .Y(men_men_n446_));
  NA2        u0424(.A(men_men_n285_), .B(men_men_n214_), .Y(men_men_n447_));
  OAI220     u0425(.A0(men_men_n447_), .A1(men_men_n444_), .B0(men_men_n446_), .B1(men_men_n357_), .Y(men_men_n448_));
  INV        u0426(.A(men_men_n448_), .Y(men_men_n449_));
  AOI210     u0427(.A0(men_men_n449_), .A1(men_men_n439_), .B0(men_men_n26_), .Y(men_men_n450_));
  NA2        u0428(.A(men_men_n332_), .B(men_men_n331_), .Y(men_men_n451_));
  AOI220     u0429(.A0(men_men_n305_), .A1(men_men_n295_), .B0(men_men_n299_), .B1(men_men_n323_), .Y(men_men_n452_));
  NO2        u0430(.A(men_men_n452_), .B(men_men_n171_), .Y(men_men_n453_));
  NO2        u0431(.A(men_men_n185_), .B(men_men_n86_), .Y(men_men_n454_));
  AOI220     u0432(.A0(men_men_n454_), .A1(men_men_n304_), .B0(men_men_n287_), .B1(men_men_n214_), .Y(men_men_n455_));
  NO2        u0433(.A(men_men_n455_), .B(i_7_), .Y(men_men_n456_));
  NO3        u0434(.A(men_men_n456_), .B(men_men_n453_), .C(men_men_n451_), .Y(men_men_n457_));
  NA2        u0435(.A(men_men_n198_), .B(men_men_n99_), .Y(men_men_n458_));
  NA3        u0436(.A(men_men_n335_), .B(men_men_n164_), .C(men_men_n86_), .Y(men_men_n459_));
  AOI210     u0437(.A0(men_men_n459_), .A1(men_men_n458_), .B0(men_men_n333_), .Y(men_men_n460_));
  NA2        u0438(.A(men_men_n195_), .B(i_10_), .Y(men_men_n461_));
  NA3        u0439(.A(men_men_n263_), .B(men_men_n64_), .C(i_2_), .Y(men_men_n462_));
  NA2        u0440(.A(men_men_n305_), .B(men_men_n239_), .Y(men_men_n463_));
  OAI220     u0441(.A0(men_men_n463_), .A1(men_men_n185_), .B0(men_men_n462_), .B1(men_men_n461_), .Y(men_men_n464_));
  NO2        u0442(.A(i_3_), .B(men_men_n48_), .Y(men_men_n465_));
  NA3        u0443(.A(men_men_n348_), .B(men_men_n347_), .C(men_men_n465_), .Y(men_men_n466_));
  NA2        u0444(.A(men_men_n325_), .B(men_men_n330_), .Y(men_men_n467_));
  OAI210     u0445(.A0(men_men_n467_), .A1(i_1_), .B0(men_men_n466_), .Y(men_men_n468_));
  NO3        u0446(.A(men_men_n468_), .B(men_men_n464_), .C(men_men_n460_), .Y(men_men_n469_));
  AOI210     u0447(.A0(men_men_n469_), .A1(men_men_n457_), .B0(men_men_n280_), .Y(men_men_n470_));
  NO4        u0448(.A(men_men_n470_), .B(men_men_n450_), .C(men_men_n430_), .D(men_men_n401_), .Y(men_men_n471_));
  NO2        u0449(.A(men_men_n63_), .B(i_4_), .Y(men_men_n472_));
  NO2        u0450(.A(men_men_n73_), .B(i_13_), .Y(men_men_n473_));
  NO2        u0451(.A(i_10_), .B(i_9_), .Y(men_men_n474_));
  NAi21      u0452(.An(i_12_), .B(i_8_), .Y(men_men_n475_));
  NO2        u0453(.A(men_men_n475_), .B(i_3_), .Y(men_men_n476_));
  NO2        u0454(.A(men_men_n46_), .B(i_4_), .Y(men_men_n477_));
  NA2        u0455(.A(men_men_n477_), .B(men_men_n107_), .Y(men_men_n478_));
  NO2        u0456(.A(men_men_n478_), .B(men_men_n207_), .Y(men_men_n479_));
  NA2        u0457(.A(men_men_n318_), .B(i_0_), .Y(men_men_n480_));
  NO3        u0458(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n481_));
  NA2        u0459(.A(men_men_n275_), .B(men_men_n100_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n482_), .B(men_men_n481_), .Y(men_men_n483_));
  NA2        u0461(.A(i_8_), .B(i_9_), .Y(men_men_n484_));
  AOI210     u0462(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n485_));
  OR2        u0463(.A(men_men_n485_), .B(men_men_n484_), .Y(men_men_n486_));
  NA2        u0464(.A(men_men_n292_), .B(men_men_n208_), .Y(men_men_n487_));
  OAI220     u0465(.A0(men_men_n487_), .A1(men_men_n486_), .B0(men_men_n483_), .B1(men_men_n480_), .Y(men_men_n488_));
  NA2        u0466(.A(men_men_n256_), .B(men_men_n317_), .Y(men_men_n489_));
  NO3        u0467(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n490_));
  INV        u0468(.A(men_men_n490_), .Y(men_men_n491_));
  NA3        u0469(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n492_));
  NA4        u0470(.A(men_men_n145_), .B(men_men_n115_), .C(men_men_n80_), .D(men_men_n23_), .Y(men_men_n493_));
  OAI220     u0471(.A0(men_men_n493_), .A1(men_men_n492_), .B0(men_men_n491_), .B1(men_men_n489_), .Y(men_men_n494_));
  NO3        u0472(.A(men_men_n494_), .B(men_men_n488_), .C(men_men_n479_), .Y(men_men_n495_));
  NA2        u0473(.A(men_men_n304_), .B(men_men_n109_), .Y(men_men_n496_));
  OR2        u0474(.A(men_men_n496_), .B(men_men_n211_), .Y(men_men_n497_));
  OR2        u0475(.A(men_men_n367_), .B(men_men_n104_), .Y(men_men_n498_));
  OA220      u0476(.A0(men_men_n498_), .A1(men_men_n163_), .B0(men_men_n497_), .B1(men_men_n236_), .Y(men_men_n499_));
  NA2        u0477(.A(men_men_n99_), .B(i_13_), .Y(men_men_n500_));
  NA2        u0478(.A(men_men_n454_), .B(men_men_n402_), .Y(men_men_n501_));
  NO2        u0479(.A(i_2_), .B(i_13_), .Y(men_men_n502_));
  NO2        u0480(.A(men_men_n501_), .B(men_men_n500_), .Y(men_men_n503_));
  NO3        u0481(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n504_));
  NO2        u0482(.A(i_6_), .B(i_7_), .Y(men_men_n505_));
  NA2        u0483(.A(men_men_n505_), .B(men_men_n504_), .Y(men_men_n506_));
  NO2        u0484(.A(i_11_), .B(i_1_), .Y(men_men_n507_));
  NO2        u0485(.A(men_men_n73_), .B(i_3_), .Y(men_men_n508_));
  OR2        u0486(.A(i_11_), .B(i_8_), .Y(men_men_n509_));
  NOi21      u0487(.An(i_2_), .B(i_7_), .Y(men_men_n510_));
  NAi31      u0488(.An(men_men_n509_), .B(men_men_n510_), .C(men_men_n508_), .Y(men_men_n511_));
  NO2        u0489(.A(men_men_n441_), .B(i_6_), .Y(men_men_n512_));
  NA3        u0490(.A(men_men_n512_), .B(men_men_n472_), .C(men_men_n75_), .Y(men_men_n513_));
  NO2        u0491(.A(men_men_n513_), .B(men_men_n511_), .Y(men_men_n514_));
  NO2        u0492(.A(i_3_), .B(men_men_n195_), .Y(men_men_n515_));
  NO2        u0493(.A(i_6_), .B(i_10_), .Y(men_men_n516_));
  NA3        u0494(.A(men_men_n516_), .B(men_men_n322_), .C(men_men_n515_), .Y(men_men_n517_));
  NO2        u0495(.A(men_men_n517_), .B(men_men_n156_), .Y(men_men_n518_));
  NA3        u0496(.A(men_men_n250_), .B(men_men_n173_), .C(men_men_n132_), .Y(men_men_n519_));
  NA2        u0497(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n520_));
  NO2        u0498(.A(men_men_n158_), .B(i_3_), .Y(men_men_n521_));
  NAi31      u0499(.An(men_men_n520_), .B(men_men_n521_), .C(men_men_n231_), .Y(men_men_n522_));
  NA3        u0500(.A(men_men_n415_), .B(men_men_n181_), .C(men_men_n149_), .Y(men_men_n523_));
  NA3        u0501(.A(men_men_n523_), .B(men_men_n522_), .C(men_men_n519_), .Y(men_men_n524_));
  NO4        u0502(.A(men_men_n524_), .B(men_men_n518_), .C(men_men_n514_), .D(men_men_n503_), .Y(men_men_n525_));
  NA2        u0503(.A(men_men_n481_), .B(men_men_n403_), .Y(men_men_n526_));
  NA2        u0504(.A(men_men_n490_), .B(men_men_n410_), .Y(men_men_n527_));
  NO2        u0505(.A(men_men_n527_), .B(men_men_n229_), .Y(men_men_n528_));
  NAi21      u0506(.An(men_men_n220_), .B(men_men_n421_), .Y(men_men_n529_));
  NO2        u0507(.A(men_men_n26_), .B(i_5_), .Y(men_men_n530_));
  NO2        u0508(.A(i_0_), .B(men_men_n86_), .Y(men_men_n531_));
  NA3        u0509(.A(men_men_n531_), .B(men_men_n530_), .C(men_men_n142_), .Y(men_men_n532_));
  OR3        u0510(.A(men_men_n312_), .B(men_men_n38_), .C(men_men_n46_), .Y(men_men_n533_));
  NO2        u0511(.A(men_men_n533_), .B(men_men_n532_), .Y(men_men_n534_));
  NA2        u0512(.A(men_men_n27_), .B(i_10_), .Y(men_men_n535_));
  NA2        u0513(.A(men_men_n322_), .B(men_men_n243_), .Y(men_men_n536_));
  OAI220     u0514(.A0(men_men_n536_), .A1(men_men_n462_), .B0(men_men_n535_), .B1(men_men_n500_), .Y(men_men_n537_));
  NA4        u0515(.A(men_men_n315_), .B(men_men_n228_), .C(men_men_n73_), .D(men_men_n241_), .Y(men_men_n538_));
  NO2        u0516(.A(men_men_n538_), .B(men_men_n506_), .Y(men_men_n539_));
  NO4        u0517(.A(men_men_n539_), .B(men_men_n537_), .C(men_men_n534_), .D(men_men_n528_), .Y(men_men_n540_));
  NA4        u0518(.A(men_men_n540_), .B(men_men_n525_), .C(men_men_n499_), .D(men_men_n495_), .Y(men_men_n541_));
  NA3        u0519(.A(men_men_n315_), .B(men_men_n178_), .C(men_men_n176_), .Y(men_men_n542_));
  OAI210     u0520(.A0(men_men_n310_), .A1(men_men_n183_), .B0(men_men_n542_), .Y(men_men_n543_));
  AN2        u0521(.A(men_men_n295_), .B(men_men_n238_), .Y(men_men_n544_));
  NA2        u0522(.A(men_men_n544_), .B(men_men_n543_), .Y(men_men_n545_));
  NA2        u0523(.A(men_men_n122_), .B(men_men_n112_), .Y(men_men_n546_));
  AN2        u0524(.A(men_men_n546_), .B(men_men_n481_), .Y(men_men_n547_));
  NA2        u0525(.A(men_men_n322_), .B(men_men_n165_), .Y(men_men_n548_));
  OAI210     u0526(.A0(men_men_n548_), .A1(men_men_n236_), .B0(men_men_n316_), .Y(men_men_n549_));
  AOI220     u0527(.A0(men_men_n549_), .A1(men_men_n334_), .B0(men_men_n547_), .B1(men_men_n318_), .Y(men_men_n550_));
  NA2        u0528(.A(men_men_n403_), .B(men_men_n230_), .Y(men_men_n551_));
  NA2        u0529(.A(men_men_n372_), .B(men_men_n73_), .Y(men_men_n552_));
  NA2        u0530(.A(men_men_n390_), .B(men_men_n382_), .Y(men_men_n553_));
  AO210      u0531(.A0(men_men_n552_), .A1(men_men_n551_), .B0(men_men_n553_), .Y(men_men_n554_));
  NO2        u0532(.A(men_men_n36_), .B(i_8_), .Y(men_men_n555_));
  NAi41      u0533(.An(men_men_n552_), .B(men_men_n516_), .C(men_men_n555_), .D(men_men_n46_), .Y(men_men_n556_));
  INV        u0534(.A(men_men_n442_), .Y(men_men_n557_));
  NA3        u0535(.A(men_men_n557_), .B(men_men_n556_), .C(men_men_n554_), .Y(men_men_n558_));
  INV        u0536(.A(men_men_n558_), .Y(men_men_n559_));
  NA2        u0537(.A(men_men_n263_), .B(men_men_n64_), .Y(men_men_n560_));
  OAI210     u0538(.A0(i_8_), .A1(men_men_n560_), .B0(men_men_n134_), .Y(men_men_n561_));
  AOI210     u0539(.A0(men_men_n196_), .A1(i_9_), .B0(men_men_n274_), .Y(men_men_n562_));
  NO2        u0540(.A(men_men_n562_), .B(men_men_n201_), .Y(men_men_n563_));
  OR2        u0541(.A(men_men_n185_), .B(i_4_), .Y(men_men_n564_));
  NO2        u0542(.A(men_men_n564_), .B(men_men_n86_), .Y(men_men_n565_));
  AOI220     u0543(.A0(men_men_n565_), .A1(men_men_n563_), .B0(men_men_n561_), .B1(men_men_n443_), .Y(men_men_n566_));
  NA4        u0544(.A(men_men_n566_), .B(men_men_n559_), .C(men_men_n550_), .D(men_men_n545_), .Y(men_men_n567_));
  NA2        u0545(.A(men_men_n409_), .B(men_men_n304_), .Y(men_men_n568_));
  NA2        u0546(.A(men_men_n170_), .B(men_men_n568_), .Y(men_men_n569_));
  NO2        u0547(.A(i_12_), .B(men_men_n195_), .Y(men_men_n570_));
  NA2        u0548(.A(men_men_n570_), .B(men_men_n230_), .Y(men_men_n571_));
  NA3        u0549(.A(men_men_n516_), .B(men_men_n176_), .C(men_men_n27_), .Y(men_men_n572_));
  NO3        u0550(.A(men_men_n572_), .B(men_men_n571_), .C(men_men_n496_), .Y(men_men_n573_));
  NOi31      u0551(.An(men_men_n325_), .B(men_men_n441_), .C(men_men_n38_), .Y(men_men_n574_));
  OAI210     u0552(.A0(men_men_n574_), .A1(men_men_n573_), .B0(men_men_n569_), .Y(men_men_n575_));
  NO2        u0553(.A(i_8_), .B(i_7_), .Y(men_men_n576_));
  OAI210     u0554(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n577_));
  NA2        u0555(.A(men_men_n577_), .B(men_men_n228_), .Y(men_men_n578_));
  AOI220     u0556(.A0(men_men_n335_), .A1(men_men_n39_), .B0(men_men_n239_), .B1(men_men_n210_), .Y(men_men_n579_));
  OAI220     u0557(.A0(men_men_n579_), .A1(men_men_n564_), .B0(men_men_n578_), .B1(men_men_n247_), .Y(men_men_n580_));
  NA2        u0558(.A(men_men_n44_), .B(i_10_), .Y(men_men_n581_));
  NO2        u0559(.A(men_men_n581_), .B(i_6_), .Y(men_men_n582_));
  NA3        u0560(.A(men_men_n582_), .B(men_men_n580_), .C(men_men_n576_), .Y(men_men_n583_));
  AOI220     u0561(.A0(men_men_n454_), .A1(men_men_n335_), .B0(men_men_n252_), .B1(men_men_n249_), .Y(men_men_n584_));
  OAI220     u0562(.A0(men_men_n584_), .A1(men_men_n271_), .B0(men_men_n500_), .B1(men_men_n133_), .Y(men_men_n585_));
  NA2        u0563(.A(men_men_n585_), .B(men_men_n274_), .Y(men_men_n586_));
  NOi31      u0564(.An(men_men_n299_), .B(men_men_n310_), .C(men_men_n183_), .Y(men_men_n587_));
  NA3        u0565(.A(men_men_n315_), .B(men_men_n176_), .C(men_men_n99_), .Y(men_men_n588_));
  NO2        u0566(.A(men_men_n226_), .B(men_men_n44_), .Y(men_men_n589_));
  NO2        u0567(.A(men_men_n158_), .B(i_5_), .Y(men_men_n590_));
  NA3        u0568(.A(men_men_n590_), .B(men_men_n431_), .C(men_men_n328_), .Y(men_men_n591_));
  OAI210     u0569(.A0(men_men_n591_), .A1(men_men_n589_), .B0(men_men_n588_), .Y(men_men_n592_));
  OAI210     u0570(.A0(men_men_n592_), .A1(men_men_n587_), .B0(men_men_n490_), .Y(men_men_n593_));
  NA4        u0571(.A(men_men_n593_), .B(men_men_n586_), .C(men_men_n583_), .D(men_men_n575_), .Y(men_men_n594_));
  NA3        u0572(.A(men_men_n222_), .B(men_men_n71_), .C(men_men_n44_), .Y(men_men_n595_));
  NA2        u0573(.A(men_men_n292_), .B(men_men_n84_), .Y(men_men_n596_));
  AOI210     u0574(.A0(men_men_n595_), .A1(men_men_n362_), .B0(men_men_n596_), .Y(men_men_n597_));
  NA2        u0575(.A(men_men_n305_), .B(men_men_n295_), .Y(men_men_n598_));
  NO2        u0576(.A(men_men_n598_), .B(men_men_n175_), .Y(men_men_n599_));
  NA2        u0577(.A(men_men_n228_), .B(men_men_n227_), .Y(men_men_n600_));
  NA2        u0578(.A(men_men_n474_), .B(men_men_n226_), .Y(men_men_n601_));
  NO2        u0579(.A(men_men_n600_), .B(men_men_n601_), .Y(men_men_n602_));
  NA2        u0580(.A(i_0_), .B(men_men_n48_), .Y(men_men_n603_));
  NA3        u0581(.A(men_men_n570_), .B(men_men_n283_), .C(men_men_n603_), .Y(men_men_n604_));
  NO2        u0582(.A(men_men_n1110_), .B(men_men_n604_), .Y(men_men_n605_));
  NO4        u0583(.A(men_men_n605_), .B(men_men_n602_), .C(men_men_n599_), .D(men_men_n597_), .Y(men_men_n606_));
  NO4        u0584(.A(men_men_n257_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n607_));
  NO3        u0585(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n608_));
  NO2        u0586(.A(men_men_n237_), .B(men_men_n36_), .Y(men_men_n609_));
  AN2        u0587(.A(men_men_n609_), .B(men_men_n608_), .Y(men_men_n610_));
  OA210      u0588(.A0(men_men_n610_), .A1(men_men_n607_), .B0(men_men_n372_), .Y(men_men_n611_));
  NO2        u0589(.A(men_men_n441_), .B(i_1_), .Y(men_men_n612_));
  NOi31      u0590(.An(men_men_n612_), .B(men_men_n482_), .C(men_men_n73_), .Y(men_men_n613_));
  AN4        u0591(.A(men_men_n613_), .B(men_men_n438_), .C(men_men_n530_), .D(i_2_), .Y(men_men_n614_));
  NO2        u0592(.A(men_men_n452_), .B(men_men_n179_), .Y(men_men_n615_));
  NO3        u0593(.A(men_men_n615_), .B(men_men_n614_), .C(men_men_n611_), .Y(men_men_n616_));
  NOi21      u0594(.An(i_10_), .B(i_6_), .Y(men_men_n617_));
  NO2        u0595(.A(men_men_n86_), .B(men_men_n25_), .Y(men_men_n618_));
  AOI220     u0596(.A0(men_men_n292_), .A1(men_men_n618_), .B0(men_men_n283_), .B1(men_men_n617_), .Y(men_men_n619_));
  NO2        u0597(.A(men_men_n619_), .B(men_men_n480_), .Y(men_men_n620_));
  NO2        u0598(.A(men_men_n114_), .B(men_men_n23_), .Y(men_men_n621_));
  NA2        u0599(.A(men_men_n325_), .B(men_men_n165_), .Y(men_men_n622_));
  AOI220     u0600(.A0(men_men_n622_), .A1(men_men_n463_), .B0(men_men_n186_), .B1(men_men_n184_), .Y(men_men_n623_));
  NO2        u0601(.A(men_men_n200_), .B(men_men_n37_), .Y(men_men_n624_));
  NOi31      u0602(.An(men_men_n146_), .B(men_men_n624_), .C(men_men_n343_), .Y(men_men_n625_));
  NO3        u0603(.A(men_men_n625_), .B(men_men_n623_), .C(men_men_n620_), .Y(men_men_n626_));
  NO2        u0604(.A(men_men_n552_), .B(men_men_n398_), .Y(men_men_n627_));
  INV        u0605(.A(men_men_n328_), .Y(men_men_n628_));
  NO2        u0606(.A(i_12_), .B(men_men_n86_), .Y(men_men_n629_));
  NA3        u0607(.A(men_men_n629_), .B(men_men_n283_), .C(men_men_n603_), .Y(men_men_n630_));
  NA3        u0608(.A(men_men_n406_), .B(men_men_n292_), .C(men_men_n222_), .Y(men_men_n631_));
  AOI210     u0609(.A0(men_men_n631_), .A1(men_men_n630_), .B0(men_men_n628_), .Y(men_men_n632_));
  NA2        u0610(.A(men_men_n176_), .B(i_0_), .Y(men_men_n633_));
  NO3        u0611(.A(men_men_n633_), .B(men_men_n354_), .C(men_men_n310_), .Y(men_men_n634_));
  OR2        u0612(.A(i_2_), .B(i_5_), .Y(men_men_n635_));
  OR2        u0613(.A(men_men_n635_), .B(men_men_n434_), .Y(men_men_n636_));
  AOI210     u0614(.A0(men_men_n392_), .A1(men_men_n249_), .B0(men_men_n200_), .Y(men_men_n637_));
  AOI210     u0615(.A0(men_men_n637_), .A1(men_men_n636_), .B0(men_men_n529_), .Y(men_men_n638_));
  NO4        u0616(.A(men_men_n638_), .B(men_men_n634_), .C(men_men_n632_), .D(men_men_n627_), .Y(men_men_n639_));
  NA4        u0617(.A(men_men_n639_), .B(men_men_n626_), .C(men_men_n616_), .D(men_men_n606_), .Y(men_men_n640_));
  NO4        u0618(.A(men_men_n640_), .B(men_men_n594_), .C(men_men_n567_), .D(men_men_n541_), .Y(men_men_n641_));
  NA4        u0619(.A(men_men_n641_), .B(men_men_n471_), .C(men_men_n371_), .D(men_men_n321_), .Y(men7));
  NO2        u0620(.A(men_men_n109_), .B(men_men_n92_), .Y(men_men_n643_));
  NA2        u0621(.A(men_men_n404_), .B(men_men_n643_), .Y(men_men_n644_));
  NA2        u0622(.A(men_men_n516_), .B(men_men_n84_), .Y(men_men_n645_));
  OAI210     u0623(.A0(men_men_n1111_), .A1(men_men_n645_), .B0(men_men_n644_), .Y(men_men_n646_));
  NA3        u0624(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n647_));
  NO2        u0625(.A(men_men_n241_), .B(i_4_), .Y(men_men_n648_));
  NA2        u0626(.A(men_men_n648_), .B(i_8_), .Y(men_men_n649_));
  AOI210     u0627(.A0(men_men_n649_), .A1(men_men_n108_), .B0(men_men_n647_), .Y(men_men_n650_));
  NA2        u0628(.A(i_2_), .B(men_men_n86_), .Y(men_men_n651_));
  OAI210     u0629(.A0(men_men_n89_), .A1(men_men_n205_), .B0(men_men_n206_), .Y(men_men_n652_));
  NO2        u0630(.A(i_7_), .B(men_men_n37_), .Y(men_men_n653_));
  NA2        u0631(.A(i_4_), .B(i_8_), .Y(men_men_n654_));
  AOI210     u0632(.A0(men_men_n654_), .A1(men_men_n315_), .B0(men_men_n653_), .Y(men_men_n655_));
  OAI220     u0633(.A0(men_men_n655_), .A1(men_men_n651_), .B0(men_men_n652_), .B1(i_13_), .Y(men_men_n656_));
  NO3        u0634(.A(men_men_n656_), .B(men_men_n650_), .C(men_men_n646_), .Y(men_men_n657_));
  AOI210     u0635(.A0(men_men_n128_), .A1(men_men_n62_), .B0(i_10_), .Y(men_men_n658_));
  AOI210     u0636(.A0(men_men_n658_), .A1(men_men_n241_), .B0(men_men_n162_), .Y(men_men_n659_));
  OR2        u0637(.A(i_6_), .B(i_10_), .Y(men_men_n660_));
  NO2        u0638(.A(men_men_n660_), .B(men_men_n23_), .Y(men_men_n661_));
  OR3        u0639(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n662_));
  NO3        u0640(.A(men_men_n662_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n663_));
  INV        u0641(.A(men_men_n202_), .Y(men_men_n664_));
  OR2        u0642(.A(men_men_n659_), .B(men_men_n276_), .Y(men_men_n665_));
  AOI210     u0643(.A0(men_men_n665_), .A1(men_men_n657_), .B0(men_men_n63_), .Y(men_men_n666_));
  NOi21      u0644(.An(i_11_), .B(i_7_), .Y(men_men_n667_));
  AO210      u0645(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n668_));
  NO2        u0646(.A(men_men_n668_), .B(men_men_n667_), .Y(men_men_n669_));
  NA2        u0647(.A(men_men_n669_), .B(men_men_n210_), .Y(men_men_n670_));
  NA3        u0648(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n671_));
  NAi31      u0649(.An(men_men_n671_), .B(men_men_n219_), .C(i_11_), .Y(men_men_n672_));
  AOI210     u0650(.A0(men_men_n672_), .A1(men_men_n670_), .B0(men_men_n63_), .Y(men_men_n673_));
  NO3        u0651(.A(men_men_n265_), .B(men_men_n212_), .C(i_8_), .Y(men_men_n674_));
  OAI210     u0652(.A0(men_men_n674_), .A1(men_men_n231_), .B0(men_men_n63_), .Y(men_men_n675_));
  NA2        u0653(.A(men_men_n435_), .B(men_men_n31_), .Y(men_men_n676_));
  OR2        u0654(.A(men_men_n212_), .B(men_men_n109_), .Y(men_men_n677_));
  INV        u0655(.A(men_men_n676_), .Y(men_men_n678_));
  NO2        u0656(.A(men_men_n63_), .B(i_9_), .Y(men_men_n679_));
  NO2        u0657(.A(men_men_n679_), .B(i_4_), .Y(men_men_n680_));
  NA2        u0658(.A(men_men_n680_), .B(men_men_n678_), .Y(men_men_n681_));
  NO2        u0659(.A(i_1_), .B(i_12_), .Y(men_men_n682_));
  NA3        u0660(.A(men_men_n682_), .B(men_men_n111_), .C(men_men_n24_), .Y(men_men_n683_));
  NA4        u0661(.A(men_men_n683_), .B(men_men_n681_), .C(men_men_n675_), .D(men_men_n398_), .Y(men_men_n684_));
  OAI210     u0662(.A0(men_men_n684_), .A1(men_men_n673_), .B0(i_6_), .Y(men_men_n685_));
  OAI210     u0663(.A0(men_men_n671_), .A1(men_men_n109_), .B0(men_men_n492_), .Y(men_men_n686_));
  NA2        u0664(.A(men_men_n686_), .B(men_men_n629_), .Y(men_men_n687_));
  NO2        u0665(.A(men_men_n241_), .B(men_men_n86_), .Y(men_men_n688_));
  NO2        u0666(.A(men_men_n688_), .B(i_11_), .Y(men_men_n689_));
  INV        u0667(.A(men_men_n687_), .Y(men_men_n690_));
  NO4        u0668(.A(men_men_n219_), .B(men_men_n128_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n691_));
  NA2        u0669(.A(men_men_n691_), .B(men_men_n679_), .Y(men_men_n692_));
  NA2        u0670(.A(men_men_n241_), .B(i_6_), .Y(men_men_n693_));
  NO3        u0671(.A(men_men_n660_), .B(men_men_n237_), .C(men_men_n23_), .Y(men_men_n694_));
  AOI210     u0672(.A0(i_1_), .A1(men_men_n266_), .B0(men_men_n694_), .Y(men_men_n695_));
  OAI210     u0673(.A0(men_men_n695_), .A1(men_men_n44_), .B0(men_men_n692_), .Y(men_men_n696_));
  NA3        u0674(.A(men_men_n576_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n697_));
  NA3        u0675(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n698_));
  NO2        u0676(.A(men_men_n46_), .B(i_1_), .Y(men_men_n699_));
  NA3        u0677(.A(men_men_n699_), .B(men_men_n275_), .C(men_men_n44_), .Y(men_men_n700_));
  NO2        u0678(.A(men_men_n700_), .B(men_men_n698_), .Y(men_men_n701_));
  NA3        u0679(.A(men_men_n679_), .B(men_men_n328_), .C(i_6_), .Y(men_men_n702_));
  NO2        u0680(.A(men_men_n702_), .B(men_men_n23_), .Y(men_men_n703_));
  AOI210     u0681(.A0(men_men_n507_), .A1(men_men_n445_), .B0(men_men_n246_), .Y(men_men_n704_));
  NO2        u0682(.A(men_men_n704_), .B(men_men_n651_), .Y(men_men_n705_));
  NAi21      u0683(.An(men_men_n697_), .B(men_men_n94_), .Y(men_men_n706_));
  NA2        u0684(.A(men_men_n699_), .B(men_men_n275_), .Y(men_men_n707_));
  NO2        u0685(.A(i_11_), .B(men_men_n37_), .Y(men_men_n708_));
  NA2        u0686(.A(men_men_n708_), .B(men_men_n24_), .Y(men_men_n709_));
  OAI210     u0687(.A0(men_men_n709_), .A1(men_men_n707_), .B0(men_men_n706_), .Y(men_men_n710_));
  OR4        u0688(.A(men_men_n710_), .B(men_men_n705_), .C(men_men_n703_), .D(men_men_n701_), .Y(men_men_n711_));
  NO3        u0689(.A(men_men_n711_), .B(men_men_n696_), .C(men_men_n690_), .Y(men_men_n712_));
  INV        u0690(.A(i_1_), .Y(men_men_n713_));
  NO2        u0691(.A(men_men_n713_), .B(men_men_n662_), .Y(men_men_n714_));
  NO2        u0692(.A(men_men_n440_), .B(men_men_n86_), .Y(men_men_n715_));
  NA2        u0693(.A(men_men_n714_), .B(men_men_n46_), .Y(men_men_n716_));
  NA2        u0694(.A(i_3_), .B(men_men_n195_), .Y(men_men_n717_));
  NO2        u0695(.A(men_men_n717_), .B(men_men_n114_), .Y(men_men_n718_));
  AN2        u0696(.A(men_men_n718_), .B(men_men_n582_), .Y(men_men_n719_));
  NO2        u0697(.A(men_men_n237_), .B(men_men_n44_), .Y(men_men_n720_));
  NO3        u0698(.A(men_men_n720_), .B(men_men_n318_), .C(men_men_n242_), .Y(men_men_n721_));
  NO2        u0699(.A(men_men_n117_), .B(men_men_n37_), .Y(men_men_n722_));
  NO2        u0700(.A(men_men_n722_), .B(i_6_), .Y(men_men_n723_));
  NO2        u0701(.A(men_men_n86_), .B(i_9_), .Y(men_men_n724_));
  NO2        u0702(.A(men_men_n724_), .B(men_men_n63_), .Y(men_men_n725_));
  NO2        u0703(.A(men_men_n725_), .B(men_men_n682_), .Y(men_men_n726_));
  NO4        u0704(.A(men_men_n726_), .B(men_men_n723_), .C(men_men_n721_), .D(i_4_), .Y(men_men_n727_));
  NA2        u0705(.A(i_1_), .B(i_3_), .Y(men_men_n728_));
  NO2        u0706(.A(men_men_n484_), .B(men_men_n95_), .Y(men_men_n729_));
  INV        u0707(.A(men_men_n729_), .Y(men_men_n730_));
  NO2        u0708(.A(men_men_n730_), .B(men_men_n728_), .Y(men_men_n731_));
  NO3        u0709(.A(men_men_n731_), .B(men_men_n727_), .C(men_men_n719_), .Y(men_men_n732_));
  NA4        u0710(.A(men_men_n732_), .B(men_men_n716_), .C(men_men_n712_), .D(men_men_n685_), .Y(men_men_n733_));
  NO3        u0711(.A(men_men_n509_), .B(i_3_), .C(i_7_), .Y(men_men_n734_));
  NOi21      u0712(.An(men_men_n734_), .B(i_10_), .Y(men_men_n735_));
  OA210      u0713(.A0(men_men_n735_), .A1(men_men_n250_), .B0(men_men_n86_), .Y(men_men_n736_));
  NA2        u0714(.A(men_men_n390_), .B(men_men_n389_), .Y(men_men_n737_));
  NO3        u0715(.A(men_men_n510_), .B(men_men_n654_), .C(men_men_n86_), .Y(men_men_n738_));
  NA2        u0716(.A(men_men_n738_), .B(men_men_n25_), .Y(men_men_n739_));
  NA2        u0717(.A(men_men_n162_), .B(men_men_n86_), .Y(men_men_n740_));
  NA3        u0718(.A(men_men_n740_), .B(men_men_n739_), .C(men_men_n737_), .Y(men_men_n741_));
  OAI210     u0719(.A0(men_men_n741_), .A1(men_men_n736_), .B0(i_1_), .Y(men_men_n742_));
  NO2        u0720(.A(men_men_n702_), .B(men_men_n475_), .Y(men_men_n743_));
  INV        u0721(.A(men_men_n743_), .Y(men_men_n744_));
  AOI210     u0722(.A0(men_men_n744_), .A1(men_men_n742_), .B0(i_13_), .Y(men_men_n745_));
  OR2        u0723(.A(i_11_), .B(i_7_), .Y(men_men_n746_));
  NA3        u0724(.A(men_men_n746_), .B(i_3_), .C(men_men_n138_), .Y(men_men_n747_));
  AOI220     u0725(.A0(men_men_n502_), .A1(men_men_n162_), .B0(men_men_n477_), .B1(men_men_n138_), .Y(men_men_n748_));
  NA2        u0726(.A(men_men_n748_), .B(men_men_n747_), .Y(men_men_n749_));
  NO2        u0727(.A(men_men_n510_), .B(men_men_n24_), .Y(men_men_n750_));
  AOI210     u0728(.A0(men_men_n750_), .A1(men_men_n715_), .B0(men_men_n250_), .Y(men_men_n751_));
  OAI220     u0729(.A0(men_men_n751_), .A1(men_men_n40_), .B0(men_men_n54_), .B1(men_men_n95_), .Y(men_men_n752_));
  AOI210     u0730(.A0(men_men_n749_), .A1(men_men_n345_), .B0(men_men_n752_), .Y(men_men_n753_));
  NA2        u0731(.A(men_men_n114_), .B(men_men_n109_), .Y(men_men_n754_));
  AOI220     u0732(.A0(men_men_n754_), .A1(men_men_n72_), .B0(men_men_n406_), .B1(men_men_n699_), .Y(men_men_n755_));
  NO2        u0733(.A(men_men_n755_), .B(men_men_n247_), .Y(men_men_n756_));
  AOI210     u0734(.A0(men_men_n475_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n757_));
  NOi21      u0735(.An(men_men_n757_), .B(men_men_n645_), .Y(men_men_n758_));
  NA2        u0736(.A(men_men_n127_), .B(i_13_), .Y(men_men_n759_));
  NO2        u0737(.A(men_men_n698_), .B(men_men_n114_), .Y(men_men_n760_));
  INV        u0738(.A(men_men_n760_), .Y(men_men_n761_));
  OAI220     u0739(.A0(men_men_n761_), .A1(men_men_n71_), .B0(men_men_n759_), .B1(men_men_n1112_), .Y(men_men_n762_));
  NO3        u0740(.A(men_men_n71_), .B(men_men_n32_), .C(men_men_n104_), .Y(men_men_n763_));
  NA2        u0741(.A(men_men_n26_), .B(men_men_n195_), .Y(men_men_n764_));
  INV        u0742(.A(men_men_n763_), .Y(men_men_n765_));
  AOI220     u0743(.A0(men_men_n406_), .A1(men_men_n699_), .B0(men_men_n94_), .B1(men_men_n105_), .Y(men_men_n766_));
  OAI220     u0744(.A0(men_men_n766_), .A1(men_men_n649_), .B0(men_men_n765_), .B1(men_men_n664_), .Y(men_men_n767_));
  NO4        u0745(.A(men_men_n767_), .B(men_men_n762_), .C(men_men_n758_), .D(men_men_n756_), .Y(men_men_n768_));
  OR2        u0746(.A(i_11_), .B(i_6_), .Y(men_men_n769_));
  NA3        u0747(.A(men_men_n648_), .B(men_men_n764_), .C(i_7_), .Y(men_men_n770_));
  AOI210     u0748(.A0(men_men_n770_), .A1(men_men_n761_), .B0(men_men_n769_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n689_), .B(i_13_), .Y(men_men_n772_));
  NA2        u0750(.A(men_men_n105_), .B(men_men_n764_), .Y(men_men_n773_));
  NAi21      u0751(.An(i_11_), .B(i_12_), .Y(men_men_n774_));
  NO3        u0752(.A(men_men_n774_), .B(i_13_), .C(men_men_n86_), .Y(men_men_n775_));
  NO3        u0753(.A(men_men_n510_), .B(men_men_n629_), .C(men_men_n654_), .Y(men_men_n776_));
  AOI220     u0754(.A0(men_men_n776_), .A1(men_men_n322_), .B0(men_men_n775_), .B1(men_men_n773_), .Y(men_men_n777_));
  NA2        u0755(.A(men_men_n777_), .B(men_men_n772_), .Y(men_men_n778_));
  OAI210     u0756(.A0(men_men_n778_), .A1(men_men_n771_), .B0(men_men_n63_), .Y(men_men_n779_));
  NO2        u0757(.A(i_2_), .B(i_12_), .Y(men_men_n780_));
  NA2        u0758(.A(men_men_n387_), .B(men_men_n780_), .Y(men_men_n781_));
  OAI210     u0759(.A0(i_8_), .A1(men_men_n389_), .B0(men_men_n387_), .Y(men_men_n782_));
  NO2        u0760(.A(men_men_n128_), .B(i_2_), .Y(men_men_n783_));
  NA2        u0761(.A(men_men_n783_), .B(men_men_n682_), .Y(men_men_n784_));
  NA3        u0762(.A(men_men_n784_), .B(men_men_n782_), .C(men_men_n781_), .Y(men_men_n785_));
  NA3        u0763(.A(men_men_n785_), .B(men_men_n45_), .C(men_men_n230_), .Y(men_men_n786_));
  NA4        u0764(.A(men_men_n786_), .B(men_men_n779_), .C(men_men_n768_), .D(men_men_n753_), .Y(men_men_n787_));
  OR4        u0765(.A(men_men_n787_), .B(men_men_n745_), .C(men_men_n733_), .D(men_men_n666_), .Y(men5));
  NA3        u0766(.A(men_men_n24_), .B(men_men_n780_), .C(men_men_n109_), .Y(men_men_n789_));
  NO2        u0767(.A(men_men_n649_), .B(i_11_), .Y(men_men_n790_));
  NA2        u0768(.A(men_men_n89_), .B(men_men_n790_), .Y(men_men_n791_));
  NA2        u0769(.A(men_men_n791_), .B(men_men_n789_), .Y(men_men_n792_));
  NO3        u0770(.A(i_11_), .B(men_men_n241_), .C(i_13_), .Y(men_men_n793_));
  NO2        u0771(.A(men_men_n124_), .B(men_men_n23_), .Y(men_men_n794_));
  NA2        u0772(.A(i_12_), .B(i_8_), .Y(men_men_n795_));
  INV        u0773(.A(men_men_n474_), .Y(men_men_n796_));
  NA2        u0774(.A(men_men_n1116_), .B(men_men_n794_), .Y(men_men_n797_));
  INV        u0775(.A(men_men_n797_), .Y(men_men_n798_));
  NO2        u0776(.A(men_men_n798_), .B(men_men_n792_), .Y(men_men_n799_));
  INV        u0777(.A(men_men_n173_), .Y(men_men_n800_));
  INV        u0778(.A(men_men_n250_), .Y(men_men_n801_));
  INV        u0779(.A(men_men_n476_), .Y(men_men_n802_));
  AOI210     u0780(.A0(men_men_n802_), .A1(men_men_n801_), .B0(men_men_n800_), .Y(men_men_n803_));
  NO2        u0781(.A(men_men_n484_), .B(men_men_n26_), .Y(men_men_n804_));
  NO2        u0782(.A(men_men_n804_), .B(men_men_n445_), .Y(men_men_n805_));
  INV        u0783(.A(men_men_n803_), .Y(men_men_n806_));
  INV        u0784(.A(men_men_n794_), .Y(men_men_n807_));
  INV        u0785(.A(men_men_n174_), .Y(men_men_n808_));
  NO3        u0786(.A(men_men_n668_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n809_));
  AOI210     u0787(.A0(men_men_n808_), .A1(men_men_n89_), .B0(men_men_n809_), .Y(men_men_n810_));
  AOI210     u0788(.A0(men_men_n810_), .A1(men_men_n807_), .B0(men_men_n195_), .Y(men_men_n811_));
  OA210      u0789(.A0(men_men_n669_), .A1(men_men_n126_), .B0(i_13_), .Y(men_men_n812_));
  NA2        u0790(.A(men_men_n202_), .B(men_men_n205_), .Y(men_men_n813_));
  NA2        u0791(.A(men_men_n152_), .B(i_8_), .Y(men_men_n814_));
  AOI210     u0792(.A0(men_men_n814_), .A1(men_men_n813_), .B0(men_men_n392_), .Y(men_men_n815_));
  NA2        u0793(.A(men_men_n212_), .B(men_men_n148_), .Y(men_men_n816_));
  NA2        u0794(.A(men_men_n816_), .B(men_men_n445_), .Y(men_men_n817_));
  NO2        u0795(.A(men_men_n105_), .B(men_men_n44_), .Y(men_men_n818_));
  NA3        u0796(.A(men_men_n104_), .B(men_men_n315_), .C(men_men_n42_), .Y(men_men_n819_));
  OAI210     u0797(.A0(men_men_n819_), .A1(men_men_n818_), .B0(men_men_n817_), .Y(men_men_n820_));
  NO4        u0798(.A(men_men_n820_), .B(men_men_n815_), .C(men_men_n812_), .D(men_men_n811_), .Y(men_men_n821_));
  NA2        u0799(.A(men_men_n621_), .B(men_men_n28_), .Y(men_men_n822_));
  NA2        u0800(.A(men_men_n793_), .B(men_men_n284_), .Y(men_men_n823_));
  NA2        u0801(.A(men_men_n823_), .B(men_men_n822_), .Y(men_men_n824_));
  NO2        u0802(.A(men_men_n62_), .B(i_12_), .Y(men_men_n825_));
  INV        u0803(.A(men_men_n824_), .Y(men_men_n826_));
  NA4        u0804(.A(men_men_n826_), .B(men_men_n821_), .C(men_men_n806_), .D(men_men_n799_), .Y(men6));
  NO2        u0805(.A(men_men_n317_), .B(i_1_), .Y(men_men_n828_));
  NO2        u0806(.A(men_men_n188_), .B(men_men_n139_), .Y(men_men_n829_));
  OAI210     u0807(.A0(men_men_n829_), .A1(men_men_n828_), .B0(men_men_n783_), .Y(men_men_n830_));
  NA4        u0808(.A(men_men_n410_), .B(men_men_n515_), .C(men_men_n71_), .D(men_men_n104_), .Y(men_men_n831_));
  INV        u0809(.A(men_men_n831_), .Y(men_men_n832_));
  NO2        u0810(.A(men_men_n225_), .B(men_men_n520_), .Y(men_men_n833_));
  NO2        u0811(.A(men_men_n832_), .B(men_men_n340_), .Y(men_men_n834_));
  AO210      u0812(.A0(men_men_n834_), .A1(men_men_n830_), .B0(i_12_), .Y(men_men_n835_));
  NA2        u0813(.A(men_men_n393_), .B(men_men_n348_), .Y(men_men_n836_));
  NA2        u0814(.A(men_men_n735_), .B(men_men_n71_), .Y(men_men_n837_));
  NA2        u0815(.A(men_men_n837_), .B(men_men_n836_), .Y(men_men_n838_));
  INV        u0816(.A(men_men_n199_), .Y(men_men_n839_));
  NO2        u0817(.A(men_men_n838_), .B(men_men_n839_), .Y(men_men_n840_));
  INV        u0818(.A(men_men_n339_), .Y(men_men_n841_));
  NA2        u0819(.A(men_men_n75_), .B(men_men_n131_), .Y(men_men_n842_));
  NO2        u0820(.A(men_men_n842_), .B(men_men_n841_), .Y(men_men_n843_));
  NO3        u0821(.A(men_men_n257_), .B(men_men_n132_), .C(i_9_), .Y(men_men_n844_));
  NA2        u0822(.A(men_men_n844_), .B(men_men_n825_), .Y(men_men_n845_));
  AOI210     u0823(.A0(men_men_n845_), .A1(men_men_n553_), .B0(men_men_n188_), .Y(men_men_n846_));
  NO2        u0824(.A(men_men_n32_), .B(i_11_), .Y(men_men_n847_));
  NAi32      u0825(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n848_));
  AOI210     u0826(.A0(men_men_n769_), .A1(men_men_n87_), .B0(men_men_n848_), .Y(men_men_n849_));
  OAI210     u0827(.A0(men_men_n734_), .A1(men_men_n609_), .B0(men_men_n608_), .Y(men_men_n850_));
  NAi21      u0828(.An(men_men_n849_), .B(men_men_n850_), .Y(men_men_n851_));
  OR3        u0829(.A(men_men_n851_), .B(men_men_n846_), .C(men_men_n843_), .Y(men_men_n852_));
  NO2        u0830(.A(men_men_n746_), .B(i_2_), .Y(men_men_n853_));
  NA2        u0831(.A(men_men_n48_), .B(men_men_n37_), .Y(men_men_n854_));
  OAI210     u0832(.A0(men_men_n854_), .A1(men_men_n434_), .B0(men_men_n377_), .Y(men_men_n855_));
  NA2        u0833(.A(men_men_n855_), .B(men_men_n853_), .Y(men_men_n856_));
  AO220      u0834(.A0(men_men_n376_), .A1(men_men_n366_), .B0(men_men_n418_), .B1(i_8_), .Y(men_men_n857_));
  NA3        u0835(.A(men_men_n857_), .B(men_men_n262_), .C(i_7_), .Y(men_men_n858_));
  OR2        u0836(.A(men_men_n669_), .B(men_men_n476_), .Y(men_men_n859_));
  NA3        u0837(.A(men_men_n859_), .B(men_men_n147_), .C(men_men_n69_), .Y(men_men_n860_));
  OR2        u0838(.A(men_men_n796_), .B(men_men_n36_), .Y(men_men_n861_));
  NA4        u0839(.A(men_men_n861_), .B(men_men_n860_), .C(men_men_n858_), .D(men_men_n856_), .Y(men_men_n862_));
  INV        u0840(.A(men_men_n87_), .Y(men_men_n863_));
  AOI220     u0841(.A0(men_men_n863_), .A1(men_men_n608_), .B0(men_men_n833_), .B1(men_men_n1115_), .Y(men_men_n864_));
  NA3        u0842(.A(men_men_n392_), .B(men_men_n243_), .C(men_men_n147_), .Y(men_men_n865_));
  NA2        u0843(.A(men_men_n418_), .B(men_men_n70_), .Y(men_men_n866_));
  NA4        u0844(.A(men_men_n866_), .B(men_men_n865_), .C(men_men_n864_), .D(men_men_n652_), .Y(men_men_n867_));
  AO210      u0845(.A0(men_men_n555_), .A1(men_men_n46_), .B0(men_men_n88_), .Y(men_men_n868_));
  NA2        u0846(.A(men_men_n868_), .B(men_men_n516_), .Y(men_men_n869_));
  AOI210     u0847(.A0(men_men_n476_), .A1(men_men_n474_), .B0(men_men_n607_), .Y(men_men_n870_));
  NO2        u0848(.A(men_men_n660_), .B(men_men_n105_), .Y(men_men_n871_));
  OAI210     u0849(.A0(men_men_n871_), .A1(men_men_n112_), .B0(men_men_n433_), .Y(men_men_n872_));
  NA2        u0850(.A(men_men_n249_), .B(men_men_n46_), .Y(men_men_n873_));
  INV        u0851(.A(men_men_n636_), .Y(men_men_n874_));
  NA3        u0852(.A(men_men_n874_), .B(men_men_n339_), .C(i_7_), .Y(men_men_n875_));
  NA4        u0853(.A(men_men_n875_), .B(men_men_n872_), .C(men_men_n870_), .D(men_men_n869_), .Y(men_men_n876_));
  NO4        u0854(.A(men_men_n876_), .B(men_men_n867_), .C(men_men_n862_), .D(men_men_n852_), .Y(men_men_n877_));
  NA4        u0855(.A(men_men_n877_), .B(men_men_n840_), .C(men_men_n835_), .D(men_men_n400_), .Y(men3));
  NA2        u0856(.A(i_12_), .B(i_10_), .Y(men_men_n879_));
  NA2        u0857(.A(i_6_), .B(i_7_), .Y(men_men_n880_));
  NO2        u0858(.A(men_men_n880_), .B(i_0_), .Y(men_men_n881_));
  NO2        u0859(.A(i_11_), .B(men_men_n241_), .Y(men_men_n882_));
  OAI210     u0860(.A0(men_men_n881_), .A1(men_men_n299_), .B0(men_men_n882_), .Y(men_men_n883_));
  NO2        u0861(.A(men_men_n883_), .B(men_men_n195_), .Y(men_men_n884_));
  NO3        u0862(.A(men_men_n480_), .B(men_men_n92_), .C(men_men_n44_), .Y(men_men_n885_));
  OA210      u0863(.A0(men_men_n885_), .A1(men_men_n884_), .B0(men_men_n176_), .Y(men_men_n886_));
  NA3        u0864(.A(men_men_n865_), .B(men_men_n652_), .C(men_men_n391_), .Y(men_men_n887_));
  NA2        u0865(.A(men_men_n887_), .B(men_men_n39_), .Y(men_men_n888_));
  NOi21      u0866(.An(men_men_n99_), .B(men_men_n805_), .Y(men_men_n889_));
  NO3        u0867(.A(men_men_n677_), .B(men_men_n484_), .C(men_men_n131_), .Y(men_men_n890_));
  NA2        u0868(.A(men_men_n435_), .B(men_men_n45_), .Y(men_men_n891_));
  AN2        u0869(.A(men_men_n482_), .B(men_men_n55_), .Y(men_men_n892_));
  NO3        u0870(.A(men_men_n892_), .B(men_men_n890_), .C(men_men_n889_), .Y(men_men_n893_));
  AOI210     u0871(.A0(men_men_n893_), .A1(men_men_n888_), .B0(men_men_n48_), .Y(men_men_n894_));
  NO4        u0872(.A(men_men_n396_), .B(men_men_n403_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n895_));
  NA2        u0873(.A(men_men_n188_), .B(men_men_n617_), .Y(men_men_n896_));
  NOi21      u0874(.An(men_men_n896_), .B(men_men_n895_), .Y(men_men_n897_));
  NA2        u0875(.A(men_men_n757_), .B(men_men_n724_), .Y(men_men_n898_));
  NA2        u0876(.A(men_men_n346_), .B(men_men_n465_), .Y(men_men_n899_));
  OAI220     u0877(.A0(men_men_n899_), .A1(men_men_n898_), .B0(men_men_n897_), .B1(men_men_n63_), .Y(men_men_n900_));
  NOi21      u0878(.An(i_5_), .B(i_9_), .Y(men_men_n901_));
  NA2        u0879(.A(men_men_n901_), .B(men_men_n473_), .Y(men_men_n902_));
  INV        u0880(.A(men_men_n738_), .Y(men_men_n903_));
  NO3        u0881(.A(men_men_n1113_), .B(men_men_n275_), .C(men_men_n73_), .Y(men_men_n904_));
  NO2        u0882(.A(men_men_n177_), .B(men_men_n148_), .Y(men_men_n905_));
  AOI210     u0883(.A0(men_men_n905_), .A1(men_men_n249_), .B0(men_men_n904_), .Y(men_men_n906_));
  OAI220     u0884(.A0(men_men_n906_), .A1(men_men_n183_), .B0(men_men_n903_), .B1(men_men_n902_), .Y(men_men_n907_));
  NO4        u0885(.A(men_men_n907_), .B(men_men_n900_), .C(men_men_n894_), .D(men_men_n886_), .Y(men_men_n908_));
  NA2        u0886(.A(men_men_n188_), .B(men_men_n24_), .Y(men_men_n909_));
  NO2        u0887(.A(men_men_n722_), .B(men_men_n643_), .Y(men_men_n910_));
  NO2        u0888(.A(men_men_n910_), .B(men_men_n909_), .Y(men_men_n911_));
  NA2        u0889(.A(men_men_n322_), .B(men_men_n129_), .Y(men_men_n912_));
  NAi21      u0890(.An(men_men_n163_), .B(men_men_n465_), .Y(men_men_n913_));
  OAI220     u0891(.A0(men_men_n913_), .A1(men_men_n873_), .B0(men_men_n912_), .B1(men_men_n424_), .Y(men_men_n914_));
  NO2        u0892(.A(men_men_n914_), .B(men_men_n911_), .Y(men_men_n915_));
  NO2        u0893(.A(men_men_n410_), .B(men_men_n303_), .Y(men_men_n916_));
  NA2        u0894(.A(men_men_n916_), .B(men_men_n760_), .Y(men_men_n917_));
  NO4        u0895(.A(men_men_n635_), .B(men_men_n219_), .C(men_men_n441_), .D(men_men_n434_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n918_), .B(i_11_), .Y(men_men_n919_));
  AN2        u0897(.A(men_men_n99_), .B(men_men_n248_), .Y(men_men_n920_));
  NA2        u0898(.A(men_men_n793_), .B(men_men_n340_), .Y(men_men_n921_));
  AOI210     u0899(.A0(men_men_n516_), .A1(men_men_n89_), .B0(men_men_n58_), .Y(men_men_n922_));
  OAI220     u0900(.A0(men_men_n922_), .A1(men_men_n921_), .B0(men_men_n709_), .B1(men_men_n578_), .Y(men_men_n923_));
  NO2        u0901(.A(men_men_n259_), .B(men_men_n154_), .Y(men_men_n924_));
  NA2        u0902(.A(i_0_), .B(i_10_), .Y(men_men_n925_));
  OAI210     u0903(.A0(men_men_n925_), .A1(men_men_n86_), .B0(men_men_n581_), .Y(men_men_n926_));
  NO4        u0904(.A(men_men_n114_), .B(men_men_n58_), .C(men_men_n717_), .D(i_5_), .Y(men_men_n927_));
  AO220      u0905(.A0(men_men_n927_), .A1(men_men_n926_), .B0(men_men_n924_), .B1(i_6_), .Y(men_men_n928_));
  AOI220     u0906(.A0(men_men_n346_), .A1(men_men_n101_), .B0(men_men_n188_), .B1(men_men_n84_), .Y(men_men_n929_));
  NA2        u0907(.A(men_men_n612_), .B(i_4_), .Y(men_men_n930_));
  NA2        u0908(.A(men_men_n191_), .B(men_men_n205_), .Y(men_men_n931_));
  OAI220     u0909(.A0(men_men_n931_), .A1(men_men_n921_), .B0(men_men_n930_), .B1(men_men_n929_), .Y(men_men_n932_));
  NO4        u0910(.A(men_men_n932_), .B(men_men_n928_), .C(men_men_n923_), .D(men_men_n920_), .Y(men_men_n933_));
  NA4        u0911(.A(men_men_n933_), .B(men_men_n919_), .C(men_men_n917_), .D(men_men_n915_), .Y(men_men_n934_));
  NO2        u0912(.A(men_men_n106_), .B(men_men_n37_), .Y(men_men_n935_));
  NA2        u0913(.A(i_11_), .B(i_9_), .Y(men_men_n936_));
  NO3        u0914(.A(i_12_), .B(men_men_n936_), .C(men_men_n651_), .Y(men_men_n937_));
  AO220      u0915(.A0(men_men_n937_), .A1(men_men_n935_), .B0(men_men_n277_), .B1(men_men_n88_), .Y(men_men_n938_));
  NO2        u0916(.A(men_men_n48_), .B(i_7_), .Y(men_men_n939_));
  NAi31      u0917(.An(men_men_n272_), .B(men_men_n489_), .C(men_men_n161_), .Y(men_men_n940_));
  NO2        u0918(.A(men_men_n936_), .B(men_men_n73_), .Y(men_men_n941_));
  NO2        u0919(.A(men_men_n177_), .B(i_0_), .Y(men_men_n942_));
  INV        u0920(.A(men_men_n942_), .Y(men_men_n943_));
  NA2        u0921(.A(men_men_n505_), .B(men_men_n235_), .Y(men_men_n944_));
  AOI210     u0922(.A0(men_men_n390_), .A1(men_men_n41_), .B0(men_men_n432_), .Y(men_men_n945_));
  OAI220     u0923(.A0(men_men_n945_), .A1(men_men_n902_), .B0(men_men_n944_), .B1(men_men_n943_), .Y(men_men_n946_));
  NO3        u0924(.A(men_men_n946_), .B(men_men_n940_), .C(men_men_n938_), .Y(men_men_n947_));
  AOI210     u0925(.A0(men_men_n475_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n948_));
  NA2        u0926(.A(men_men_n173_), .B(men_men_n106_), .Y(men_men_n949_));
  NOi32      u0927(.An(men_men_n948_), .Bn(men_men_n191_), .C(men_men_n949_), .Y(men_men_n950_));
  AOI210     u0928(.A0(men_men_n653_), .A1(men_men_n340_), .B0(men_men_n248_), .Y(men_men_n951_));
  NO2        u0929(.A(men_men_n951_), .B(men_men_n891_), .Y(men_men_n952_));
  NO2        u0930(.A(men_men_n952_), .B(men_men_n950_), .Y(men_men_n953_));
  NOi21      u0931(.An(i_7_), .B(i_5_), .Y(men_men_n954_));
  NOi31      u0932(.An(men_men_n954_), .B(i_0_), .C(men_men_n774_), .Y(men_men_n955_));
  NA3        u0933(.A(men_men_n955_), .B(men_men_n404_), .C(i_6_), .Y(men_men_n956_));
  OA210      u0934(.A0(men_men_n949_), .A1(men_men_n553_), .B0(men_men_n956_), .Y(men_men_n957_));
  NO3        u0935(.A(men_men_n427_), .B(men_men_n379_), .C(men_men_n375_), .Y(men_men_n958_));
  NO2        u0936(.A(men_men_n269_), .B(men_men_n329_), .Y(men_men_n959_));
  NO2        u0937(.A(men_men_n774_), .B(men_men_n264_), .Y(men_men_n960_));
  AOI210     u0938(.A0(men_men_n960_), .A1(men_men_n959_), .B0(men_men_n958_), .Y(men_men_n961_));
  NA4        u0939(.A(men_men_n961_), .B(men_men_n957_), .C(men_men_n953_), .D(men_men_n947_), .Y(men_men_n962_));
  NO2        u0940(.A(men_men_n909_), .B(men_men_n244_), .Y(men_men_n963_));
  AN2        u0941(.A(men_men_n345_), .B(men_men_n340_), .Y(men_men_n964_));
  AO220      u0942(.A0(men_men_n964_), .A1(men_men_n905_), .B0(men_men_n361_), .B1(men_men_n27_), .Y(men_men_n965_));
  OAI210     u0943(.A0(men_men_n965_), .A1(men_men_n963_), .B0(i_10_), .Y(men_men_n966_));
  NO2        u0944(.A(men_men_n879_), .B(men_men_n328_), .Y(men_men_n967_));
  OA210      u0945(.A0(men_men_n505_), .A1(men_men_n228_), .B0(men_men_n504_), .Y(men_men_n968_));
  NA2        u0946(.A(men_men_n967_), .B(men_men_n941_), .Y(men_men_n969_));
  NA3        u0947(.A(men_men_n504_), .B(men_men_n435_), .C(men_men_n45_), .Y(men_men_n970_));
  OAI210     u0948(.A0(men_men_n913_), .A1(i_7_), .B0(men_men_n970_), .Y(men_men_n971_));
  NO2        u0949(.A(men_men_n262_), .B(men_men_n46_), .Y(men_men_n972_));
  NA2        u0950(.A(men_men_n941_), .B(men_men_n315_), .Y(men_men_n973_));
  OAI210     u0951(.A0(men_men_n972_), .A1(men_men_n190_), .B0(men_men_n973_), .Y(men_men_n974_));
  AOI220     u0952(.A0(men_men_n974_), .A1(men_men_n505_), .B0(men_men_n971_), .B1(men_men_n73_), .Y(men_men_n975_));
  NA3        u0953(.A(men_men_n854_), .B(men_men_n402_), .C(men_men_n688_), .Y(men_men_n976_));
  NA2        u0954(.A(men_men_n95_), .B(men_men_n44_), .Y(men_men_n977_));
  NO2        u0955(.A(men_men_n75_), .B(men_men_n795_), .Y(men_men_n978_));
  AOI220     u0956(.A0(men_men_n978_), .A1(men_men_n977_), .B0(men_men_n176_), .B1(men_men_n643_), .Y(men_men_n979_));
  AOI210     u0957(.A0(men_men_n979_), .A1(men_men_n976_), .B0(men_men_n47_), .Y(men_men_n980_));
  NO3        u0958(.A(men_men_n635_), .B(men_men_n374_), .C(men_men_n24_), .Y(men_men_n981_));
  AOI210     u0959(.A0(men_men_n750_), .A1(men_men_n590_), .B0(men_men_n981_), .Y(men_men_n982_));
  NAi21      u0960(.An(i_9_), .B(i_5_), .Y(men_men_n983_));
  NO2        u0961(.A(men_men_n983_), .B(men_men_n427_), .Y(men_men_n984_));
  NO2        u0962(.A(men_men_n647_), .B(men_men_n108_), .Y(men_men_n985_));
  AOI220     u0963(.A0(men_men_n985_), .A1(i_0_), .B0(men_men_n984_), .B1(men_men_n669_), .Y(men_men_n986_));
  OAI220     u0964(.A0(men_men_n986_), .A1(men_men_n86_), .B0(men_men_n982_), .B1(men_men_n174_), .Y(men_men_n987_));
  NO3        u0965(.A(men_men_n987_), .B(men_men_n980_), .C(men_men_n558_), .Y(men_men_n988_));
  NA4        u0966(.A(men_men_n988_), .B(men_men_n975_), .C(men_men_n969_), .D(men_men_n966_), .Y(men_men_n989_));
  NO3        u0967(.A(men_men_n989_), .B(men_men_n962_), .C(men_men_n934_), .Y(men_men_n990_));
  NO2        u0968(.A(i_0_), .B(men_men_n774_), .Y(men_men_n991_));
  NA2        u0969(.A(men_men_n73_), .B(men_men_n44_), .Y(men_men_n992_));
  NO3        u0970(.A(men_men_n108_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n993_));
  AO220      u0971(.A0(men_men_n993_), .A1(men_men_n73_), .B0(men_men_n991_), .B1(men_men_n176_), .Y(men_men_n994_));
  NO2        u0972(.A(men_men_n737_), .B(men_men_n949_), .Y(men_men_n995_));
  AOI210     u0973(.A0(men_men_n994_), .A1(men_men_n363_), .B0(men_men_n995_), .Y(men_men_n996_));
  NA2        u0974(.A(men_men_n783_), .B(men_men_n146_), .Y(men_men_n997_));
  INV        u0975(.A(men_men_n997_), .Y(men_men_n998_));
  NA3        u0976(.A(men_men_n998_), .B(men_men_n724_), .C(men_men_n73_), .Y(men_men_n999_));
  NO2        u0977(.A(men_men_n850_), .B(men_men_n427_), .Y(men_men_n1000_));
  NA3        u0978(.A(men_men_n881_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n1001_));
  NA2        u0979(.A(men_men_n882_), .B(i_9_), .Y(men_men_n1002_));
  AOI210     u0980(.A0(men_men_n1001_), .A1(men_men_n532_), .B0(men_men_n1002_), .Y(men_men_n1003_));
  NO2        u0981(.A(men_men_n1003_), .B(men_men_n1000_), .Y(men_men_n1004_));
  NA3        u0982(.A(men_men_n1004_), .B(men_men_n999_), .C(men_men_n996_), .Y(men_men_n1005_));
  NA2        u0983(.A(men_men_n964_), .B(men_men_n392_), .Y(men_men_n1006_));
  AOI210     u0984(.A0(men_men_n310_), .A1(men_men_n163_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  NA2        u0985(.A(men_men_n939_), .B(men_men_n521_), .Y(men_men_n1008_));
  AOI210     u0986(.A0(i_11_), .A1(men_men_n163_), .B0(men_men_n1008_), .Y(men_men_n1009_));
  NO2        u0987(.A(men_men_n1009_), .B(men_men_n1007_), .Y(men_men_n1010_));
  NO3        u0988(.A(men_men_n925_), .B(men_men_n901_), .C(men_men_n192_), .Y(men_men_n1011_));
  AOI220     u0989(.A0(men_men_n1011_), .A1(i_11_), .B0(men_men_n613_), .B1(men_men_n75_), .Y(men_men_n1012_));
  NO3        u0990(.A(men_men_n213_), .B(men_men_n403_), .C(i_0_), .Y(men_men_n1013_));
  OAI210     u0991(.A0(men_men_n1013_), .A1(men_men_n76_), .B0(i_13_), .Y(men_men_n1014_));
  INV        u0992(.A(men_men_n222_), .Y(men_men_n1015_));
  OAI220     u0993(.A0(men_men_n571_), .A1(men_men_n139_), .B0(men_men_n693_), .B1(men_men_n664_), .Y(men_men_n1016_));
  NA3        u0994(.A(men_men_n1016_), .B(men_men_n419_), .C(men_men_n1015_), .Y(men_men_n1017_));
  NA4        u0995(.A(men_men_n1017_), .B(men_men_n1014_), .C(men_men_n1012_), .D(men_men_n1010_), .Y(men_men_n1018_));
  NO2        u0996(.A(men_men_n247_), .B(men_men_n95_), .Y(men_men_n1019_));
  AOI210     u0997(.A0(men_men_n1019_), .A1(men_men_n991_), .B0(men_men_n110_), .Y(men_men_n1020_));
  AOI220     u0998(.A0(men_men_n954_), .A1(men_men_n521_), .B0(men_men_n881_), .B1(men_men_n164_), .Y(men_men_n1021_));
  NA2        u0999(.A(men_men_n366_), .B(men_men_n178_), .Y(men_men_n1022_));
  OA220      u1000(.A0(men_men_n1022_), .A1(men_men_n1021_), .B0(men_men_n1020_), .B1(i_5_), .Y(men_men_n1023_));
  AOI210     u1001(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n177_), .Y(men_men_n1024_));
  NA2        u1002(.A(men_men_n1024_), .B(men_men_n968_), .Y(men_men_n1025_));
  NA3        u1003(.A(men_men_n661_), .B(men_men_n188_), .C(men_men_n84_), .Y(men_men_n1026_));
  NA2        u1004(.A(men_men_n1026_), .B(men_men_n588_), .Y(men_men_n1027_));
  NO3        u1005(.A(men_men_n891_), .B(men_men_n54_), .C(men_men_n48_), .Y(men_men_n1028_));
  NA2        u1006(.A(men_men_n526_), .B(men_men_n519_), .Y(men_men_n1029_));
  NO3        u1007(.A(men_men_n1029_), .B(men_men_n1028_), .C(men_men_n1027_), .Y(men_men_n1030_));
  NA3        u1008(.A(men_men_n410_), .B(men_men_n173_), .C(men_men_n172_), .Y(men_men_n1031_));
  NA3        u1009(.A(men_men_n939_), .B(men_men_n299_), .C(i_10_), .Y(men_men_n1032_));
  NA2        u1010(.A(men_men_n1032_), .B(men_men_n1031_), .Y(men_men_n1033_));
  NA3        u1011(.A(men_men_n410_), .B(men_men_n347_), .C(men_men_n226_), .Y(men_men_n1034_));
  INV        u1012(.A(men_men_n1034_), .Y(men_men_n1035_));
  NOi31      u1013(.An(men_men_n409_), .B(men_men_n992_), .C(men_men_n244_), .Y(men_men_n1036_));
  NO3        u1014(.A(men_men_n936_), .B(men_men_n222_), .C(men_men_n192_), .Y(men_men_n1037_));
  NO4        u1015(.A(men_men_n1037_), .B(men_men_n1036_), .C(men_men_n1035_), .D(men_men_n1033_), .Y(men_men_n1038_));
  NA4        u1016(.A(men_men_n1038_), .B(men_men_n1030_), .C(men_men_n1025_), .D(men_men_n1023_), .Y(men_men_n1039_));
  AOI210     u1017(.A0(men_men_n612_), .A1(men_men_n570_), .B0(men_men_n663_), .Y(men_men_n1040_));
  NO3        u1018(.A(men_men_n1040_), .B(men_men_n603_), .C(men_men_n360_), .Y(men_men_n1041_));
  NA3        u1019(.A(men_men_n882_), .B(men_men_n111_), .C(men_men_n124_), .Y(men_men_n1042_));
  INV        u1020(.A(men_men_n1042_), .Y(men_men_n1043_));
  AOI210     u1021(.A0(men_men_n1043_), .A1(men_men_n1114_), .B0(men_men_n1041_), .Y(men_men_n1044_));
  NA3        u1022(.A(men_men_n315_), .B(i_5_), .C(men_men_n195_), .Y(men_men_n1045_));
  NAi31      u1023(.An(men_men_n246_), .B(men_men_n1045_), .C(men_men_n247_), .Y(men_men_n1046_));
  NO4        u1024(.A(men_men_n244_), .B(men_men_n213_), .C(i_0_), .D(i_12_), .Y(men_men_n1047_));
  AOI220     u1025(.A0(men_men_n1047_), .A1(men_men_n1046_), .B0(men_men_n832_), .B1(men_men_n178_), .Y(men_men_n1048_));
  AN2        u1026(.A(men_men_n925_), .B(men_men_n154_), .Y(men_men_n1049_));
  NO4        u1027(.A(men_men_n1049_), .B(i_12_), .C(men_men_n697_), .D(men_men_n131_), .Y(men_men_n1050_));
  NA2        u1028(.A(men_men_n1050_), .B(men_men_n222_), .Y(men_men_n1051_));
  NA3        u1029(.A(men_men_n101_), .B(men_men_n617_), .C(i_11_), .Y(men_men_n1052_));
  NO2        u1030(.A(men_men_n1052_), .B(men_men_n156_), .Y(men_men_n1053_));
  NA2        u1031(.A(men_men_n954_), .B(men_men_n502_), .Y(men_men_n1054_));
  OAI220     u1032(.A0(i_7_), .A1(men_men_n1045_), .B0(men_men_n1054_), .B1(men_men_n725_), .Y(men_men_n1055_));
  AOI210     u1033(.A0(men_men_n1055_), .A1(men_men_n942_), .B0(men_men_n1053_), .Y(men_men_n1056_));
  NA4        u1034(.A(men_men_n1056_), .B(men_men_n1051_), .C(men_men_n1048_), .D(men_men_n1044_), .Y(men_men_n1057_));
  NO4        u1035(.A(men_men_n1057_), .B(men_men_n1039_), .C(men_men_n1018_), .D(men_men_n1005_), .Y(men_men_n1058_));
  OAI210     u1036(.A0(men_men_n853_), .A1(men_men_n847_), .B0(men_men_n37_), .Y(men_men_n1059_));
  NA3        u1037(.A(men_men_n948_), .B(men_men_n387_), .C(i_5_), .Y(men_men_n1060_));
  NA3        u1038(.A(men_men_n1060_), .B(men_men_n1059_), .C(men_men_n659_), .Y(men_men_n1061_));
  NA2        u1039(.A(men_men_n1061_), .B(men_men_n210_), .Y(men_men_n1062_));
  AN2        u1040(.A(men_men_n746_), .B(men_men_n388_), .Y(men_men_n1063_));
  NA2        u1041(.A(men_men_n189_), .B(men_men_n191_), .Y(men_men_n1064_));
  AO210      u1042(.A0(men_men_n1063_), .A1(men_men_n33_), .B0(men_men_n1064_), .Y(men_men_n1065_));
  OAI210     u1043(.A0(men_men_n663_), .A1(men_men_n661_), .B0(men_men_n328_), .Y(men_men_n1066_));
  NAi31      u1044(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1067_));
  NO2        u1045(.A(men_men_n70_), .B(men_men_n1067_), .Y(men_men_n1068_));
  NO2        u1046(.A(men_men_n1068_), .B(men_men_n694_), .Y(men_men_n1069_));
  NA3        u1047(.A(men_men_n1069_), .B(men_men_n1066_), .C(men_men_n1065_), .Y(men_men_n1070_));
  NO2        u1048(.A(men_men_n492_), .B(men_men_n275_), .Y(men_men_n1071_));
  NO4        u1049(.A(men_men_n237_), .B(men_men_n145_), .C(men_men_n728_), .D(men_men_n37_), .Y(men_men_n1072_));
  NO3        u1050(.A(men_men_n1072_), .B(men_men_n1071_), .C(men_men_n918_), .Y(men_men_n1073_));
  OAI210     u1051(.A0(men_men_n1052_), .A1(men_men_n148_), .B0(men_men_n1073_), .Y(men_men_n1074_));
  AOI210     u1052(.A0(men_men_n1070_), .A1(men_men_n48_), .B0(men_men_n1074_), .Y(men_men_n1075_));
  AOI210     u1053(.A0(men_men_n1075_), .A1(men_men_n1062_), .B0(men_men_n73_), .Y(men_men_n1076_));
  NO2        u1054(.A(men_men_n610_), .B(men_men_n399_), .Y(men_men_n1077_));
  NO2        u1055(.A(men_men_n1077_), .B(men_men_n800_), .Y(men_men_n1078_));
  OAI210     u1056(.A0(men_men_n80_), .A1(men_men_n54_), .B0(men_men_n109_), .Y(men_men_n1079_));
  NA2        u1057(.A(men_men_n1079_), .B(men_men_n76_), .Y(men_men_n1080_));
  AOI210     u1058(.A0(men_men_n1024_), .A1(men_men_n939_), .B0(men_men_n955_), .Y(men_men_n1081_));
  AOI210     u1059(.A0(men_men_n1081_), .A1(men_men_n1080_), .B0(men_men_n728_), .Y(men_men_n1082_));
  NA2        u1060(.A(men_men_n269_), .B(men_men_n57_), .Y(men_men_n1083_));
  AOI220     u1061(.A0(men_men_n1083_), .A1(men_men_n76_), .B0(men_men_n361_), .B1(men_men_n261_), .Y(men_men_n1084_));
  NO2        u1062(.A(men_men_n1084_), .B(men_men_n241_), .Y(men_men_n1085_));
  NA3        u1063(.A(men_men_n99_), .B(men_men_n317_), .C(men_men_n31_), .Y(men_men_n1086_));
  INV        u1064(.A(men_men_n1086_), .Y(men_men_n1087_));
  NO3        u1065(.A(men_men_n1087_), .B(men_men_n1085_), .C(men_men_n1082_), .Y(men_men_n1088_));
  OAI210     u1066(.A0(men_men_n277_), .A1(men_men_n159_), .B0(men_men_n89_), .Y(men_men_n1089_));
  NA3        u1067(.A(men_men_n804_), .B(men_men_n299_), .C(men_men_n80_), .Y(men_men_n1090_));
  AOI210     u1068(.A0(men_men_n1090_), .A1(men_men_n1089_), .B0(i_11_), .Y(men_men_n1091_));
  NA2        u1069(.A(men_men_n654_), .B(men_men_n219_), .Y(men_men_n1092_));
  OAI210     u1070(.A0(men_men_n1092_), .A1(men_men_n948_), .B0(men_men_n210_), .Y(men_men_n1093_));
  NA2        u1071(.A(men_men_n165_), .B(i_5_), .Y(men_men_n1094_));
  AOI210     u1072(.A0(men_men_n1093_), .A1(men_men_n813_), .B0(men_men_n1094_), .Y(men_men_n1095_));
  NO3        u1073(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1096_));
  OAI210     u1074(.A0(men_men_n959_), .A1(men_men_n317_), .B0(men_men_n1096_), .Y(men_men_n1097_));
  NO2        u1075(.A(men_men_n1097_), .B(men_men_n774_), .Y(men_men_n1098_));
  NO4        u1076(.A(men_men_n983_), .B(men_men_n509_), .C(men_men_n258_), .D(men_men_n257_), .Y(men_men_n1099_));
  NO2        u1077(.A(men_men_n1099_), .B(men_men_n607_), .Y(men_men_n1100_));
  NO2        u1078(.A(men_men_n849_), .B(men_men_n380_), .Y(men_men_n1101_));
  AOI210     u1079(.A0(men_men_n1101_), .A1(men_men_n1100_), .B0(men_men_n40_), .Y(men_men_n1102_));
  NO4        u1080(.A(men_men_n1102_), .B(men_men_n1098_), .C(men_men_n1095_), .D(men_men_n1091_), .Y(men_men_n1103_));
  OAI210     u1081(.A0(men_men_n1088_), .A1(i_4_), .B0(men_men_n1103_), .Y(men_men_n1104_));
  NO3        u1082(.A(men_men_n1104_), .B(men_men_n1078_), .C(men_men_n1076_), .Y(men_men_n1105_));
  NA4        u1083(.A(men_men_n1105_), .B(men_men_n1058_), .C(men_men_n990_), .D(men_men_n908_), .Y(men4));
  INV        u1084(.A(i_5_), .Y(men_men_n1109_));
  INV        u1085(.A(men_men_n383_), .Y(men_men_n1110_));
  INV        u1086(.A(men_men_n144_), .Y(men_men_n1111_));
  INV        u1087(.A(i_1_), .Y(men_men_n1112_));
  INV        u1088(.A(i_9_), .Y(men_men_n1113_));
  INV        u1089(.A(i_5_), .Y(men_men_n1114_));
  INV        u1090(.A(i_7_), .Y(men_men_n1115_));
  INV        u1091(.A(i_3_), .Y(men_men_n1116_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule