// Benchmark "top" written by ABC on Fri Jun 21 17:49:24 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n129_, new_new_n130_, new_new_n131_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n674_,
    new_new_n675_, new_new_n676_, new_new_n677_, new_new_n678_,
    new_new_n679_, new_new_n680_, new_new_n681_, new_new_n682_,
    new_new_n683_, new_new_n684_, new_new_n685_, new_new_n686_,
    new_new_n687_, new_new_n688_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n722_, new_new_n723_,
    new_new_n724_, new_new_n725_, new_new_n726_, new_new_n727_,
    new_new_n728_, new_new_n729_, new_new_n730_, new_new_n731_,
    new_new_n732_, new_new_n733_, new_new_n734_, new_new_n735_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n964_, new_new_n965_, new_new_n966_, new_new_n967_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NO2        g028(.A(new_new_n47_), .B(new_new_n46_), .Y(new_new_n51_));
  NA2        g029(.A(i_0_), .B(i_2_), .Y(new_new_n52_));
  NA2        g030(.A(i_7_), .B(i_9_), .Y(new_new_n53_));
  NA2        g031(.A(new_new_n51_), .B(new_new_n45_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  NAi21      g034(.An(i_2_), .B(i_7_), .Y(new_new_n57_));
  INV        g035(.A(i_1_), .Y(new_new_n58_));
  NA2        g036(.A(i_1_), .B(i_10_), .Y(new_new_n59_));
  NO2        g037(.A(new_new_n59_), .B(i_6_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n50_), .B(i_2_), .Y(new_new_n61_));
  AOI210     g039(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_6_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(new_new_n25_), .Y(new_new_n64_));
  INV        g042(.A(i_0_), .Y(new_new_n65_));
  NAi21      g043(.An(i_5_), .B(i_10_), .Y(new_new_n66_));
  NA2        g044(.A(i_5_), .B(i_9_), .Y(new_new_n67_));
  AOI210     g045(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n65_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n64_), .Y(new_new_n69_));
  OAI210     g047(.A0(new_new_n62_), .A1(new_new_n61_), .B0(new_new_n69_), .Y(new_new_n70_));
  OAI210     g048(.A0(new_new_n70_), .A1(new_new_n60_), .B0(i_0_), .Y(new_new_n71_));
  NA2        g049(.A(i_12_), .B(i_5_), .Y(new_new_n72_));
  NO2        g050(.A(i_3_), .B(i_9_), .Y(new_new_n73_));
  NO2        g051(.A(i_3_), .B(i_7_), .Y(new_new_n74_));
  NO3        g052(.A(new_new_n74_), .B(new_new_n73_), .C(new_new_n58_), .Y(new_new_n75_));
  INV        g053(.A(i_6_), .Y(new_new_n76_));
  OR4        g054(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n77_));
  INV        g055(.A(new_new_n77_), .Y(new_new_n78_));
  NO2        g056(.A(i_2_), .B(i_7_), .Y(new_new_n79_));
  NO2        g057(.A(new_new_n78_), .B(new_new_n79_), .Y(new_new_n80_));
  NA2        g058(.A(new_new_n75_), .B(new_new_n80_), .Y(new_new_n81_));
  NAi21      g059(.An(i_6_), .B(i_10_), .Y(new_new_n82_));
  NA2        g060(.A(i_6_), .B(i_9_), .Y(new_new_n83_));
  AOI210     g061(.A0(new_new_n83_), .A1(new_new_n82_), .B0(new_new_n58_), .Y(new_new_n84_));
  NA2        g062(.A(i_2_), .B(i_6_), .Y(new_new_n85_));
  INV        g063(.A(new_new_n84_), .Y(new_new_n86_));
  AOI210     g064(.A0(new_new_n86_), .A1(new_new_n81_), .B0(new_new_n72_), .Y(new_new_n87_));
  AN3        g065(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_11_), .Y(new_new_n89_));
  NO2        g067(.A(i_5_), .B(i_8_), .Y(new_new_n90_));
  NOi21      g068(.An(new_new_n90_), .B(new_new_n89_), .Y(new_new_n91_));
  AOI220     g069(.A0(new_new_n91_), .A1(new_new_n57_), .B0(new_new_n88_), .B1(new_new_n32_), .Y(new_new_n92_));
  INV        g070(.A(i_7_), .Y(new_new_n93_));
  NA2        g071(.A(new_new_n46_), .B(new_new_n93_), .Y(new_new_n94_));
  NO2        g072(.A(i_0_), .B(i_5_), .Y(new_new_n95_));
  NO2        g073(.A(new_new_n95_), .B(new_new_n76_), .Y(new_new_n96_));
  NA2        g074(.A(i_12_), .B(i_3_), .Y(new_new_n97_));
  INV        g075(.A(new_new_n97_), .Y(new_new_n98_));
  NA3        g076(.A(new_new_n98_), .B(new_new_n96_), .C(new_new_n94_), .Y(new_new_n99_));
  NAi21      g077(.An(i_7_), .B(i_11_), .Y(new_new_n100_));
  AN2        g078(.A(i_2_), .B(i_10_), .Y(new_new_n101_));
  NO2        g079(.A(new_new_n101_), .B(i_7_), .Y(new_new_n102_));
  OR2        g080(.A(new_new_n72_), .B(new_new_n55_), .Y(new_new_n103_));
  NO2        g081(.A(i_8_), .B(new_new_n93_), .Y(new_new_n104_));
  NO3        g082(.A(new_new_n104_), .B(new_new_n103_), .C(new_new_n102_), .Y(new_new_n105_));
  NA2        g083(.A(i_12_), .B(i_7_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n58_), .B(new_new_n26_), .Y(new_new_n107_));
  NA2        g085(.A(new_new_n107_), .B(i_0_), .Y(new_new_n108_));
  NA2        g086(.A(i_11_), .B(i_12_), .Y(new_new_n109_));
  OAI210     g087(.A0(new_new_n108_), .A1(new_new_n106_), .B0(new_new_n109_), .Y(new_new_n110_));
  NO2        g088(.A(new_new_n110_), .B(new_new_n105_), .Y(new_new_n111_));
  NA3        g089(.A(new_new_n111_), .B(new_new_n99_), .C(new_new_n92_), .Y(new_new_n112_));
  NOi21      g090(.An(i_1_), .B(i_5_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n113_), .B(i_11_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n93_), .B(new_new_n37_), .Y(new_new_n115_));
  NA2        g093(.A(i_7_), .B(new_new_n25_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(new_new_n115_), .Y(new_new_n117_));
  NO2        g095(.A(new_new_n117_), .B(new_new_n46_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n83_), .B(new_new_n82_), .Y(new_new_n119_));
  NAi21      g097(.An(i_3_), .B(i_8_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(new_new_n57_), .Y(new_new_n121_));
  NOi31      g099(.An(new_new_n121_), .B(new_new_n119_), .C(new_new_n118_), .Y(new_new_n122_));
  NO2        g100(.A(i_1_), .B(new_new_n76_), .Y(new_new_n123_));
  NO2        g101(.A(i_6_), .B(i_5_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(i_3_), .Y(new_new_n125_));
  OAI220     g103(.A0(new_new_n125_), .A1(new_new_n100_), .B0(new_new_n122_), .B1(new_new_n114_), .Y(new_new_n126_));
  NO3        g104(.A(new_new_n126_), .B(new_new_n112_), .C(new_new_n87_), .Y(new_new_n127_));
  NA3        g105(.A(new_new_n127_), .B(new_new_n71_), .C(new_new_n54_), .Y(mai2));
  NO2        g106(.A(new_new_n58_), .B(new_new_n37_), .Y(new_new_n129_));
  NA2        g107(.A(i_6_), .B(new_new_n25_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(new_new_n129_), .Y(new_new_n131_));
  NA4        g109(.A(new_new_n131_), .B(new_new_n69_), .C(new_new_n61_), .D(new_new_n30_), .Y(mai0));
  AN2        g110(.A(i_8_), .B(i_7_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n133_), .B(i_6_), .Y(new_new_n134_));
  NO2        g112(.A(i_12_), .B(i_13_), .Y(new_new_n135_));
  NAi21      g113(.An(i_5_), .B(i_11_), .Y(new_new_n136_));
  NOi21      g114(.An(new_new_n135_), .B(new_new_n136_), .Y(new_new_n137_));
  NO2        g115(.A(i_0_), .B(i_1_), .Y(new_new_n138_));
  NA2        g116(.A(i_2_), .B(i_3_), .Y(new_new_n139_));
  NO2        g117(.A(new_new_n139_), .B(i_4_), .Y(new_new_n140_));
  NA3        g118(.A(new_new_n140_), .B(new_new_n138_), .C(new_new_n137_), .Y(new_new_n141_));
  AN2        g119(.A(new_new_n135_), .B(new_new_n73_), .Y(new_new_n142_));
  NA2        g120(.A(i_1_), .B(i_5_), .Y(new_new_n143_));
  NO2        g121(.A(new_new_n65_), .B(new_new_n46_), .Y(new_new_n144_));
  NA2        g122(.A(new_new_n144_), .B(new_new_n36_), .Y(new_new_n145_));
  NO3        g123(.A(new_new_n145_), .B(new_new_n143_), .C(i_13_), .Y(new_new_n146_));
  OR2        g124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NO3        g125(.A(new_new_n147_), .B(new_new_n72_), .C(i_13_), .Y(new_new_n148_));
  NAi32      g126(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n149_));
  NAi21      g127(.An(new_new_n149_), .B(new_new_n148_), .Y(new_new_n150_));
  NOi21      g128(.An(i_4_), .B(i_10_), .Y(new_new_n151_));
  NA2        g129(.A(new_new_n151_), .B(new_new_n40_), .Y(new_new_n152_));
  NO2        g130(.A(i_3_), .B(i_5_), .Y(new_new_n153_));
  NO3        g131(.A(new_new_n65_), .B(i_2_), .C(i_1_), .Y(new_new_n154_));
  NA2        g132(.A(new_new_n154_), .B(new_new_n153_), .Y(new_new_n155_));
  OAI210     g133(.A0(new_new_n155_), .A1(new_new_n152_), .B0(new_new_n150_), .Y(new_new_n156_));
  NO2        g134(.A(new_new_n156_), .B(new_new_n146_), .Y(new_new_n157_));
  AOI210     g135(.A0(new_new_n157_), .A1(new_new_n141_), .B0(new_new_n134_), .Y(new_new_n158_));
  NA2        g136(.A(i_3_), .B(new_new_n48_), .Y(new_new_n159_));
  NOi21      g137(.An(i_4_), .B(i_9_), .Y(new_new_n160_));
  NOi21      g138(.An(i_11_), .B(i_13_), .Y(new_new_n161_));
  NA2        g139(.A(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  OR2        g140(.A(new_new_n162_), .B(new_new_n159_), .Y(new_new_n163_));
  NO2        g141(.A(i_4_), .B(i_5_), .Y(new_new_n164_));
  NAi21      g142(.An(i_12_), .B(i_11_), .Y(new_new_n165_));
  NO2        g143(.A(new_new_n165_), .B(i_13_), .Y(new_new_n166_));
  NA3        g144(.A(new_new_n166_), .B(new_new_n164_), .C(new_new_n73_), .Y(new_new_n167_));
  NA2        g145(.A(new_new_n167_), .B(new_new_n163_), .Y(new_new_n168_));
  NO2        g146(.A(new_new_n65_), .B(new_new_n58_), .Y(new_new_n169_));
  NA2        g147(.A(new_new_n169_), .B(new_new_n46_), .Y(new_new_n170_));
  NAi31      g148(.An(new_new_n965_), .B(new_new_n142_), .C(i_11_), .Y(new_new_n171_));
  NA2        g149(.A(i_3_), .B(i_5_), .Y(new_new_n172_));
  AOI210     g150(.A0(new_new_n162_), .A1(new_new_n171_), .B0(new_new_n170_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n65_), .B(i_5_), .Y(new_new_n174_));
  NO2        g152(.A(i_13_), .B(i_10_), .Y(new_new_n175_));
  NA3        g153(.A(new_new_n175_), .B(new_new_n174_), .C(new_new_n44_), .Y(new_new_n176_));
  NO2        g154(.A(i_2_), .B(i_1_), .Y(new_new_n177_));
  NA2        g155(.A(new_new_n177_), .B(i_3_), .Y(new_new_n178_));
  NAi21      g156(.An(i_4_), .B(i_12_), .Y(new_new_n179_));
  NO3        g157(.A(new_new_n179_), .B(new_new_n178_), .C(new_new_n176_), .Y(new_new_n180_));
  NO3        g158(.A(new_new_n180_), .B(new_new_n173_), .C(new_new_n168_), .Y(new_new_n181_));
  INV        g159(.A(i_8_), .Y(new_new_n182_));
  NO2        g160(.A(new_new_n182_), .B(i_7_), .Y(new_new_n183_));
  NA2        g161(.A(new_new_n183_), .B(i_6_), .Y(new_new_n184_));
  NO3        g162(.A(i_3_), .B(new_new_n76_), .C(new_new_n48_), .Y(new_new_n185_));
  NA2        g163(.A(new_new_n185_), .B(new_new_n104_), .Y(new_new_n186_));
  NO3        g164(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n187_));
  NA3        g165(.A(new_new_n187_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n188_));
  NO3        g166(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n189_));
  INV        g167(.A(new_new_n189_), .Y(new_new_n190_));
  AOI210     g168(.A0(new_new_n190_), .A1(new_new_n188_), .B0(new_new_n186_), .Y(new_new_n191_));
  NO2        g169(.A(i_3_), .B(i_8_), .Y(new_new_n192_));
  NO3        g170(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n193_));
  NA3        g171(.A(new_new_n193_), .B(new_new_n192_), .C(new_new_n40_), .Y(new_new_n194_));
  NO2        g172(.A(new_new_n95_), .B(new_new_n55_), .Y(new_new_n195_));
  NO2        g173(.A(i_13_), .B(i_9_), .Y(new_new_n196_));
  NA3        g174(.A(new_new_n196_), .B(i_6_), .C(new_new_n182_), .Y(new_new_n197_));
  BUFFER     g175(.A(new_new_n197_), .Y(new_new_n198_));
  NO2        g176(.A(new_new_n44_), .B(i_5_), .Y(new_new_n199_));
  NO3        g177(.A(i_0_), .B(i_2_), .C(new_new_n58_), .Y(new_new_n200_));
  NA3        g178(.A(new_new_n200_), .B(new_new_n199_), .C(i_10_), .Y(new_new_n201_));
  OAI210     g179(.A0(new_new_n201_), .A1(new_new_n198_), .B0(new_new_n194_), .Y(new_new_n202_));
  AOI210     g180(.A0(new_new_n202_), .A1(i_7_), .B0(new_new_n191_), .Y(new_new_n203_));
  OAI220     g181(.A0(new_new_n203_), .A1(i_4_), .B0(new_new_n184_), .B1(new_new_n181_), .Y(new_new_n204_));
  NA3        g182(.A(i_13_), .B(new_new_n182_), .C(i_10_), .Y(new_new_n205_));
  NO2        g183(.A(new_new_n205_), .B(i_12_), .Y(new_new_n206_));
  NA2        g184(.A(i_0_), .B(i_5_), .Y(new_new_n207_));
  OAI220     g185(.A0(new_new_n76_), .A1(new_new_n178_), .B0(new_new_n170_), .B1(new_new_n125_), .Y(new_new_n208_));
  NAi31      g186(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n36_), .B(i_13_), .Y(new_new_n210_));
  NO2        g188(.A(new_new_n46_), .B(new_new_n58_), .Y(new_new_n211_));
  NA3        g189(.A(new_new_n211_), .B(i_3_), .C(new_new_n210_), .Y(new_new_n212_));
  INV        g190(.A(i_13_), .Y(new_new_n213_));
  NO2        g191(.A(i_12_), .B(new_new_n213_), .Y(new_new_n214_));
  NA3        g192(.A(new_new_n214_), .B(new_new_n187_), .C(new_new_n185_), .Y(new_new_n215_));
  OAI210     g193(.A0(new_new_n212_), .A1(new_new_n209_), .B0(new_new_n215_), .Y(new_new_n216_));
  AOI220     g194(.A0(new_new_n216_), .A1(new_new_n133_), .B0(new_new_n208_), .B1(new_new_n206_), .Y(new_new_n217_));
  NO2        g195(.A(i_12_), .B(new_new_n37_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n172_), .B(i_4_), .Y(new_new_n219_));
  NA2        g197(.A(new_new_n219_), .B(new_new_n218_), .Y(new_new_n220_));
  OR2        g198(.A(i_8_), .B(i_7_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n221_), .B(new_new_n76_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n52_), .B(i_1_), .Y(new_new_n223_));
  INV        g201(.A(i_12_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n44_), .B(new_new_n224_), .Y(new_new_n225_));
  NO3        g203(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n226_));
  NA2        g204(.A(i_2_), .B(i_1_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n52_), .B(new_new_n220_), .Y(new_new_n228_));
  NO3        g206(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n229_));
  NAi21      g207(.An(i_4_), .B(i_3_), .Y(new_new_n230_));
  INV        g208(.A(new_new_n67_), .Y(new_new_n231_));
  NO2        g209(.A(i_0_), .B(i_6_), .Y(new_new_n232_));
  NOi41      g210(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n233_));
  NA2        g211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  NO2        g212(.A(new_new_n227_), .B(new_new_n172_), .Y(new_new_n235_));
  NAi21      g213(.An(new_new_n234_), .B(new_new_n235_), .Y(new_new_n236_));
  INV        g214(.A(new_new_n236_), .Y(new_new_n237_));
  AOI220     g215(.A0(new_new_n237_), .A1(new_new_n40_), .B0(new_new_n228_), .B1(new_new_n196_), .Y(new_new_n238_));
  NO2        g216(.A(i_11_), .B(new_new_n213_), .Y(new_new_n239_));
  NOi21      g217(.An(i_1_), .B(i_6_), .Y(new_new_n240_));
  NAi21      g218(.An(i_3_), .B(i_7_), .Y(new_new_n241_));
  NA2        g219(.A(new_new_n224_), .B(i_9_), .Y(new_new_n242_));
  NO2        g220(.A(i_12_), .B(i_3_), .Y(new_new_n243_));
  NA3        g221(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n244_));
  INV        g222(.A(new_new_n134_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n224_), .B(i_13_), .Y(new_new_n246_));
  NO2        g224(.A(new_new_n246_), .B(new_new_n67_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n247_), .B(new_new_n245_), .Y(new_new_n248_));
  NO2        g226(.A(new_new_n221_), .B(new_new_n37_), .Y(new_new_n249_));
  NA2        g227(.A(i_12_), .B(i_6_), .Y(new_new_n250_));
  OR2        g228(.A(i_13_), .B(i_9_), .Y(new_new_n251_));
  NO3        g229(.A(new_new_n251_), .B(new_new_n250_), .C(new_new_n48_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n230_), .B(i_2_), .Y(new_new_n253_));
  NA3        g231(.A(new_new_n253_), .B(new_new_n252_), .C(new_new_n44_), .Y(new_new_n254_));
  NA2        g232(.A(new_new_n239_), .B(i_9_), .Y(new_new_n255_));
  OAI210     g233(.A0(new_new_n58_), .A1(new_new_n255_), .B0(new_new_n254_), .Y(new_new_n256_));
  NO3        g234(.A(i_11_), .B(new_new_n213_), .C(new_new_n25_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n241_), .B(i_8_), .Y(new_new_n258_));
  NO2        g236(.A(i_6_), .B(new_new_n48_), .Y(new_new_n259_));
  NA3        g237(.A(new_new_n259_), .B(new_new_n258_), .C(new_new_n257_), .Y(new_new_n260_));
  NO3        g238(.A(new_new_n26_), .B(new_new_n76_), .C(i_5_), .Y(new_new_n261_));
  NA3        g239(.A(new_new_n261_), .B(new_new_n249_), .C(new_new_n214_), .Y(new_new_n262_));
  AOI210     g240(.A0(new_new_n262_), .A1(new_new_n260_), .B0(i_1_), .Y(new_new_n263_));
  AOI210     g241(.A0(new_new_n256_), .A1(new_new_n249_), .B0(new_new_n263_), .Y(new_new_n264_));
  NA4        g242(.A(new_new_n264_), .B(new_new_n248_), .C(new_new_n238_), .D(new_new_n217_), .Y(new_new_n265_));
  NO3        g243(.A(i_12_), .B(new_new_n213_), .C(new_new_n37_), .Y(new_new_n266_));
  INV        g244(.A(new_new_n266_), .Y(new_new_n267_));
  NA2        g245(.A(i_8_), .B(new_new_n93_), .Y(new_new_n268_));
  NO3        g246(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n269_));
  AOI220     g247(.A0(new_new_n269_), .A1(new_new_n185_), .B0(new_new_n153_), .B1(new_new_n223_), .Y(new_new_n270_));
  NO2        g248(.A(new_new_n270_), .B(new_new_n268_), .Y(new_new_n271_));
  NO3        g249(.A(i_0_), .B(i_2_), .C(new_new_n58_), .Y(new_new_n272_));
  NO2        g250(.A(new_new_n227_), .B(i_0_), .Y(new_new_n273_));
  AOI220     g251(.A0(new_new_n273_), .A1(new_new_n183_), .B0(new_new_n272_), .B1(new_new_n133_), .Y(new_new_n274_));
  NA2        g252(.A(new_new_n259_), .B(new_new_n26_), .Y(new_new_n275_));
  NO2        g253(.A(new_new_n275_), .B(new_new_n274_), .Y(new_new_n276_));
  NA2        g254(.A(i_0_), .B(i_1_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n277_), .B(i_2_), .Y(new_new_n278_));
  NO2        g256(.A(new_new_n56_), .B(i_6_), .Y(new_new_n279_));
  NA3        g257(.A(new_new_n279_), .B(new_new_n278_), .C(new_new_n153_), .Y(new_new_n280_));
  OAI210     g258(.A0(new_new_n155_), .A1(new_new_n134_), .B0(new_new_n280_), .Y(new_new_n281_));
  NO3        g259(.A(new_new_n281_), .B(new_new_n276_), .C(new_new_n271_), .Y(new_new_n282_));
  NO2        g260(.A(i_3_), .B(i_10_), .Y(new_new_n283_));
  NA3        g261(.A(new_new_n283_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n284_));
  NO2        g262(.A(i_2_), .B(new_new_n93_), .Y(new_new_n285_));
  NA2        g263(.A(i_1_), .B(new_new_n36_), .Y(new_new_n286_));
  NO2        g264(.A(new_new_n286_), .B(i_8_), .Y(new_new_n287_));
  INV        g265(.A(new_new_n287_), .Y(new_new_n288_));
  AN2        g266(.A(i_3_), .B(i_10_), .Y(new_new_n289_));
  NA4        g267(.A(new_new_n289_), .B(new_new_n187_), .C(new_new_n166_), .D(new_new_n164_), .Y(new_new_n290_));
  NO2        g268(.A(i_5_), .B(new_new_n37_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n292_));
  OR2        g270(.A(new_new_n288_), .B(new_new_n284_), .Y(new_new_n293_));
  OAI220     g271(.A0(new_new_n293_), .A1(i_6_), .B0(new_new_n282_), .B1(new_new_n267_), .Y(new_new_n294_));
  NO4        g272(.A(new_new_n294_), .B(new_new_n265_), .C(new_new_n204_), .D(new_new_n158_), .Y(new_new_n295_));
  NO3        g273(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n296_));
  NO3        g274(.A(i_6_), .B(new_new_n182_), .C(i_7_), .Y(new_new_n297_));
  AOI210     g275(.A0(new_new_n967_), .A1(new_new_n227_), .B0(new_new_n159_), .Y(new_new_n298_));
  NO2        g276(.A(i_2_), .B(i_3_), .Y(new_new_n299_));
  OR2        g277(.A(i_0_), .B(i_5_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n207_), .B(new_new_n300_), .Y(new_new_n301_));
  NA4        g279(.A(new_new_n301_), .B(new_new_n222_), .C(new_new_n299_), .D(i_1_), .Y(new_new_n302_));
  NA3        g280(.A(new_new_n273_), .B(new_new_n153_), .C(new_new_n104_), .Y(new_new_n303_));
  NAi21      g281(.An(i_8_), .B(i_7_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n304_), .B(i_6_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n147_), .B(new_new_n46_), .Y(new_new_n306_));
  NA3        g284(.A(new_new_n306_), .B(new_new_n305_), .C(new_new_n153_), .Y(new_new_n307_));
  NA3        g285(.A(new_new_n307_), .B(new_new_n303_), .C(new_new_n302_), .Y(new_new_n308_));
  OAI210     g286(.A0(new_new_n308_), .A1(new_new_n298_), .B0(i_4_), .Y(new_new_n309_));
  NO2        g287(.A(i_12_), .B(i_10_), .Y(new_new_n310_));
  NOi21      g288(.An(i_5_), .B(i_0_), .Y(new_new_n311_));
  NO3        g289(.A(new_new_n286_), .B(new_new_n311_), .C(new_new_n120_), .Y(new_new_n312_));
  NA4        g290(.A(new_new_n74_), .B(new_new_n36_), .C(new_new_n76_), .D(i_8_), .Y(new_new_n313_));
  NA2        g291(.A(new_new_n312_), .B(new_new_n310_), .Y(new_new_n314_));
  NO2        g292(.A(i_6_), .B(i_8_), .Y(new_new_n315_));
  AN2        g293(.A(i_0_), .B(new_new_n315_), .Y(new_new_n316_));
  NO2        g294(.A(i_1_), .B(i_7_), .Y(new_new_n317_));
  AO220      g295(.A0(new_new_n317_), .A1(new_new_n316_), .B0(new_new_n305_), .B1(new_new_n223_), .Y(new_new_n318_));
  NA2        g296(.A(new_new_n318_), .B(i_4_), .Y(new_new_n319_));
  NA3        g297(.A(new_new_n319_), .B(new_new_n314_), .C(new_new_n309_), .Y(new_new_n320_));
  NO3        g298(.A(new_new_n221_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n321_));
  NO3        g299(.A(new_new_n304_), .B(i_2_), .C(i_1_), .Y(new_new_n322_));
  OAI210     g300(.A0(new_new_n322_), .A1(new_new_n321_), .B0(i_6_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n240_), .B(new_new_n285_), .Y(new_new_n324_));
  NA2        g302(.A(new_new_n324_), .B(new_new_n323_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n325_), .B(i_3_), .Y(new_new_n326_));
  INV        g304(.A(new_new_n74_), .Y(new_new_n327_));
  NA2        g305(.A(i_2_), .B(new_new_n124_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n85_), .B(new_new_n182_), .Y(new_new_n329_));
  AOI210     g307(.A0(new_new_n85_), .A1(new_new_n328_), .B0(new_new_n327_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n182_), .B(i_9_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n331_), .B(new_new_n195_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n330_), .B(new_new_n276_), .Y(new_new_n333_));
  AOI210     g311(.A0(new_new_n333_), .A1(new_new_n326_), .B0(new_new_n152_), .Y(new_new_n334_));
  AOI210     g312(.A0(new_new_n320_), .A1(new_new_n296_), .B0(new_new_n334_), .Y(new_new_n335_));
  NOi32      g313(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n336_));
  INV        g314(.A(new_new_n336_), .Y(new_new_n337_));
  NAi21      g315(.An(i_0_), .B(i_6_), .Y(new_new_n338_));
  NAi21      g316(.An(i_1_), .B(i_5_), .Y(new_new_n339_));
  NA2        g317(.A(new_new_n339_), .B(new_new_n338_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n340_), .B(new_new_n25_), .Y(new_new_n341_));
  OAI210     g319(.A0(new_new_n341_), .A1(new_new_n149_), .B0(new_new_n234_), .Y(new_new_n342_));
  NAi41      g320(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n343_));
  OAI220     g321(.A0(new_new_n343_), .A1(new_new_n339_), .B0(new_new_n209_), .B1(new_new_n149_), .Y(new_new_n344_));
  AOI210     g322(.A0(new_new_n343_), .A1(new_new_n149_), .B0(new_new_n147_), .Y(new_new_n345_));
  OR2        g323(.A(new_new_n345_), .B(new_new_n344_), .Y(new_new_n346_));
  NO2        g324(.A(i_1_), .B(new_new_n93_), .Y(new_new_n347_));
  NAi21      g325(.An(i_3_), .B(i_4_), .Y(new_new_n348_));
  NA2        g326(.A(i_2_), .B(i_7_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n348_), .B(i_10_), .Y(new_new_n350_));
  AOI210     g328(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n351_));
  OAI210     g329(.A0(new_new_n351_), .A1(new_new_n177_), .B0(new_new_n350_), .Y(new_new_n352_));
  AOI220     g330(.A0(new_new_n350_), .A1(new_new_n317_), .B0(new_new_n226_), .B1(new_new_n177_), .Y(new_new_n353_));
  AOI210     g331(.A0(new_new_n353_), .A1(new_new_n352_), .B0(i_5_), .Y(new_new_n354_));
  NO3        g332(.A(new_new_n354_), .B(new_new_n346_), .C(new_new_n342_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n355_), .B(new_new_n337_), .Y(new_new_n356_));
  NO2        g334(.A(new_new_n56_), .B(new_new_n25_), .Y(new_new_n357_));
  AN2        g335(.A(i_12_), .B(i_5_), .Y(new_new_n358_));
  NO2        g336(.A(i_4_), .B(new_new_n26_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n359_), .B(new_new_n358_), .Y(new_new_n360_));
  NO2        g338(.A(i_11_), .B(i_6_), .Y(new_new_n361_));
  NA3        g339(.A(new_new_n361_), .B(new_new_n306_), .C(new_new_n213_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n362_), .B(new_new_n360_), .Y(new_new_n363_));
  NO2        g341(.A(new_new_n230_), .B(i_5_), .Y(new_new_n364_));
  NO2        g342(.A(i_5_), .B(i_10_), .Y(new_new_n365_));
  AOI220     g343(.A0(new_new_n365_), .A1(new_new_n253_), .B0(new_new_n364_), .B1(new_new_n187_), .Y(new_new_n366_));
  NA2        g344(.A(new_new_n135_), .B(new_new_n45_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n367_), .B(new_new_n366_), .Y(new_new_n368_));
  OAI210     g346(.A0(new_new_n368_), .A1(new_new_n363_), .B0(new_new_n357_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n370_));
  NO2        g348(.A(new_new_n141_), .B(new_new_n76_), .Y(new_new_n371_));
  OAI210     g349(.A0(new_new_n371_), .A1(new_new_n363_), .B0(new_new_n370_), .Y(new_new_n372_));
  NO3        g350(.A(new_new_n76_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n373_));
  NA3        g351(.A(new_new_n283_), .B(new_new_n83_), .C(new_new_n53_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n374_), .B(i_12_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n365_), .B(new_new_n224_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n36_), .B(new_new_n209_), .Y(new_new_n377_));
  NAi21      g355(.An(i_13_), .B(i_0_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n378_), .B(new_new_n227_), .Y(new_new_n379_));
  OAI210     g357(.A0(new_new_n377_), .A1(new_new_n375_), .B0(new_new_n379_), .Y(new_new_n380_));
  NA3        g358(.A(new_new_n380_), .B(new_new_n372_), .C(new_new_n369_), .Y(new_new_n381_));
  NA2        g359(.A(new_new_n44_), .B(new_new_n213_), .Y(new_new_n382_));
  NO2        g360(.A(i_0_), .B(i_11_), .Y(new_new_n383_));
  INV        g361(.A(i_5_), .Y(new_new_n384_));
  AN2        g362(.A(i_1_), .B(i_6_), .Y(new_new_n385_));
  NOi21      g363(.An(i_2_), .B(i_12_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n386_), .B(new_new_n385_), .Y(new_new_n387_));
  NO2        g365(.A(new_new_n387_), .B(new_new_n384_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n133_), .B(i_9_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n389_), .B(i_4_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n388_), .B(new_new_n390_), .Y(new_new_n391_));
  NAi21      g369(.An(i_9_), .B(i_4_), .Y(new_new_n392_));
  OR2        g370(.A(i_13_), .B(i_10_), .Y(new_new_n393_));
  NO3        g371(.A(new_new_n393_), .B(new_new_n109_), .C(new_new_n392_), .Y(new_new_n394_));
  BUFFER     g372(.A(new_new_n205_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n93_), .B(new_new_n25_), .Y(new_new_n396_));
  NA2        g374(.A(new_new_n259_), .B(new_new_n200_), .Y(new_new_n397_));
  NO2        g375(.A(new_new_n397_), .B(new_new_n395_), .Y(new_new_n398_));
  INV        g376(.A(new_new_n398_), .Y(new_new_n399_));
  AOI210     g377(.A0(new_new_n399_), .A1(new_new_n391_), .B0(new_new_n26_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n303_), .B(new_new_n302_), .Y(new_new_n401_));
  AOI220     g379(.A0(new_new_n279_), .A1(new_new_n269_), .B0(new_new_n273_), .B1(i_6_), .Y(new_new_n402_));
  NO2        g380(.A(new_new_n402_), .B(new_new_n159_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n172_), .B(new_new_n76_), .Y(new_new_n404_));
  AOI220     g382(.A0(new_new_n404_), .A1(new_new_n278_), .B0(new_new_n261_), .B1(new_new_n200_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n405_), .B(new_new_n268_), .Y(new_new_n406_));
  NO3        g384(.A(new_new_n406_), .B(new_new_n403_), .C(new_new_n401_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n185_), .B(new_new_n88_), .Y(new_new_n408_));
  NA3        g386(.A(new_new_n306_), .B(new_new_n153_), .C(new_new_n76_), .Y(new_new_n409_));
  AOI210     g387(.A0(new_new_n409_), .A1(new_new_n408_), .B0(new_new_n304_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n279_), .B(new_new_n223_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n411_), .B(new_new_n172_), .Y(new_new_n412_));
  NA3        g390(.A(new_new_n317_), .B(new_new_n316_), .C(i_5_), .Y(new_new_n413_));
  INV        g391(.A(new_new_n297_), .Y(new_new_n414_));
  OAI210     g392(.A0(new_new_n414_), .A1(new_new_n178_), .B0(new_new_n413_), .Y(new_new_n415_));
  NO3        g393(.A(new_new_n415_), .B(new_new_n412_), .C(new_new_n410_), .Y(new_new_n416_));
  AOI210     g394(.A0(new_new_n416_), .A1(new_new_n407_), .B0(new_new_n255_), .Y(new_new_n417_));
  NO4        g395(.A(new_new_n417_), .B(new_new_n400_), .C(new_new_n381_), .D(new_new_n356_), .Y(new_new_n418_));
  NO2        g396(.A(i_10_), .B(i_9_), .Y(new_new_n419_));
  NAi21      g397(.An(i_12_), .B(i_8_), .Y(new_new_n420_));
  NO2        g398(.A(new_new_n420_), .B(i_3_), .Y(new_new_n421_));
  NA2        g399(.A(i_2_), .B(new_new_n96_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n422_), .B(new_new_n194_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n292_), .B(i_0_), .Y(new_new_n424_));
  NO3        g402(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n425_));
  NA2        g403(.A(new_new_n250_), .B(new_new_n89_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n426_), .B(new_new_n425_), .Y(new_new_n427_));
  NA2        g405(.A(i_8_), .B(i_9_), .Y(new_new_n428_));
  NO2        g406(.A(i_7_), .B(i_2_), .Y(new_new_n429_));
  OR2        g407(.A(new_new_n429_), .B(new_new_n428_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n266_), .B(new_new_n195_), .Y(new_new_n431_));
  NO2        g409(.A(new_new_n431_), .B(new_new_n430_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n239_), .B(new_new_n291_), .Y(new_new_n433_));
  NO3        g411(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n434_));
  INV        g412(.A(new_new_n434_), .Y(new_new_n435_));
  NA3        g413(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n436_));
  NA4        g414(.A(new_new_n136_), .B(new_new_n107_), .C(new_new_n72_), .D(new_new_n23_), .Y(new_new_n437_));
  OAI220     g415(.A0(new_new_n437_), .A1(new_new_n436_), .B0(new_new_n435_), .B1(new_new_n433_), .Y(new_new_n438_));
  NO3        g416(.A(new_new_n438_), .B(new_new_n432_), .C(new_new_n423_), .Y(new_new_n439_));
  OR2        g417(.A(new_new_n277_), .B(new_new_n197_), .Y(new_new_n440_));
  OA210      g418(.A0(new_new_n332_), .A1(new_new_n93_), .B0(new_new_n280_), .Y(new_new_n441_));
  OA220      g419(.A0(new_new_n441_), .A1(new_new_n152_), .B0(new_new_n440_), .B1(new_new_n220_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n88_), .B(i_13_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n404_), .B(new_new_n357_), .Y(new_new_n444_));
  NO2        g422(.A(i_2_), .B(i_13_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n444_), .B(new_new_n443_), .Y(new_new_n446_));
  NO3        g424(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n447_));
  NO2        g425(.A(i_6_), .B(i_7_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n448_), .B(new_new_n447_), .Y(new_new_n449_));
  NO2        g427(.A(i_11_), .B(i_1_), .Y(new_new_n450_));
  NOi21      g428(.An(i_2_), .B(i_7_), .Y(new_new_n451_));
  NO2        g429(.A(i_3_), .B(new_new_n182_), .Y(new_new_n452_));
  NO2        g430(.A(i_6_), .B(i_10_), .Y(new_new_n453_));
  NA3        g431(.A(new_new_n453_), .B(new_new_n296_), .C(new_new_n452_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n454_), .B(new_new_n145_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n456_));
  NO2        g434(.A(new_new_n147_), .B(i_3_), .Y(new_new_n457_));
  NAi31      g435(.An(new_new_n456_), .B(new_new_n457_), .C(new_new_n214_), .Y(new_new_n458_));
  NA3        g436(.A(new_new_n370_), .B(new_new_n169_), .C(new_new_n140_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n459_), .B(new_new_n458_), .Y(new_new_n460_));
  NO3        g438(.A(new_new_n460_), .B(new_new_n455_), .C(new_new_n446_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n425_), .B(new_new_n358_), .Y(new_new_n462_));
  NA2        g440(.A(new_new_n434_), .B(new_new_n365_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n463_), .B(new_new_n212_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n26_), .B(i_5_), .Y(new_new_n465_));
  NA3        g443(.A(new_new_n966_), .B(new_new_n465_), .C(new_new_n133_), .Y(new_new_n466_));
  OR3        g444(.A(new_new_n286_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n467_), .B(new_new_n466_), .Y(new_new_n468_));
  NA2        g446(.A(new_new_n27_), .B(i_10_), .Y(new_new_n469_));
  NO2        g447(.A(new_new_n469_), .B(new_new_n443_), .Y(new_new_n470_));
  NA3        g448(.A(new_new_n289_), .B(new_new_n211_), .C(new_new_n65_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n471_), .B(new_new_n449_), .Y(new_new_n472_));
  NO4        g450(.A(new_new_n472_), .B(new_new_n470_), .C(new_new_n468_), .D(new_new_n464_), .Y(new_new_n473_));
  NA4        g451(.A(new_new_n473_), .B(new_new_n461_), .C(new_new_n442_), .D(new_new_n439_), .Y(new_new_n474_));
  AN2        g452(.A(new_new_n269_), .B(new_new_n222_), .Y(new_new_n475_));
  NA2        g453(.A(new_new_n475_), .B(new_new_n166_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n114_), .B(new_new_n103_), .Y(new_new_n477_));
  AN2        g455(.A(new_new_n477_), .B(new_new_n425_), .Y(new_new_n478_));
  NA2        g456(.A(new_new_n296_), .B(new_new_n154_), .Y(new_new_n479_));
  OAI210     g457(.A0(new_new_n479_), .A1(new_new_n220_), .B0(new_new_n290_), .Y(new_new_n480_));
  AOI220     g458(.A0(new_new_n480_), .A1(new_new_n305_), .B0(new_new_n478_), .B1(new_new_n292_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n336_), .B(new_new_n65_), .Y(new_new_n482_));
  NO2        g460(.A(new_new_n36_), .B(i_8_), .Y(new_new_n483_));
  AOI210     g461(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n394_), .Y(new_new_n484_));
  NO2        g462(.A(i_7_), .B(new_new_n188_), .Y(new_new_n485_));
  OR2        g463(.A(new_new_n172_), .B(i_4_), .Y(new_new_n486_));
  INV        g464(.A(new_new_n486_), .Y(new_new_n487_));
  NA2        g465(.A(new_new_n487_), .B(new_new_n485_), .Y(new_new_n488_));
  NA4        g466(.A(new_new_n488_), .B(new_new_n484_), .C(new_new_n481_), .D(new_new_n476_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n364_), .B(new_new_n278_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n360_), .B(new_new_n490_), .Y(new_new_n491_));
  NO2        g469(.A(i_12_), .B(new_new_n182_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n453_), .B(new_new_n27_), .Y(new_new_n493_));
  NO2        g471(.A(new_new_n493_), .B(i_12_), .Y(new_new_n494_));
  NOi31      g472(.An(new_new_n297_), .B(new_new_n393_), .C(new_new_n38_), .Y(new_new_n495_));
  OAI210     g473(.A0(new_new_n495_), .A1(new_new_n494_), .B0(new_new_n491_), .Y(new_new_n496_));
  NO2        g474(.A(i_8_), .B(i_7_), .Y(new_new_n497_));
  OAI210     g475(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n498_));
  NA2        g476(.A(new_new_n498_), .B(new_new_n211_), .Y(new_new_n499_));
  OAI220     g477(.A0(new_new_n46_), .A1(new_new_n486_), .B0(new_new_n499_), .B1(new_new_n230_), .Y(new_new_n500_));
  NA2        g478(.A(new_new_n44_), .B(i_10_), .Y(new_new_n501_));
  NO2        g479(.A(new_new_n501_), .B(i_6_), .Y(new_new_n502_));
  NA3        g480(.A(new_new_n502_), .B(new_new_n500_), .C(new_new_n497_), .Y(new_new_n503_));
  AOI220     g481(.A0(new_new_n404_), .A1(new_new_n306_), .B0(new_new_n235_), .B1(new_new_n232_), .Y(new_new_n504_));
  OAI220     g482(.A0(new_new_n504_), .A1(new_new_n246_), .B0(new_new_n443_), .B1(new_new_n125_), .Y(new_new_n505_));
  NA2        g483(.A(new_new_n505_), .B(new_new_n249_), .Y(new_new_n506_));
  NA3        g484(.A(new_new_n289_), .B(new_new_n164_), .C(new_new_n88_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n210_), .B(new_new_n44_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n147_), .B(i_5_), .Y(new_new_n509_));
  NA3        g487(.A(new_new_n509_), .B(new_new_n382_), .C(new_new_n299_), .Y(new_new_n510_));
  OAI210     g488(.A0(new_new_n510_), .A1(new_new_n508_), .B0(new_new_n507_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n511_), .B(new_new_n434_), .Y(new_new_n512_));
  NA4        g490(.A(new_new_n512_), .B(new_new_n506_), .C(new_new_n503_), .D(new_new_n496_), .Y(new_new_n513_));
  NA3        g491(.A(new_new_n207_), .B(new_new_n63_), .C(new_new_n44_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n266_), .B(new_new_n74_), .Y(new_new_n515_));
  AOI210     g493(.A0(new_new_n514_), .A1(new_new_n328_), .B0(new_new_n515_), .Y(new_new_n516_));
  NO2        g494(.A(new_new_n46_), .B(new_new_n163_), .Y(new_new_n517_));
  AOI210     g495(.A0(i_6_), .A1(new_new_n46_), .B0(new_new_n347_), .Y(new_new_n518_));
  NA2        g496(.A(i_0_), .B(new_new_n48_), .Y(new_new_n519_));
  NA3        g497(.A(new_new_n492_), .B(new_new_n257_), .C(new_new_n519_), .Y(new_new_n520_));
  NO2        g498(.A(new_new_n518_), .B(new_new_n520_), .Y(new_new_n521_));
  NO3        g499(.A(new_new_n521_), .B(new_new_n517_), .C(new_new_n516_), .Y(new_new_n522_));
  NO4        g500(.A(new_new_n240_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n523_));
  NO3        g501(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n524_));
  NO2        g502(.A(new_new_n221_), .B(new_new_n36_), .Y(new_new_n525_));
  AN2        g503(.A(new_new_n525_), .B(new_new_n524_), .Y(new_new_n526_));
  OA210      g504(.A0(new_new_n526_), .A1(new_new_n523_), .B0(new_new_n336_), .Y(new_new_n527_));
  NO2        g505(.A(new_new_n393_), .B(i_1_), .Y(new_new_n528_));
  NOi31      g506(.An(new_new_n528_), .B(new_new_n426_), .C(new_new_n65_), .Y(new_new_n529_));
  AN4        g507(.A(new_new_n529_), .B(new_new_n390_), .C(new_new_n465_), .D(i_2_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n402_), .B(new_new_n167_), .Y(new_new_n531_));
  NO3        g509(.A(new_new_n531_), .B(new_new_n530_), .C(new_new_n527_), .Y(new_new_n532_));
  NOi21      g510(.An(i_10_), .B(i_6_), .Y(new_new_n533_));
  NO2        g511(.A(new_new_n76_), .B(new_new_n25_), .Y(new_new_n534_));
  AOI220     g512(.A0(new_new_n266_), .A1(new_new_n534_), .B0(new_new_n257_), .B1(new_new_n533_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n535_), .B(new_new_n424_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n106_), .B(new_new_n23_), .Y(new_new_n537_));
  NA2        g515(.A(new_new_n297_), .B(new_new_n154_), .Y(new_new_n538_));
  AOI220     g516(.A0(new_new_n538_), .A1(new_new_n411_), .B0(new_new_n162_), .B1(new_new_n171_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n187_), .B(new_new_n37_), .Y(new_new_n540_));
  NOi31      g518(.An(new_new_n137_), .B(new_new_n540_), .C(new_new_n313_), .Y(new_new_n541_));
  NO3        g519(.A(new_new_n541_), .B(new_new_n539_), .C(new_new_n536_), .Y(new_new_n542_));
  NO2        g520(.A(new_new_n482_), .B(new_new_n353_), .Y(new_new_n543_));
  NO2        g521(.A(i_12_), .B(new_new_n76_), .Y(new_new_n544_));
  NO3        g522(.A(i_4_), .B(new_new_n323_), .C(new_new_n284_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n545_), .B(new_new_n543_), .Y(new_new_n546_));
  NA4        g524(.A(new_new_n546_), .B(new_new_n542_), .C(new_new_n532_), .D(new_new_n522_), .Y(new_new_n547_));
  NO4        g525(.A(new_new_n547_), .B(new_new_n513_), .C(new_new_n489_), .D(new_new_n474_), .Y(new_new_n548_));
  NA4        g526(.A(new_new_n548_), .B(new_new_n418_), .C(new_new_n335_), .D(new_new_n295_), .Y(mai7));
  NO2        g527(.A(new_new_n100_), .B(new_new_n82_), .Y(new_new_n550_));
  NA2        g528(.A(new_new_n453_), .B(new_new_n74_), .Y(new_new_n551_));
  NA2        g529(.A(i_11_), .B(new_new_n182_), .Y(new_new_n552_));
  NA3        g530(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n224_), .B(i_4_), .Y(new_new_n554_));
  NA2        g532(.A(new_new_n554_), .B(i_8_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n97_), .B(new_new_n553_), .Y(new_new_n556_));
  NA2        g534(.A(i_2_), .B(new_new_n76_), .Y(new_new_n557_));
  OAI210     g535(.A0(new_new_n79_), .A1(new_new_n192_), .B0(new_new_n193_), .Y(new_new_n558_));
  NO2        g536(.A(i_7_), .B(new_new_n37_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n558_), .B(i_13_), .Y(new_new_n560_));
  NO3        g538(.A(new_new_n560_), .B(new_new_n556_), .C(new_new_n550_), .Y(new_new_n561_));
  AOI210     g539(.A0(new_new_n120_), .A1(new_new_n57_), .B0(i_10_), .Y(new_new_n562_));
  AOI210     g540(.A0(new_new_n562_), .A1(new_new_n224_), .B0(new_new_n151_), .Y(new_new_n563_));
  OR2        g541(.A(i_6_), .B(i_10_), .Y(new_new_n564_));
  NO2        g542(.A(new_new_n564_), .B(new_new_n23_), .Y(new_new_n565_));
  OR3        g543(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n566_));
  NO3        g544(.A(new_new_n566_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n567_));
  INV        g545(.A(new_new_n189_), .Y(new_new_n568_));
  NO2        g546(.A(new_new_n567_), .B(new_new_n565_), .Y(new_new_n569_));
  OA220      g547(.A0(new_new_n569_), .A1(i_2_), .B0(new_new_n563_), .B1(new_new_n251_), .Y(new_new_n570_));
  AOI210     g548(.A0(new_new_n570_), .A1(new_new_n561_), .B0(new_new_n58_), .Y(new_new_n571_));
  NOi21      g549(.An(i_11_), .B(i_7_), .Y(new_new_n572_));
  AO210      g550(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n573_));
  NO2        g551(.A(new_new_n573_), .B(new_new_n572_), .Y(new_new_n574_));
  NA2        g552(.A(new_new_n574_), .B(new_new_n196_), .Y(new_new_n575_));
  NA3        g553(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n576_));
  NAi31      g554(.An(new_new_n576_), .B(i_12_), .C(i_11_), .Y(new_new_n577_));
  AOI210     g555(.A0(new_new_n577_), .A1(new_new_n575_), .B0(new_new_n58_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n78_), .B(new_new_n58_), .Y(new_new_n579_));
  AO210      g557(.A0(new_new_n579_), .A1(new_new_n353_), .B0(new_new_n41_), .Y(new_new_n580_));
  NA2        g558(.A(new_new_n214_), .B(new_new_n58_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n58_), .B(i_9_), .Y(new_new_n582_));
  NO2        g560(.A(i_1_), .B(i_12_), .Y(new_new_n583_));
  NA2        g561(.A(new_new_n581_), .B(new_new_n580_), .Y(new_new_n584_));
  OAI210     g562(.A0(new_new_n584_), .A1(new_new_n578_), .B0(i_6_), .Y(new_new_n585_));
  NO2        g563(.A(new_new_n576_), .B(new_new_n100_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n586_), .B(new_new_n544_), .Y(new_new_n587_));
  NO2        g565(.A(new_new_n224_), .B(new_new_n76_), .Y(new_new_n588_));
  NO2        g566(.A(new_new_n588_), .B(i_11_), .Y(new_new_n589_));
  NA2        g567(.A(new_new_n587_), .B(new_new_n427_), .Y(new_new_n590_));
  NO4        g568(.A(i_12_), .B(new_new_n120_), .C(i_13_), .D(new_new_n76_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n591_), .B(new_new_n582_), .Y(new_new_n592_));
  NA2        g570(.A(new_new_n224_), .B(i_6_), .Y(new_new_n593_));
  INV        g571(.A(new_new_n592_), .Y(new_new_n594_));
  NA3        g572(.A(new_new_n497_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n129_), .B(i_9_), .Y(new_new_n596_));
  NA2        g574(.A(i_3_), .B(i_9_), .Y(new_new_n597_));
  NO2        g575(.A(new_new_n46_), .B(i_1_), .Y(new_new_n598_));
  NO2        g576(.A(new_new_n596_), .B(new_new_n964_), .Y(new_new_n599_));
  NA3        g577(.A(new_new_n582_), .B(new_new_n299_), .C(i_6_), .Y(new_new_n600_));
  NO2        g578(.A(new_new_n600_), .B(new_new_n23_), .Y(new_new_n601_));
  AOI210     g579(.A0(new_new_n450_), .A1(new_new_n396_), .B0(new_new_n229_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n602_), .B(new_new_n557_), .Y(new_new_n603_));
  NA2        g581(.A(new_new_n598_), .B(new_new_n250_), .Y(new_new_n604_));
  NO2        g582(.A(i_11_), .B(new_new_n37_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n605_), .B(new_new_n24_), .Y(new_new_n606_));
  NO2        g584(.A(new_new_n606_), .B(new_new_n604_), .Y(new_new_n607_));
  OR4        g585(.A(new_new_n607_), .B(new_new_n603_), .C(new_new_n601_), .D(new_new_n599_), .Y(new_new_n608_));
  NO3        g586(.A(new_new_n608_), .B(new_new_n594_), .C(new_new_n590_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n224_), .B(new_new_n93_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n610_), .B(new_new_n572_), .Y(new_new_n611_));
  NO2        g589(.A(new_new_n392_), .B(new_new_n76_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n221_), .B(new_new_n44_), .Y(new_new_n613_));
  NO3        g591(.A(new_new_n613_), .B(new_new_n292_), .C(new_new_n225_), .Y(new_new_n614_));
  NO2        g592(.A(new_new_n109_), .B(new_new_n37_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n615_), .B(i_6_), .Y(new_new_n616_));
  NO2        g594(.A(new_new_n76_), .B(i_9_), .Y(new_new_n617_));
  NO2        g595(.A(new_new_n617_), .B(new_new_n58_), .Y(new_new_n618_));
  NO2        g596(.A(new_new_n618_), .B(new_new_n583_), .Y(new_new_n619_));
  NO4        g597(.A(new_new_n619_), .B(new_new_n616_), .C(new_new_n614_), .D(i_4_), .Y(new_new_n620_));
  NA2        g598(.A(i_1_), .B(i_3_), .Y(new_new_n621_));
  INV        g599(.A(new_new_n620_), .Y(new_new_n622_));
  NA3        g600(.A(new_new_n622_), .B(new_new_n609_), .C(new_new_n585_), .Y(new_new_n623_));
  NO3        g601(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n624_));
  NOi21      g602(.An(new_new_n624_), .B(i_10_), .Y(new_new_n625_));
  OA210      g603(.A0(new_new_n625_), .A1(new_new_n233_), .B0(new_new_n76_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n626_), .B(i_1_), .Y(new_new_n627_));
  AOI210     g605(.A0(new_new_n250_), .A1(new_new_n89_), .B0(i_1_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n348_), .B(i_2_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n629_), .B(new_new_n628_), .Y(new_new_n630_));
  AOI210     g608(.A0(new_new_n630_), .A1(new_new_n627_), .B0(i_13_), .Y(new_new_n631_));
  OR2        g609(.A(i_11_), .B(i_7_), .Y(new_new_n632_));
  NA3        g610(.A(new_new_n632_), .B(new_new_n98_), .C(new_new_n129_), .Y(new_new_n633_));
  AOI220     g611(.A0(new_new_n445_), .A1(new_new_n151_), .B0(i_2_), .B1(new_new_n129_), .Y(new_new_n634_));
  OAI210     g612(.A0(new_new_n634_), .A1(new_new_n44_), .B0(new_new_n633_), .Y(new_new_n635_));
  NO2        g613(.A(new_new_n53_), .B(i_12_), .Y(new_new_n636_));
  INV        g614(.A(new_new_n636_), .Y(new_new_n637_));
  NO2        g615(.A(new_new_n451_), .B(new_new_n24_), .Y(new_new_n638_));
  NA2        g616(.A(new_new_n638_), .B(new_new_n612_), .Y(new_new_n639_));
  OAI220     g617(.A0(new_new_n639_), .A1(new_new_n41_), .B0(new_new_n637_), .B1(new_new_n85_), .Y(new_new_n640_));
  AOI210     g618(.A0(new_new_n635_), .A1(new_new_n315_), .B0(new_new_n640_), .Y(new_new_n641_));
  INV        g619(.A(new_new_n106_), .Y(new_new_n642_));
  AOI220     g620(.A0(new_new_n642_), .A1(new_new_n64_), .B0(new_new_n361_), .B1(new_new_n598_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n643_), .B(new_new_n230_), .Y(new_new_n644_));
  AOI210     g622(.A0(new_new_n420_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n645_));
  NOi31      g623(.An(new_new_n645_), .B(new_new_n551_), .C(new_new_n44_), .Y(new_new_n646_));
  NA2        g624(.A(new_new_n119_), .B(i_13_), .Y(new_new_n647_));
  NO2        g625(.A(new_new_n597_), .B(new_new_n106_), .Y(new_new_n648_));
  INV        g626(.A(new_new_n648_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n647_), .B(new_new_n628_), .Y(new_new_n650_));
  AOI220     g628(.A0(new_new_n361_), .A1(new_new_n598_), .B0(new_new_n84_), .B1(new_new_n94_), .Y(new_new_n651_));
  NO2        g629(.A(new_new_n651_), .B(new_new_n555_), .Y(new_new_n652_));
  NO4        g630(.A(new_new_n652_), .B(new_new_n650_), .C(new_new_n646_), .D(new_new_n644_), .Y(new_new_n653_));
  OR2        g631(.A(i_11_), .B(i_6_), .Y(new_new_n654_));
  NA2        g632(.A(new_new_n554_), .B(i_7_), .Y(new_new_n655_));
  AOI210     g633(.A0(new_new_n655_), .A1(new_new_n649_), .B0(new_new_n654_), .Y(new_new_n656_));
  NA3        g634(.A(new_new_n386_), .B(new_new_n559_), .C(new_new_n89_), .Y(new_new_n657_));
  NA2        g635(.A(new_new_n589_), .B(i_13_), .Y(new_new_n658_));
  NAi21      g636(.An(i_11_), .B(i_12_), .Y(new_new_n659_));
  NOi41      g637(.An(new_new_n102_), .B(new_new_n659_), .C(i_13_), .D(new_new_n76_), .Y(new_new_n660_));
  NA2        g638(.A(new_new_n660_), .B(new_new_n46_), .Y(new_new_n661_));
  NA3        g639(.A(new_new_n661_), .B(new_new_n658_), .C(new_new_n657_), .Y(new_new_n662_));
  OAI210     g640(.A0(new_new_n662_), .A1(new_new_n656_), .B0(new_new_n58_), .Y(new_new_n663_));
  NO2        g641(.A(i_2_), .B(i_12_), .Y(new_new_n664_));
  NA2        g642(.A(new_new_n347_), .B(new_new_n664_), .Y(new_new_n665_));
  NO3        g643(.A(i_9_), .B(new_new_n359_), .C(new_new_n554_), .Y(new_new_n666_));
  NA2        g644(.A(new_new_n666_), .B(new_new_n347_), .Y(new_new_n667_));
  NO2        g645(.A(new_new_n120_), .B(i_2_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n668_), .B(new_new_n583_), .Y(new_new_n669_));
  NA3        g647(.A(new_new_n669_), .B(new_new_n667_), .C(new_new_n665_), .Y(new_new_n670_));
  NA3        g648(.A(new_new_n670_), .B(new_new_n45_), .C(new_new_n213_), .Y(new_new_n671_));
  NA4        g649(.A(new_new_n671_), .B(new_new_n663_), .C(new_new_n653_), .D(new_new_n641_), .Y(new_new_n672_));
  OR4        g650(.A(new_new_n672_), .B(new_new_n631_), .C(new_new_n623_), .D(new_new_n571_), .Y(mai5));
  NA2        g651(.A(new_new_n611_), .B(new_new_n253_), .Y(new_new_n674_));
  AN2        g652(.A(new_new_n24_), .B(i_10_), .Y(new_new_n675_));
  NA3        g653(.A(new_new_n675_), .B(new_new_n664_), .C(new_new_n100_), .Y(new_new_n676_));
  NO2        g654(.A(new_new_n555_), .B(i_11_), .Y(new_new_n677_));
  NA2        g655(.A(new_new_n79_), .B(new_new_n677_), .Y(new_new_n678_));
  NA3        g656(.A(new_new_n678_), .B(new_new_n676_), .C(new_new_n674_), .Y(new_new_n679_));
  NO3        g657(.A(i_11_), .B(new_new_n224_), .C(i_13_), .Y(new_new_n680_));
  NO2        g658(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n681_));
  NA2        g659(.A(i_12_), .B(i_8_), .Y(new_new_n682_));
  OAI210     g660(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n682_), .Y(new_new_n683_));
  INV        g661(.A(new_new_n419_), .Y(new_new_n684_));
  AOI220     g662(.A0(new_new_n299_), .A1(new_new_n537_), .B0(new_new_n683_), .B1(new_new_n681_), .Y(new_new_n685_));
  INV        g663(.A(new_new_n685_), .Y(new_new_n686_));
  NO2        g664(.A(new_new_n686_), .B(new_new_n679_), .Y(new_new_n687_));
  INV        g665(.A(new_new_n161_), .Y(new_new_n688_));
  INV        g666(.A(new_new_n233_), .Y(new_new_n689_));
  OAI210     g667(.A0(new_new_n629_), .A1(new_new_n421_), .B0(new_new_n102_), .Y(new_new_n690_));
  AOI210     g668(.A0(new_new_n690_), .A1(new_new_n689_), .B0(new_new_n688_), .Y(new_new_n691_));
  NO2        g669(.A(new_new_n428_), .B(new_new_n26_), .Y(new_new_n692_));
  NO2        g670(.A(new_new_n692_), .B(new_new_n396_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n693_), .B(i_2_), .Y(new_new_n694_));
  INV        g672(.A(new_new_n694_), .Y(new_new_n695_));
  AOI210     g673(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n393_), .Y(new_new_n696_));
  AOI210     g674(.A0(new_new_n696_), .A1(new_new_n695_), .B0(new_new_n691_), .Y(new_new_n697_));
  NO2        g675(.A(new_new_n179_), .B(new_new_n117_), .Y(new_new_n698_));
  OAI210     g676(.A0(new_new_n698_), .A1(new_new_n681_), .B0(i_2_), .Y(new_new_n699_));
  INV        g677(.A(new_new_n162_), .Y(new_new_n700_));
  NO3        g678(.A(new_new_n573_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n701_));
  AOI210     g679(.A0(new_new_n700_), .A1(new_new_n79_), .B0(new_new_n701_), .Y(new_new_n702_));
  AOI210     g680(.A0(new_new_n702_), .A1(new_new_n699_), .B0(new_new_n182_), .Y(new_new_n703_));
  OA210      g681(.A0(new_new_n574_), .A1(new_new_n118_), .B0(i_13_), .Y(new_new_n704_));
  INV        g682(.A(new_new_n142_), .Y(new_new_n705_));
  NO2        g683(.A(new_new_n705_), .B(new_new_n349_), .Y(new_new_n706_));
  NO2        g684(.A(new_new_n139_), .B(new_new_n483_), .Y(new_new_n707_));
  NA2        g685(.A(new_new_n707_), .B(new_new_n396_), .Y(new_new_n708_));
  NO2        g686(.A(new_new_n94_), .B(new_new_n44_), .Y(new_new_n709_));
  INV        g687(.A(new_new_n285_), .Y(new_new_n710_));
  NA4        g688(.A(new_new_n710_), .B(new_new_n289_), .C(new_new_n116_), .D(new_new_n42_), .Y(new_new_n711_));
  OAI210     g689(.A0(new_new_n711_), .A1(new_new_n709_), .B0(new_new_n708_), .Y(new_new_n712_));
  NO4        g690(.A(new_new_n712_), .B(new_new_n706_), .C(new_new_n704_), .D(new_new_n703_), .Y(new_new_n713_));
  NA2        g691(.A(new_new_n537_), .B(new_new_n28_), .Y(new_new_n714_));
  NA2        g692(.A(new_new_n680_), .B(new_new_n258_), .Y(new_new_n715_));
  NA2        g693(.A(new_new_n715_), .B(new_new_n714_), .Y(new_new_n716_));
  NO2        g694(.A(new_new_n57_), .B(i_12_), .Y(new_new_n717_));
  NO2        g695(.A(new_new_n717_), .B(new_new_n118_), .Y(new_new_n718_));
  NO2        g696(.A(new_new_n718_), .B(new_new_n552_), .Y(new_new_n719_));
  AOI220     g697(.A0(new_new_n719_), .A1(new_new_n36_), .B0(new_new_n716_), .B1(new_new_n46_), .Y(new_new_n720_));
  NA4        g698(.A(new_new_n720_), .B(new_new_n713_), .C(new_new_n697_), .D(new_new_n687_), .Y(mai6));
  NO3        g699(.A(i_9_), .B(new_new_n291_), .C(i_1_), .Y(new_new_n722_));
  NO2        g700(.A(new_new_n174_), .B(new_new_n130_), .Y(new_new_n723_));
  OAI210     g701(.A0(new_new_n723_), .A1(new_new_n722_), .B0(new_new_n668_), .Y(new_new_n724_));
  NA4        g702(.A(new_new_n365_), .B(new_new_n452_), .C(new_new_n63_), .D(new_new_n93_), .Y(new_new_n725_));
  INV        g703(.A(new_new_n725_), .Y(new_new_n726_));
  NO2        g704(.A(i_11_), .B(i_9_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n726_), .B(new_new_n311_), .Y(new_new_n728_));
  AO210      g706(.A0(new_new_n728_), .A1(new_new_n724_), .B0(i_12_), .Y(new_new_n729_));
  NA2        g707(.A(new_new_n350_), .B(new_new_n317_), .Y(new_new_n730_));
  NA2        g708(.A(new_new_n544_), .B(new_new_n58_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n625_), .B(new_new_n63_), .Y(new_new_n732_));
  BUFFER     g710(.A(new_new_n579_), .Y(new_new_n733_));
  NA4        g711(.A(new_new_n733_), .B(new_new_n732_), .C(new_new_n731_), .D(new_new_n730_), .Y(new_new_n734_));
  INV        g712(.A(new_new_n186_), .Y(new_new_n735_));
  AOI220     g713(.A0(new_new_n735_), .A1(new_new_n727_), .B0(new_new_n734_), .B1(new_new_n65_), .Y(new_new_n736_));
  INV        g714(.A(new_new_n310_), .Y(new_new_n737_));
  NA2        g715(.A(new_new_n67_), .B(new_new_n123_), .Y(new_new_n738_));
  INV        g716(.A(new_new_n116_), .Y(new_new_n739_));
  NA2        g717(.A(new_new_n739_), .B(new_new_n46_), .Y(new_new_n740_));
  AOI210     g718(.A0(new_new_n740_), .A1(new_new_n738_), .B0(new_new_n737_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n240_), .B(i_9_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n742_), .B(new_new_n717_), .Y(new_new_n743_));
  NO2        g721(.A(new_new_n743_), .B(new_new_n174_), .Y(new_new_n744_));
  NO2        g722(.A(new_new_n32_), .B(i_11_), .Y(new_new_n745_));
  NA3        g723(.A(new_new_n745_), .B(new_new_n448_), .C(new_new_n365_), .Y(new_new_n746_));
  OAI210     g724(.A0(new_new_n624_), .A1(new_new_n525_), .B0(new_new_n524_), .Y(new_new_n747_));
  NA2        g725(.A(new_new_n747_), .B(new_new_n746_), .Y(new_new_n748_));
  OR3        g726(.A(new_new_n748_), .B(new_new_n744_), .C(new_new_n741_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n632_), .B(i_2_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n751_));
  OAI210     g729(.A0(new_new_n751_), .A1(new_new_n385_), .B0(new_new_n341_), .Y(new_new_n752_));
  NA2        g730(.A(new_new_n752_), .B(new_new_n750_), .Y(new_new_n753_));
  AO210      g731(.A0(new_new_n340_), .A1(new_new_n331_), .B0(new_new_n373_), .Y(new_new_n754_));
  NA3        g732(.A(new_new_n754_), .B(new_new_n243_), .C(i_7_), .Y(new_new_n755_));
  OR2        g733(.A(new_new_n574_), .B(new_new_n421_), .Y(new_new_n756_));
  NA3        g734(.A(new_new_n756_), .B(new_new_n138_), .C(new_new_n61_), .Y(new_new_n757_));
  AO210      g735(.A0(new_new_n463_), .A1(new_new_n684_), .B0(new_new_n36_), .Y(new_new_n758_));
  NA4        g736(.A(new_new_n758_), .B(new_new_n757_), .C(new_new_n755_), .D(new_new_n753_), .Y(new_new_n759_));
  OAI210     g737(.A0(new_new_n588_), .A1(i_11_), .B0(new_new_n77_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n760_), .B(new_new_n524_), .Y(new_new_n761_));
  NA2        g739(.A(new_new_n373_), .B(new_new_n62_), .Y(new_new_n762_));
  NA3        g740(.A(new_new_n762_), .B(new_new_n761_), .C(new_new_n558_), .Y(new_new_n763_));
  AO210      g741(.A0(new_new_n483_), .A1(new_new_n46_), .B0(new_new_n78_), .Y(new_new_n764_));
  NA3        g742(.A(new_new_n764_), .B(new_new_n453_), .C(new_new_n207_), .Y(new_new_n765_));
  AOI210     g743(.A0(new_new_n421_), .A1(new_new_n419_), .B0(new_new_n523_), .Y(new_new_n766_));
  NA2        g744(.A(new_new_n103_), .B(new_new_n383_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n232_), .B(new_new_n46_), .Y(new_new_n768_));
  NA3        g746(.A(new_new_n767_), .B(new_new_n766_), .C(new_new_n765_), .Y(new_new_n769_));
  NO4        g747(.A(new_new_n769_), .B(new_new_n763_), .C(new_new_n759_), .D(new_new_n749_), .Y(new_new_n770_));
  NA4        g748(.A(new_new_n770_), .B(new_new_n736_), .C(new_new_n729_), .D(new_new_n355_), .Y(mai3));
  NA2        g749(.A(i_6_), .B(i_7_), .Y(new_new_n772_));
  NO2        g750(.A(new_new_n772_), .B(i_0_), .Y(new_new_n773_));
  NO2        g751(.A(i_11_), .B(new_new_n224_), .Y(new_new_n774_));
  OAI210     g752(.A0(new_new_n773_), .A1(new_new_n273_), .B0(new_new_n774_), .Y(new_new_n775_));
  INV        g753(.A(new_new_n775_), .Y(new_new_n776_));
  NO3        g754(.A(new_new_n424_), .B(new_new_n82_), .C(new_new_n44_), .Y(new_new_n777_));
  OA210      g755(.A0(new_new_n777_), .A1(new_new_n776_), .B0(new_new_n164_), .Y(new_new_n778_));
  NA2        g756(.A(new_new_n386_), .B(new_new_n45_), .Y(new_new_n779_));
  NO4        g757(.A(new_new_n351_), .B(new_new_n358_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n780_));
  INV        g758(.A(new_new_n780_), .Y(new_new_n781_));
  NA2        g759(.A(new_new_n645_), .B(new_new_n617_), .Y(new_new_n782_));
  NA2        g760(.A(i_0_), .B(i_5_), .Y(new_new_n783_));
  OAI220     g761(.A0(new_new_n783_), .A1(new_new_n782_), .B0(new_new_n781_), .B1(new_new_n58_), .Y(new_new_n784_));
  NO2        g762(.A(new_new_n165_), .B(new_new_n139_), .Y(new_new_n785_));
  NA2        g763(.A(new_new_n785_), .B(new_new_n232_), .Y(new_new_n786_));
  NO2        g764(.A(new_new_n786_), .B(new_new_n965_), .Y(new_new_n787_));
  NO3        g765(.A(new_new_n787_), .B(new_new_n784_), .C(new_new_n778_), .Y(new_new_n788_));
  NA2        g766(.A(new_new_n174_), .B(new_new_n24_), .Y(new_new_n789_));
  NO2        g767(.A(new_new_n615_), .B(new_new_n550_), .Y(new_new_n790_));
  NO2        g768(.A(new_new_n790_), .B(new_new_n789_), .Y(new_new_n791_));
  NA2        g769(.A(new_new_n296_), .B(new_new_n121_), .Y(new_new_n792_));
  OAI220     g770(.A0(new_new_n152_), .A1(new_new_n768_), .B0(new_new_n792_), .B1(new_new_n376_), .Y(new_new_n793_));
  NO2        g771(.A(new_new_n793_), .B(new_new_n791_), .Y(new_new_n794_));
  NO2        g772(.A(new_new_n365_), .B(new_new_n277_), .Y(new_new_n795_));
  NA2        g773(.A(new_new_n795_), .B(new_new_n648_), .Y(new_new_n796_));
  INV        g774(.A(new_new_n448_), .Y(new_new_n797_));
  AN2        g775(.A(new_new_n88_), .B(new_new_n231_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n680_), .B(new_new_n311_), .Y(new_new_n799_));
  INV        g777(.A(new_new_n55_), .Y(new_new_n800_));
  OAI220     g778(.A0(new_new_n800_), .A1(new_new_n799_), .B0(new_new_n606_), .B1(new_new_n499_), .Y(new_new_n801_));
  NO2        g779(.A(new_new_n242_), .B(new_new_n143_), .Y(new_new_n802_));
  NA2        g780(.A(i_0_), .B(i_10_), .Y(new_new_n803_));
  AN2        g781(.A(new_new_n802_), .B(i_6_), .Y(new_new_n804_));
  NA2        g782(.A(new_new_n174_), .B(new_new_n74_), .Y(new_new_n805_));
  NA2        g783(.A(new_new_n528_), .B(i_4_), .Y(new_new_n806_));
  NA2        g784(.A(new_new_n177_), .B(new_new_n192_), .Y(new_new_n807_));
  OAI220     g785(.A0(new_new_n807_), .A1(new_new_n799_), .B0(new_new_n806_), .B1(new_new_n805_), .Y(new_new_n808_));
  NO4        g786(.A(new_new_n808_), .B(new_new_n804_), .C(new_new_n801_), .D(new_new_n798_), .Y(new_new_n809_));
  NA3        g787(.A(new_new_n809_), .B(new_new_n796_), .C(new_new_n794_), .Y(new_new_n810_));
  NA2        g788(.A(i_11_), .B(i_9_), .Y(new_new_n811_));
  NO2        g789(.A(new_new_n48_), .B(i_7_), .Y(new_new_n812_));
  NA2        g790(.A(new_new_n370_), .B(new_new_n169_), .Y(new_new_n813_));
  NA2        g791(.A(new_new_n813_), .B(new_new_n150_), .Y(new_new_n814_));
  NO2        g792(.A(new_new_n811_), .B(new_new_n65_), .Y(new_new_n815_));
  NO2        g793(.A(new_new_n165_), .B(i_0_), .Y(new_new_n816_));
  INV        g794(.A(new_new_n816_), .Y(new_new_n817_));
  NA2        g795(.A(new_new_n448_), .B(new_new_n219_), .Y(new_new_n818_));
  NO2        g796(.A(new_new_n818_), .B(new_new_n817_), .Y(new_new_n819_));
  NO2        g797(.A(new_new_n819_), .B(new_new_n814_), .Y(new_new_n820_));
  NA2        g798(.A(new_new_n605_), .B(new_new_n113_), .Y(new_new_n821_));
  NO2        g799(.A(i_6_), .B(new_new_n821_), .Y(new_new_n822_));
  AOI210     g800(.A0(new_new_n420_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n823_));
  NA2        g801(.A(new_new_n161_), .B(new_new_n95_), .Y(new_new_n824_));
  NOi32      g802(.An(new_new_n823_), .Bn(new_new_n177_), .C(new_new_n824_), .Y(new_new_n825_));
  NA2        g803(.A(new_new_n559_), .B(new_new_n311_), .Y(new_new_n826_));
  NO2        g804(.A(new_new_n826_), .B(new_new_n779_), .Y(new_new_n827_));
  NO3        g805(.A(new_new_n827_), .B(new_new_n825_), .C(new_new_n822_), .Y(new_new_n828_));
  NOi21      g806(.An(i_7_), .B(i_5_), .Y(new_new_n829_));
  NOi31      g807(.An(new_new_n829_), .B(i_0_), .C(new_new_n659_), .Y(new_new_n830_));
  NO3        g808(.A(new_new_n378_), .B(new_new_n343_), .C(new_new_n339_), .Y(new_new_n831_));
  NO2        g809(.A(new_new_n244_), .B(new_new_n300_), .Y(new_new_n832_));
  INV        g810(.A(new_new_n659_), .Y(new_new_n833_));
  AOI210     g811(.A0(new_new_n833_), .A1(new_new_n832_), .B0(new_new_n831_), .Y(new_new_n834_));
  NA3        g812(.A(new_new_n834_), .B(new_new_n828_), .C(new_new_n820_), .Y(new_new_n835_));
  NO2        g813(.A(new_new_n789_), .B(new_new_n227_), .Y(new_new_n836_));
  AN2        g814(.A(new_new_n315_), .B(new_new_n311_), .Y(new_new_n837_));
  AN2        g815(.A(new_new_n837_), .B(new_new_n785_), .Y(new_new_n838_));
  OAI210     g816(.A0(new_new_n838_), .A1(new_new_n836_), .B0(i_10_), .Y(new_new_n839_));
  NA3        g817(.A(new_new_n447_), .B(new_new_n386_), .C(new_new_n45_), .Y(new_new_n840_));
  OAI210     g818(.A0(new_new_n152_), .A1(new_new_n797_), .B0(new_new_n840_), .Y(new_new_n841_));
  NO2        g819(.A(new_new_n243_), .B(new_new_n46_), .Y(new_new_n842_));
  NA2        g820(.A(new_new_n815_), .B(new_new_n289_), .Y(new_new_n843_));
  OAI210     g821(.A0(new_new_n842_), .A1(new_new_n176_), .B0(new_new_n843_), .Y(new_new_n844_));
  AOI220     g822(.A0(new_new_n844_), .A1(new_new_n448_), .B0(new_new_n841_), .B1(new_new_n65_), .Y(new_new_n845_));
  NA3        g823(.A(new_new_n751_), .B(new_new_n357_), .C(new_new_n588_), .Y(new_new_n846_));
  NA2        g824(.A(new_new_n85_), .B(new_new_n44_), .Y(new_new_n847_));
  NO2        g825(.A(new_new_n67_), .B(new_new_n682_), .Y(new_new_n848_));
  AOI220     g826(.A0(new_new_n848_), .A1(new_new_n847_), .B0(new_new_n164_), .B1(new_new_n550_), .Y(new_new_n849_));
  AOI210     g827(.A0(new_new_n849_), .A1(new_new_n846_), .B0(new_new_n47_), .Y(new_new_n850_));
  NO3        g828(.A(i_5_), .B(new_new_n338_), .C(new_new_n24_), .Y(new_new_n851_));
  AOI210     g829(.A0(new_new_n638_), .A1(new_new_n509_), .B0(new_new_n851_), .Y(new_new_n852_));
  NAi21      g830(.An(i_9_), .B(i_5_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n553_), .B(new_new_n97_), .Y(new_new_n854_));
  NA2        g832(.A(new_new_n854_), .B(i_0_), .Y(new_new_n855_));
  OAI220     g833(.A0(new_new_n855_), .A1(new_new_n76_), .B0(new_new_n852_), .B1(new_new_n162_), .Y(new_new_n856_));
  NO3        g834(.A(new_new_n856_), .B(new_new_n850_), .C(new_new_n394_), .Y(new_new_n857_));
  NA3        g835(.A(new_new_n857_), .B(new_new_n845_), .C(new_new_n839_), .Y(new_new_n858_));
  NO3        g836(.A(new_new_n858_), .B(new_new_n835_), .C(new_new_n810_), .Y(new_new_n859_));
  NO2        g837(.A(i_0_), .B(new_new_n659_), .Y(new_new_n860_));
  NO3        g838(.A(new_new_n97_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n861_));
  AO220      g839(.A0(new_new_n861_), .A1(new_new_n44_), .B0(new_new_n860_), .B1(new_new_n164_), .Y(new_new_n862_));
  NO2        g840(.A(new_new_n731_), .B(new_new_n824_), .Y(new_new_n863_));
  AOI210     g841(.A0(new_new_n862_), .A1(new_new_n329_), .B0(new_new_n863_), .Y(new_new_n864_));
  NA3        g842(.A(new_new_n137_), .B(new_new_n617_), .C(new_new_n65_), .Y(new_new_n865_));
  NO2        g843(.A(new_new_n747_), .B(new_new_n378_), .Y(new_new_n866_));
  NA3        g844(.A(new_new_n773_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n867_));
  NA2        g845(.A(new_new_n774_), .B(i_9_), .Y(new_new_n868_));
  AOI210     g846(.A0(new_new_n867_), .A1(new_new_n466_), .B0(new_new_n868_), .Y(new_new_n869_));
  NO2        g847(.A(new_new_n869_), .B(new_new_n866_), .Y(new_new_n870_));
  NA3        g848(.A(new_new_n870_), .B(new_new_n865_), .C(new_new_n864_), .Y(new_new_n871_));
  NA2        g849(.A(new_new_n837_), .B(new_new_n349_), .Y(new_new_n872_));
  AOI210     g850(.A0(new_new_n284_), .A1(new_new_n152_), .B0(new_new_n872_), .Y(new_new_n873_));
  NA3        g851(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n874_));
  NA2        g852(.A(new_new_n812_), .B(new_new_n457_), .Y(new_new_n875_));
  AOI210     g853(.A0(new_new_n874_), .A1(new_new_n152_), .B0(new_new_n875_), .Y(new_new_n876_));
  NO2        g854(.A(new_new_n876_), .B(new_new_n873_), .Y(new_new_n877_));
  NO2        g855(.A(new_new_n803_), .B(new_new_n179_), .Y(new_new_n878_));
  AOI220     g856(.A0(new_new_n878_), .A1(i_11_), .B0(new_new_n529_), .B1(new_new_n67_), .Y(new_new_n879_));
  NO3        g857(.A(new_new_n199_), .B(new_new_n358_), .C(i_0_), .Y(new_new_n880_));
  OAI210     g858(.A0(new_new_n880_), .A1(new_new_n68_), .B0(i_13_), .Y(new_new_n881_));
  INV        g859(.A(new_new_n207_), .Y(new_new_n882_));
  NO2        g860(.A(new_new_n593_), .B(new_new_n568_), .Y(new_new_n883_));
  NA2        g861(.A(new_new_n883_), .B(new_new_n882_), .Y(new_new_n884_));
  NA4        g862(.A(new_new_n884_), .B(new_new_n881_), .C(new_new_n879_), .D(new_new_n877_), .Y(new_new_n885_));
  NA2        g863(.A(new_new_n829_), .B(new_new_n457_), .Y(new_new_n886_));
  INV        g864(.A(new_new_n166_), .Y(new_new_n887_));
  OR2        g865(.A(new_new_n887_), .B(new_new_n886_), .Y(new_new_n888_));
  AOI210     g866(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n165_), .Y(new_new_n889_));
  NA3        g867(.A(new_new_n565_), .B(new_new_n174_), .C(new_new_n74_), .Y(new_new_n890_));
  NA2        g868(.A(new_new_n890_), .B(new_new_n507_), .Y(new_new_n891_));
  NO3        g869(.A(new_new_n779_), .B(new_new_n53_), .C(new_new_n48_), .Y(new_new_n892_));
  INV        g870(.A(new_new_n462_), .Y(new_new_n893_));
  NO3        g871(.A(new_new_n893_), .B(new_new_n892_), .C(new_new_n891_), .Y(new_new_n894_));
  NA3        g872(.A(new_new_n812_), .B(new_new_n273_), .C(new_new_n218_), .Y(new_new_n895_));
  INV        g873(.A(new_new_n895_), .Y(new_new_n896_));
  NA3        g874(.A(new_new_n365_), .B(new_new_n316_), .C(new_new_n210_), .Y(new_new_n897_));
  INV        g875(.A(new_new_n897_), .Y(new_new_n898_));
  NO3        g876(.A(new_new_n811_), .B(new_new_n207_), .C(new_new_n179_), .Y(new_new_n899_));
  NO3        g877(.A(new_new_n899_), .B(new_new_n898_), .C(new_new_n896_), .Y(new_new_n900_));
  NA3        g878(.A(new_new_n900_), .B(new_new_n894_), .C(new_new_n888_), .Y(new_new_n901_));
  INV        g879(.A(new_new_n567_), .Y(new_new_n902_));
  NO3        g880(.A(new_new_n902_), .B(new_new_n519_), .C(new_new_n327_), .Y(new_new_n903_));
  INV        g881(.A(new_new_n903_), .Y(new_new_n904_));
  NA3        g882(.A(new_new_n289_), .B(i_5_), .C(new_new_n182_), .Y(new_new_n905_));
  NA2        g883(.A(new_new_n905_), .B(new_new_n230_), .Y(new_new_n906_));
  NO4        g884(.A(new_new_n227_), .B(new_new_n199_), .C(i_0_), .D(i_12_), .Y(new_new_n907_));
  AOI220     g885(.A0(new_new_n907_), .A1(new_new_n906_), .B0(new_new_n726_), .B1(new_new_n166_), .Y(new_new_n908_));
  AN2        g886(.A(new_new_n803_), .B(new_new_n143_), .Y(new_new_n909_));
  NO4        g887(.A(new_new_n909_), .B(i_12_), .C(new_new_n595_), .D(new_new_n123_), .Y(new_new_n910_));
  NA2        g888(.A(new_new_n910_), .B(new_new_n207_), .Y(new_new_n911_));
  NA3        g889(.A(new_new_n90_), .B(new_new_n533_), .C(i_11_), .Y(new_new_n912_));
  NO2        g890(.A(new_new_n912_), .B(new_new_n145_), .Y(new_new_n913_));
  NA2        g891(.A(new_new_n829_), .B(new_new_n445_), .Y(new_new_n914_));
  OAI220     g892(.A0(i_7_), .A1(new_new_n905_), .B0(new_new_n914_), .B1(new_new_n618_), .Y(new_new_n915_));
  AOI210     g893(.A0(new_new_n915_), .A1(new_new_n816_), .B0(new_new_n913_), .Y(new_new_n916_));
  NA4        g894(.A(new_new_n916_), .B(new_new_n911_), .C(new_new_n908_), .D(new_new_n904_), .Y(new_new_n917_));
  NO4        g895(.A(new_new_n917_), .B(new_new_n901_), .C(new_new_n885_), .D(new_new_n871_), .Y(new_new_n918_));
  OAI210     g896(.A0(new_new_n750_), .A1(new_new_n745_), .B0(new_new_n37_), .Y(new_new_n919_));
  NA3        g897(.A(new_new_n823_), .B(new_new_n347_), .C(i_5_), .Y(new_new_n920_));
  NA3        g898(.A(new_new_n920_), .B(new_new_n919_), .C(new_new_n563_), .Y(new_new_n921_));
  NA2        g899(.A(new_new_n921_), .B(new_new_n196_), .Y(new_new_n922_));
  NA2        g900(.A(new_new_n175_), .B(new_new_n177_), .Y(new_new_n923_));
  AO210      g901(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n923_), .Y(new_new_n924_));
  OAI210     g902(.A0(new_new_n567_), .A1(new_new_n565_), .B0(new_new_n299_), .Y(new_new_n925_));
  NAi31      g903(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n926_));
  NO2        g904(.A(new_new_n62_), .B(new_new_n926_), .Y(new_new_n927_));
  INV        g905(.A(new_new_n927_), .Y(new_new_n928_));
  NA3        g906(.A(new_new_n928_), .B(new_new_n925_), .C(new_new_n924_), .Y(new_new_n929_));
  NO2        g907(.A(new_new_n436_), .B(new_new_n250_), .Y(new_new_n930_));
  NO4        g908(.A(new_new_n221_), .B(new_new_n136_), .C(new_new_n621_), .D(new_new_n37_), .Y(new_new_n931_));
  NO2        g909(.A(new_new_n931_), .B(new_new_n930_), .Y(new_new_n932_));
  OAI210     g910(.A0(new_new_n912_), .A1(new_new_n139_), .B0(new_new_n932_), .Y(new_new_n933_));
  AOI210     g911(.A0(new_new_n929_), .A1(new_new_n48_), .B0(new_new_n933_), .Y(new_new_n934_));
  AOI210     g912(.A0(new_new_n934_), .A1(new_new_n922_), .B0(new_new_n65_), .Y(new_new_n935_));
  NO2        g913(.A(new_new_n526_), .B(new_new_n354_), .Y(new_new_n936_));
  NO2        g914(.A(new_new_n936_), .B(new_new_n688_), .Y(new_new_n937_));
  INV        g915(.A(new_new_n100_), .Y(new_new_n938_));
  NA2        g916(.A(new_new_n938_), .B(new_new_n68_), .Y(new_new_n939_));
  AOI210     g917(.A0(new_new_n889_), .A1(new_new_n812_), .B0(new_new_n830_), .Y(new_new_n940_));
  AOI210     g918(.A0(new_new_n940_), .A1(new_new_n939_), .B0(new_new_n621_), .Y(new_new_n941_));
  INV        g919(.A(new_new_n244_), .Y(new_new_n942_));
  NA2        g920(.A(new_new_n942_), .B(new_new_n68_), .Y(new_new_n943_));
  NO2        g921(.A(new_new_n943_), .B(new_new_n224_), .Y(new_new_n944_));
  NA3        g922(.A(new_new_n88_), .B(new_new_n291_), .C(new_new_n31_), .Y(new_new_n945_));
  INV        g923(.A(new_new_n945_), .Y(new_new_n946_));
  NO3        g924(.A(new_new_n946_), .B(new_new_n944_), .C(new_new_n941_), .Y(new_new_n947_));
  OAI210     g925(.A0(new_new_n252_), .A1(new_new_n148_), .B0(new_new_n79_), .Y(new_new_n948_));
  NA3        g926(.A(new_new_n692_), .B(new_new_n273_), .C(new_new_n72_), .Y(new_new_n949_));
  AOI210     g927(.A0(new_new_n949_), .A1(new_new_n948_), .B0(i_11_), .Y(new_new_n950_));
  INV        g928(.A(new_new_n196_), .Y(new_new_n951_));
  NA2        g929(.A(new_new_n154_), .B(i_5_), .Y(new_new_n952_));
  NO2        g930(.A(new_new_n951_), .B(new_new_n952_), .Y(new_new_n953_));
  NO3        g931(.A(new_new_n853_), .B(i_11_), .C(new_new_n241_), .Y(new_new_n954_));
  NO2        g932(.A(new_new_n954_), .B(new_new_n523_), .Y(new_new_n955_));
  INV        g933(.A(new_new_n344_), .Y(new_new_n956_));
  AOI210     g934(.A0(new_new_n956_), .A1(new_new_n955_), .B0(new_new_n41_), .Y(new_new_n957_));
  NO3        g935(.A(new_new_n957_), .B(new_new_n953_), .C(new_new_n950_), .Y(new_new_n958_));
  OAI210     g936(.A0(new_new_n947_), .A1(i_4_), .B0(new_new_n958_), .Y(new_new_n959_));
  NO3        g937(.A(new_new_n959_), .B(new_new_n937_), .C(new_new_n935_), .Y(new_new_n960_));
  NA4        g938(.A(new_new_n960_), .B(new_new_n918_), .C(new_new_n859_), .D(new_new_n788_), .Y(mai4));
  INV        g939(.A(i_2_), .Y(new_new_n964_));
  INV        g940(.A(i_5_), .Y(new_new_n965_));
  INV        g941(.A(i_0_), .Y(new_new_n966_));
  INV        g942(.A(new_new_n187_), .Y(new_new_n967_));
endmodule


