//Benchmark atmr_9sym_175_0.125

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n60_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n138_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, ori00, mai00, men00;
  INV        o00(.A(i_3_), .Y(ori_ori_n11_));
  INV        o01(.A(i_6_), .Y(ori_ori_n12_));
  INV        o02(.A(i_5_), .Y(ori_ori_n13_));
  INV        o03(.A(i_0_), .Y(ori_ori_n14_));
  INV        o04(.A(i_4_), .Y(ori_ori_n15_));
  NA2        o05(.A(i_0_), .B(ori_ori_n15_), .Y(ori_ori_n16_));
  INV        o06(.A(i_5_), .Y(ori_ori_n17_));
  NO2        o07(.A(ori_ori_n17_), .B(ori_ori_n16_), .Y(ori_ori_n18_));
  NA2        o08(.A(ori_ori_n18_), .B(ori_ori_n11_), .Y(ori_ori_n19_));
  NA2        o09(.A(ori_ori_n14_), .B(i_5_), .Y(ori_ori_n20_));
  INV        o10(.A(i_2_), .Y(ori_ori_n21_));
  NA3        o11(.A(ori_ori_n21_), .B(i_6_), .C(i_8_), .Y(ori_ori_n22_));
  AOI210     o12(.A0(ori_ori_n20_), .A1(i_5_), .B0(ori_ori_n22_), .Y(ori_ori_n23_));
  INV        o13(.A(i_2_), .Y(ori_ori_n24_));
  NO3        o14(.A(i_0_), .B(ori_ori_n24_), .C(i_4_), .Y(ori_ori_n25_));
  NO2        o15(.A(ori_ori_n25_), .B(ori_ori_n23_), .Y(ori_ori_n26_));
  NA2        o16(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n27_));
  NOi21      o17(.An(i_4_), .B(i_3_), .Y(ori_ori_n28_));
  AN2        o18(.A(i_8_), .B(i_7_), .Y(ori_ori_n29_));
  NA2        o19(.A(ori_ori_n28_), .B(i_6_), .Y(ori_ori_n30_));
  INV        o20(.A(ori_ori_n30_), .Y(ori_ori_n31_));
  NA2        o21(.A(ori_ori_n31_), .B(ori_ori_n24_), .Y(ori_ori_n32_));
  NA4        o22(.A(ori_ori_n32_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n19_), .Y(ori_ori_n33_));
  NA2        o23(.A(i_2_), .B(ori_ori_n13_), .Y(ori_ori_n34_));
  NA2        o24(.A(i_2_), .B(ori_ori_n12_), .Y(ori_ori_n35_));
  NA2        o25(.A(ori_ori_n35_), .B(ori_ori_n34_), .Y(ori_ori_n36_));
  NA2        o26(.A(ori_ori_n24_), .B(i_3_), .Y(ori_ori_n37_));
  NO2        o27(.A(ori_ori_n16_), .B(ori_ori_n37_), .Y(ori_ori_n38_));
  NOi21      o28(.An(i_4_), .B(i_6_), .Y(ori_ori_n39_));
  INV        o29(.A(ori_ori_n38_), .Y(ori_ori_n40_));
  NOi21      o30(.An(i_3_), .B(i_1_), .Y(ori_ori_n41_));
  NA2        o31(.A(ori_ori_n41_), .B(i_4_), .Y(ori_ori_n42_));
  AOI210     o32(.A0(i_8_), .A1(i_7_), .B0(ori_ori_n42_), .Y(ori_ori_n43_));
  INV        o33(.A(ori_ori_n43_), .Y(ori_ori_n44_));
  NA2        o34(.A(ori_ori_n44_), .B(ori_ori_n40_), .Y(ori_ori_n45_));
  NO2        o35(.A(i_3_), .B(ori_ori_n20_), .Y(ori_ori_n46_));
  NA2        o36(.A(ori_ori_n29_), .B(ori_ori_n12_), .Y(ori_ori_n47_));
  INV        o37(.A(ori_ori_n47_), .Y(ori_ori_n48_));
  BUFFER     o38(.A(i_0_), .Y(ori_ori_n49_));
  NO2        o39(.A(ori_ori_n48_), .B(ori_ori_n46_), .Y(ori_ori_n50_));
  NO2        o40(.A(i_8_), .B(i_7_), .Y(ori_ori_n51_));
  AN2        o41(.A(i_2_), .B(ori_ori_n51_), .Y(ori_ori_n52_));
  NA2        o42(.A(ori_ori_n49_), .B(ori_ori_n39_), .Y(ori_ori_n53_));
  OAI210     o43(.A0(ori_ori_n37_), .A1(ori_ori_n20_), .B0(ori_ori_n53_), .Y(ori_ori_n54_));
  INV        o44(.A(ori_ori_n54_), .Y(ori_ori_n55_));
  NA3        o45(.A(ori_ori_n55_), .B(ori_ori_n60_), .C(ori_ori_n50_), .Y(ori_ori_n56_));
  OR4        o46(.A(ori_ori_n56_), .B(ori_ori_n45_), .C(ori_ori_n36_), .D(ori_ori_n33_), .Y(ori00));
  INV        o47(.A(ori_ori_n52_), .Y(ori_ori_n60_));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  INV        m002(.A(i_5_), .Y(mai_mai_n13_));
  NOi21      m003(.An(i_3_), .B(i_7_), .Y(mai_mai_n14_));
  INV        m004(.A(i_0_), .Y(mai_mai_n15_));
  NOi21      m005(.An(i_1_), .B(i_3_), .Y(mai_mai_n16_));
  INV        m006(.A(i_4_), .Y(mai_mai_n17_));
  NA2        m007(.A(i_0_), .B(mai_mai_n17_), .Y(mai_mai_n18_));
  INV        m008(.A(i_7_), .Y(mai_mai_n19_));
  NA3        m009(.A(i_6_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n20_));
  NOi21      m010(.An(i_8_), .B(i_6_), .Y(mai_mai_n21_));
  NA2        m011(.A(mai_mai_n21_), .B(i_5_), .Y(mai_mai_n22_));
  AOI210     m012(.A0(mai_mai_n22_), .A1(mai_mai_n20_), .B0(mai_mai_n18_), .Y(mai_mai_n23_));
  NA2        m013(.A(mai_mai_n23_), .B(mai_mai_n11_), .Y(mai_mai_n24_));
  INV        m014(.A(i_2_), .Y(mai_mai_n25_));
  NOi21      m015(.An(i_5_), .B(i_0_), .Y(mai_mai_n26_));
  NOi21      m016(.An(i_6_), .B(i_8_), .Y(mai_mai_n27_));
  NOi21      m017(.An(i_7_), .B(i_1_), .Y(mai_mai_n28_));
  NOi21      m018(.An(i_5_), .B(i_6_), .Y(mai_mai_n29_));
  AOI220     m019(.A0(mai_mai_n29_), .A1(mai_mai_n28_), .B0(mai_mai_n27_), .B1(mai_mai_n26_), .Y(mai_mai_n30_));
  NO3        m020(.A(mai_mai_n30_), .B(mai_mai_n25_), .C(i_4_), .Y(mai_mai_n31_));
  NOi21      m021(.An(i_0_), .B(i_4_), .Y(mai_mai_n32_));
  XO2        m022(.A(i_1_), .B(i_3_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_7_), .B(i_5_), .Y(mai_mai_n34_));
  AN3        m024(.A(mai_mai_n34_), .B(mai_mai_n33_), .C(mai_mai_n32_), .Y(mai_mai_n35_));
  INV        m025(.A(i_1_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_3_), .B(i_0_), .Y(mai_mai_n37_));
  NA2        m027(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  AOI210     m028(.A0(mai_mai_n138_), .A1(mai_mai_n20_), .B0(mai_mai_n38_), .Y(mai_mai_n39_));
  NO3        m029(.A(mai_mai_n39_), .B(mai_mai_n35_), .C(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m030(.A(i_8_), .Y(mai_mai_n41_));
  NOi21      m031(.An(i_4_), .B(i_0_), .Y(mai_mai_n42_));
  AOI210     m032(.A0(mai_mai_n42_), .A1(mai_mai_n21_), .B0(mai_mai_n14_), .Y(mai_mai_n43_));
  NA2        m033(.A(i_1_), .B(mai_mai_n13_), .Y(mai_mai_n44_));
  NOi21      m034(.An(i_2_), .B(i_8_), .Y(mai_mai_n45_));
  NO3        m035(.A(mai_mai_n45_), .B(mai_mai_n42_), .C(mai_mai_n32_), .Y(mai_mai_n46_));
  NO3        m036(.A(mai_mai_n46_), .B(mai_mai_n44_), .C(mai_mai_n43_), .Y(mai_mai_n47_));
  INV        m037(.A(mai_mai_n47_), .Y(mai_mai_n48_));
  NOi31      m038(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n49_));
  NOi21      m039(.An(i_4_), .B(i_3_), .Y(mai_mai_n50_));
  NOi21      m040(.An(i_1_), .B(i_4_), .Y(mai_mai_n51_));
  OAI210     m041(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(mai_mai_n45_), .Y(mai_mai_n52_));
  INV        m042(.A(mai_mai_n52_), .Y(mai_mai_n53_));
  AN2        m043(.A(i_8_), .B(i_7_), .Y(mai_mai_n54_));
  NA2        m044(.A(mai_mai_n54_), .B(mai_mai_n12_), .Y(mai_mai_n55_));
  NOi21      m045(.An(i_8_), .B(i_7_), .Y(mai_mai_n56_));
  NO2        m046(.A(mai_mai_n55_), .B(mai_mai_n44_), .Y(mai_mai_n57_));
  AOI220     m047(.A0(mai_mai_n57_), .A1(mai_mai_n25_), .B0(mai_mai_n53_), .B1(mai_mai_n29_), .Y(mai_mai_n58_));
  NA4        m048(.A(mai_mai_n58_), .B(mai_mai_n48_), .C(mai_mai_n40_), .D(mai_mai_n24_), .Y(mai_mai_n59_));
  NA2        m049(.A(i_8_), .B(mai_mai_n19_), .Y(mai_mai_n60_));
  AOI220     m050(.A0(mai_mai_n37_), .A1(i_1_), .B0(mai_mai_n33_), .B1(i_2_), .Y(mai_mai_n61_));
  NOi21      m051(.An(i_1_), .B(i_2_), .Y(mai_mai_n62_));
  NA3        m052(.A(mai_mai_n62_), .B(mai_mai_n42_), .C(i_6_), .Y(mai_mai_n63_));
  OAI210     m053(.A0(mai_mai_n61_), .A1(mai_mai_n60_), .B0(mai_mai_n63_), .Y(mai_mai_n64_));
  NA2        m054(.A(mai_mai_n64_), .B(mai_mai_n13_), .Y(mai_mai_n65_));
  NOi32      m055(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n66_));
  NA2        m056(.A(mai_mai_n66_), .B(i_3_), .Y(mai_mai_n67_));
  NA3        m057(.A(mai_mai_n16_), .B(i_2_), .C(i_6_), .Y(mai_mai_n68_));
  NA2        m058(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  NO2        m059(.A(i_0_), .B(i_4_), .Y(mai_mai_n70_));
  AOI220     m060(.A0(mai_mai_n70_), .A1(mai_mai_n69_), .B0(mai_mai_n56_), .B1(mai_mai_n50_), .Y(mai_mai_n71_));
  NA2        m061(.A(mai_mai_n71_), .B(mai_mai_n65_), .Y(mai_mai_n72_));
  NAi21      m062(.An(i_3_), .B(i_6_), .Y(mai_mai_n73_));
  NO3        m063(.A(mai_mai_n73_), .B(i_0_), .C(mai_mai_n41_), .Y(mai_mai_n74_));
  NA2        m064(.A(mai_mai_n27_), .B(mai_mai_n26_), .Y(mai_mai_n75_));
  NOi21      m065(.An(i_7_), .B(i_8_), .Y(mai_mai_n76_));
  NOi31      m066(.An(i_6_), .B(i_5_), .C(i_7_), .Y(mai_mai_n77_));
  AOI210     m067(.A0(mai_mai_n76_), .A1(mai_mai_n12_), .B0(mai_mai_n77_), .Y(mai_mai_n78_));
  OAI210     m068(.A0(mai_mai_n78_), .A1(mai_mai_n11_), .B0(mai_mai_n75_), .Y(mai_mai_n79_));
  OAI210     m069(.A0(mai_mai_n79_), .A1(mai_mai_n74_), .B0(mai_mai_n62_), .Y(mai_mai_n80_));
  NA3        m070(.A(mai_mai_n56_), .B(mai_mai_n25_), .C(i_3_), .Y(mai_mai_n81_));
  AOI210     m071(.A0(i_1_), .A1(mai_mai_n18_), .B0(mai_mai_n81_), .Y(mai_mai_n82_));
  NAi21      m072(.An(i_6_), .B(i_0_), .Y(mai_mai_n83_));
  NA3        m073(.A(mai_mai_n51_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n84_));
  NOi21      m074(.An(i_4_), .B(i_6_), .Y(mai_mai_n85_));
  NOi21      m075(.An(i_5_), .B(i_3_), .Y(mai_mai_n86_));
  NA3        m076(.A(mai_mai_n86_), .B(mai_mai_n62_), .C(mai_mai_n85_), .Y(mai_mai_n87_));
  OAI210     m077(.A0(mai_mai_n84_), .A1(mai_mai_n83_), .B0(mai_mai_n87_), .Y(mai_mai_n88_));
  NA2        m078(.A(mai_mai_n62_), .B(mai_mai_n27_), .Y(mai_mai_n89_));
  NOi21      m079(.An(mai_mai_n34_), .B(mai_mai_n89_), .Y(mai_mai_n90_));
  NO3        m080(.A(mai_mai_n90_), .B(mai_mai_n88_), .C(mai_mai_n82_), .Y(mai_mai_n91_));
  NA2        m081(.A(mai_mai_n56_), .B(mai_mai_n12_), .Y(mai_mai_n92_));
  NA2        m082(.A(mai_mai_n27_), .B(mai_mai_n13_), .Y(mai_mai_n93_));
  NOi21      m083(.An(i_3_), .B(i_1_), .Y(mai_mai_n94_));
  NA2        m084(.A(mai_mai_n94_), .B(i_4_), .Y(mai_mai_n95_));
  AOI210     m085(.A0(mai_mai_n93_), .A1(mai_mai_n92_), .B0(mai_mai_n95_), .Y(mai_mai_n96_));
  INV        m086(.A(mai_mai_n96_), .Y(mai_mai_n97_));
  NA3        m087(.A(mai_mai_n97_), .B(mai_mai_n91_), .C(mai_mai_n80_), .Y(mai_mai_n98_));
  NOi31      m088(.An(i_6_), .B(i_1_), .C(i_8_), .Y(mai_mai_n99_));
  NA2        m089(.A(mai_mai_n27_), .B(mai_mai_n32_), .Y(mai_mai_n100_));
  NA3        m090(.A(mai_mai_n56_), .B(mai_mai_n49_), .C(i_6_), .Y(mai_mai_n101_));
  INV        m091(.A(mai_mai_n101_), .Y(mai_mai_n102_));
  NOi21      m092(.An(i_0_), .B(i_2_), .Y(mai_mai_n103_));
  NA3        m093(.A(mai_mai_n103_), .B(mai_mai_n28_), .C(mai_mai_n85_), .Y(mai_mai_n104_));
  NA3        m094(.A(mai_mai_n42_), .B(mai_mai_n34_), .C(mai_mai_n16_), .Y(mai_mai_n105_));
  NOi32      m095(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(mai_mai_n106_));
  NA2        m096(.A(mai_mai_n106_), .B(mai_mai_n99_), .Y(mai_mai_n107_));
  NA3        m097(.A(mai_mai_n103_), .B(mai_mai_n50_), .C(mai_mai_n27_), .Y(mai_mai_n108_));
  NA4        m098(.A(mai_mai_n108_), .B(mai_mai_n107_), .C(mai_mai_n105_), .D(mai_mai_n104_), .Y(mai_mai_n109_));
  NA4        m099(.A(mai_mai_n49_), .B(i_6_), .C(mai_mai_n13_), .D(i_7_), .Y(mai_mai_n110_));
  NA4        m100(.A(mai_mai_n51_), .B(mai_mai_n29_), .C(mai_mai_n15_), .D(i_8_), .Y(mai_mai_n111_));
  NA2        m101(.A(mai_mai_n111_), .B(mai_mai_n110_), .Y(mai_mai_n112_));
  NO3        m102(.A(mai_mai_n112_), .B(mai_mai_n109_), .C(mai_mai_n102_), .Y(mai_mai_n113_));
  NO4        m103(.A(i_2_), .B(mai_mai_n17_), .C(mai_mai_n11_), .D(mai_mai_n13_), .Y(mai_mai_n114_));
  NA2        m104(.A(i_2_), .B(i_4_), .Y(mai_mai_n115_));
  AOI210     m105(.A0(mai_mai_n83_), .A1(mai_mai_n73_), .B0(mai_mai_n115_), .Y(mai_mai_n116_));
  NO2        m106(.A(i_8_), .B(i_7_), .Y(mai_mai_n117_));
  OA210      m107(.A0(mai_mai_n116_), .A1(mai_mai_n114_), .B0(mai_mai_n117_), .Y(mai_mai_n118_));
  NA3        m108(.A(mai_mai_n94_), .B(i_0_), .C(i_5_), .Y(mai_mai_n119_));
  NO2        m109(.A(mai_mai_n119_), .B(i_4_), .Y(mai_mai_n120_));
  NO2        m110(.A(mai_mai_n120_), .B(mai_mai_n118_), .Y(mai_mai_n121_));
  NA2        m111(.A(mai_mai_n76_), .B(mai_mai_n12_), .Y(mai_mai_n122_));
  NA3        m112(.A(i_2_), .B(i_1_), .C(mai_mai_n13_), .Y(mai_mai_n123_));
  INV        m113(.A(mai_mai_n42_), .Y(mai_mai_n124_));
  AOI210     m114(.A0(mai_mai_n124_), .A1(mai_mai_n123_), .B0(mai_mai_n122_), .Y(mai_mai_n125_));
  NA3        m115(.A(mai_mai_n103_), .B(mai_mai_n56_), .C(mai_mai_n85_), .Y(mai_mai_n126_));
  OAI210     m116(.A0(mai_mai_n81_), .A1(i_0_), .B0(mai_mai_n126_), .Y(mai_mai_n127_));
  NA3        m117(.A(mai_mai_n86_), .B(mai_mai_n54_), .C(mai_mai_n36_), .Y(mai_mai_n128_));
  NA3        m118(.A(mai_mai_n45_), .B(mai_mai_n26_), .C(mai_mai_n14_), .Y(mai_mai_n129_));
  NOi31      m119(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n130_));
  OAI210     m120(.A0(mai_mai_n106_), .A1(mai_mai_n66_), .B0(mai_mai_n130_), .Y(mai_mai_n131_));
  NA3        m121(.A(mai_mai_n131_), .B(mai_mai_n129_), .C(mai_mai_n128_), .Y(mai_mai_n132_));
  NO3        m122(.A(mai_mai_n132_), .B(mai_mai_n127_), .C(mai_mai_n125_), .Y(mai_mai_n133_));
  NA4        m123(.A(mai_mai_n133_), .B(mai_mai_n121_), .C(mai_mai_n113_), .D(mai_mai_n100_), .Y(mai_mai_n134_));
  OR4        m124(.A(mai_mai_n134_), .B(mai_mai_n98_), .C(mai_mai_n72_), .D(mai_mai_n59_), .Y(mai00));
  INV        m125(.A(i_7_), .Y(mai_mai_n138_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NA3        u013(.A(i_6_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n24_));
  NOi21      u014(.An(i_8_), .B(i_6_), .Y(men_men_n25_));
  NOi21      u015(.An(i_1_), .B(i_8_), .Y(men_men_n26_));
  AOI220     u016(.A0(men_men_n26_), .A1(i_2_), .B0(men_men_n25_), .B1(i_5_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n22_), .Y(men_men_n28_));
  AOI210     u018(.A0(men_men_n28_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n29_));
  NA2        u019(.A(i_0_), .B(men_men_n14_), .Y(men_men_n30_));
  NA2        u020(.A(men_men_n17_), .B(i_5_), .Y(men_men_n31_));
  NO2        u021(.A(i_2_), .B(i_4_), .Y(men_men_n32_));
  NA3        u022(.A(men_men_n32_), .B(i_6_), .C(i_8_), .Y(men_men_n33_));
  AOI210     u023(.A0(men_men_n31_), .A1(men_men_n30_), .B0(men_men_n33_), .Y(men_men_n34_));
  INV        u024(.A(i_2_), .Y(men_men_n35_));
  NOi21      u025(.An(i_5_), .B(i_0_), .Y(men_men_n36_));
  NOi21      u026(.An(i_6_), .B(i_8_), .Y(men_men_n37_));
  NOi21      u027(.An(i_7_), .B(i_1_), .Y(men_men_n38_));
  NOi21      u028(.An(i_5_), .B(i_6_), .Y(men_men_n39_));
  AOI220     u029(.A0(men_men_n39_), .A1(men_men_n38_), .B0(men_men_n37_), .B1(men_men_n36_), .Y(men_men_n40_));
  NO3        u030(.A(men_men_n40_), .B(men_men_n35_), .C(i_4_), .Y(men_men_n41_));
  NOi21      u031(.An(i_0_), .B(i_4_), .Y(men_men_n42_));
  XO2        u032(.A(i_1_), .B(i_3_), .Y(men_men_n43_));
  NOi21      u033(.An(i_7_), .B(i_5_), .Y(men_men_n44_));
  INV        u034(.A(i_1_), .Y(men_men_n45_));
  NOi21      u035(.An(i_3_), .B(i_0_), .Y(men_men_n46_));
  NA2        u036(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NA3        u037(.A(i_6_), .B(men_men_n14_), .C(i_7_), .Y(men_men_n48_));
  AOI210     u038(.A0(men_men_n48_), .A1(men_men_n24_), .B0(men_men_n47_), .Y(men_men_n49_));
  NO3        u039(.A(men_men_n49_), .B(men_men_n41_), .C(men_men_n34_), .Y(men_men_n50_));
  INV        u040(.A(i_8_), .Y(men_men_n51_));
  NA2        u041(.A(i_1_), .B(men_men_n11_), .Y(men_men_n52_));
  NO4        u042(.A(men_men_n52_), .B(men_men_n30_), .C(i_2_), .D(men_men_n51_), .Y(men_men_n53_));
  NOi21      u043(.An(i_4_), .B(i_0_), .Y(men_men_n54_));
  AOI210     u044(.A0(men_men_n54_), .A1(men_men_n25_), .B0(men_men_n15_), .Y(men_men_n55_));
  NA2        u045(.A(i_1_), .B(men_men_n14_), .Y(men_men_n56_));
  NOi21      u046(.An(i_2_), .B(i_8_), .Y(men_men_n57_));
  NO3        u047(.A(men_men_n57_), .B(men_men_n54_), .C(men_men_n42_), .Y(men_men_n58_));
  NO3        u048(.A(men_men_n58_), .B(men_men_n56_), .C(men_men_n55_), .Y(men_men_n59_));
  NO2        u049(.A(men_men_n59_), .B(men_men_n53_), .Y(men_men_n60_));
  NOi31      u050(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n61_));
  NA2        u051(.A(men_men_n61_), .B(i_0_), .Y(men_men_n62_));
  NOi21      u052(.An(i_4_), .B(i_3_), .Y(men_men_n63_));
  NOi21      u053(.An(i_1_), .B(i_4_), .Y(men_men_n64_));
  OAI210     u054(.A0(men_men_n64_), .A1(men_men_n63_), .B0(men_men_n57_), .Y(men_men_n65_));
  NA2        u055(.A(men_men_n65_), .B(men_men_n62_), .Y(men_men_n66_));
  AN2        u056(.A(i_8_), .B(i_7_), .Y(men_men_n67_));
  NOi21      u057(.An(i_8_), .B(i_7_), .Y(men_men_n68_));
  NA2        u058(.A(men_men_n66_), .B(men_men_n39_), .Y(men_men_n69_));
  NA4        u059(.A(men_men_n69_), .B(men_men_n60_), .C(men_men_n50_), .D(men_men_n29_), .Y(men_men_n70_));
  NA2        u060(.A(i_8_), .B(i_7_), .Y(men_men_n71_));
  NO3        u061(.A(men_men_n71_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n72_));
  NA2        u062(.A(i_8_), .B(men_men_n23_), .Y(men_men_n73_));
  AOI220     u063(.A0(men_men_n46_), .A1(i_1_), .B0(men_men_n43_), .B1(i_2_), .Y(men_men_n74_));
  NOi21      u064(.An(i_1_), .B(i_2_), .Y(men_men_n75_));
  NO2        u065(.A(men_men_n74_), .B(men_men_n73_), .Y(men_men_n76_));
  OAI210     u066(.A0(men_men_n76_), .A1(men_men_n72_), .B0(men_men_n14_), .Y(men_men_n77_));
  NA3        u067(.A(men_men_n68_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n78_));
  NA3        u068(.A(men_men_n26_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n79_));
  NA2        u069(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NA2        u070(.A(men_men_n80_), .B(men_men_n63_), .Y(men_men_n81_));
  NA2        u071(.A(men_men_n81_), .B(men_men_n77_), .Y(men_men_n82_));
  NAi21      u072(.An(i_3_), .B(i_6_), .Y(men_men_n83_));
  NO3        u073(.A(men_men_n83_), .B(i_0_), .C(men_men_n51_), .Y(men_men_n84_));
  NA2        u074(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n85_));
  NOi21      u075(.An(i_7_), .B(i_8_), .Y(men_men_n86_));
  NA2        u076(.A(men_men_n86_), .B(men_men_n12_), .Y(men_men_n87_));
  OAI210     u077(.A0(men_men_n87_), .A1(men_men_n11_), .B0(men_men_n85_), .Y(men_men_n88_));
  OAI210     u078(.A0(men_men_n88_), .A1(men_men_n84_), .B0(men_men_n75_), .Y(men_men_n89_));
  NA3        u079(.A(men_men_n25_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n90_));
  AOI210     u080(.A0(men_men_n22_), .A1(men_men_n52_), .B0(men_men_n90_), .Y(men_men_n91_));
  AOI220     u081(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n18_), .B1(men_men_n35_), .Y(men_men_n92_));
  NA3        u082(.A(men_men_n21_), .B(i_5_), .C(i_7_), .Y(men_men_n93_));
  OAI210     u083(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n94_));
  NA3        u084(.A(men_men_n71_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n95_));
  OAI220     u085(.A0(men_men_n95_), .A1(men_men_n94_), .B0(men_men_n93_), .B1(men_men_n92_), .Y(men_men_n96_));
  NO2        u086(.A(men_men_n96_), .B(men_men_n91_), .Y(men_men_n97_));
  NA2        u087(.A(men_men_n45_), .B(i_6_), .Y(men_men_n98_));
  NOi21      u088(.An(i_2_), .B(i_1_), .Y(men_men_n99_));
  NAi21      u089(.An(i_6_), .B(i_0_), .Y(men_men_n100_));
  NA2        u090(.A(men_men_n75_), .B(men_men_n37_), .Y(men_men_n101_));
  NOi21      u091(.An(men_men_n44_), .B(men_men_n101_), .Y(men_men_n102_));
  INV        u092(.A(men_men_n102_), .Y(men_men_n103_));
  NOi21      u093(.An(i_6_), .B(i_1_), .Y(men_men_n104_));
  AOI220     u094(.A0(men_men_n104_), .A1(i_7_), .B0(men_men_n25_), .B1(i_5_), .Y(men_men_n105_));
  NOi31      u095(.An(men_men_n54_), .B(men_men_n105_), .C(i_2_), .Y(men_men_n106_));
  AOI220     u096(.A0(men_men_n86_), .A1(men_men_n14_), .B0(i_4_), .B1(men_men_n23_), .Y(men_men_n107_));
  NOi31      u097(.An(men_men_n46_), .B(men_men_n107_), .C(men_men_n35_), .Y(men_men_n108_));
  NO2        u098(.A(men_men_n108_), .B(men_men_n106_), .Y(men_men_n109_));
  NA4        u099(.A(men_men_n109_), .B(men_men_n103_), .C(men_men_n97_), .D(men_men_n89_), .Y(men_men_n110_));
  NA2        u100(.A(men_men_n57_), .B(men_men_n15_), .Y(men_men_n111_));
  NOi31      u101(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n112_));
  NOi31      u102(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n113_));
  OAI210     u103(.A0(men_men_n113_), .A1(men_men_n112_), .B0(i_7_), .Y(men_men_n114_));
  NA3        u104(.A(men_men_n114_), .B(men_men_n111_), .C(men_men_n101_), .Y(men_men_n115_));
  NA2        u105(.A(men_men_n115_), .B(men_men_n42_), .Y(men_men_n116_));
  NO2        u106(.A(men_men_n78_), .B(men_men_n31_), .Y(men_men_n117_));
  NA4        u107(.A(men_men_n67_), .B(men_men_n99_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n118_));
  NAi31      u108(.An(men_men_n100_), .B(men_men_n86_), .C(men_men_n99_), .Y(men_men_n119_));
  NA3        u109(.A(men_men_n68_), .B(men_men_n61_), .C(i_6_), .Y(men_men_n120_));
  NA3        u110(.A(men_men_n120_), .B(men_men_n119_), .C(men_men_n118_), .Y(men_men_n121_));
  NOi21      u111(.An(i_0_), .B(i_2_), .Y(men_men_n122_));
  NA2        u112(.A(men_men_n122_), .B(men_men_n38_), .Y(men_men_n123_));
  NA3        u113(.A(men_men_n54_), .B(men_men_n44_), .C(men_men_n18_), .Y(men_men_n124_));
  NOi32      u114(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n125_));
  NA2        u115(.A(men_men_n125_), .B(men_men_n112_), .Y(men_men_n126_));
  NA3        u116(.A(men_men_n126_), .B(men_men_n124_), .C(men_men_n123_), .Y(men_men_n127_));
  NA4        u117(.A(men_men_n61_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n128_));
  NA4        u118(.A(men_men_n64_), .B(men_men_n39_), .C(men_men_n17_), .D(i_8_), .Y(men_men_n129_));
  NA4        u119(.A(men_men_n64_), .B(men_men_n46_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n130_));
  NA3        u120(.A(men_men_n130_), .B(men_men_n129_), .C(men_men_n128_), .Y(men_men_n131_));
  NO4        u121(.A(men_men_n131_), .B(men_men_n127_), .C(men_men_n121_), .D(men_men_n117_), .Y(men_men_n132_));
  NOi21      u122(.An(i_5_), .B(i_2_), .Y(men_men_n133_));
  AOI220     u123(.A0(men_men_n133_), .A1(men_men_n86_), .B0(men_men_n67_), .B1(men_men_n32_), .Y(men_men_n134_));
  AOI210     u124(.A0(men_men_n134_), .A1(men_men_n111_), .B0(men_men_n98_), .Y(men_men_n135_));
  NO4        u125(.A(i_2_), .B(men_men_n21_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n136_));
  NA2        u126(.A(i_2_), .B(i_4_), .Y(men_men_n137_));
  AOI210     u127(.A0(men_men_n100_), .A1(men_men_n83_), .B0(men_men_n137_), .Y(men_men_n138_));
  NO2        u128(.A(i_8_), .B(i_7_), .Y(men_men_n139_));
  OA210      u129(.A0(men_men_n138_), .A1(men_men_n136_), .B0(men_men_n139_), .Y(men_men_n140_));
  NA4        u130(.A(i_3_), .B(i_0_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n141_));
  NO2        u131(.A(men_men_n141_), .B(i_4_), .Y(men_men_n142_));
  NO3        u132(.A(men_men_n142_), .B(men_men_n140_), .C(men_men_n135_), .Y(men_men_n143_));
  NA2        u133(.A(men_men_n122_), .B(men_men_n68_), .Y(men_men_n144_));
  NA4        u134(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n132_), .D(men_men_n116_), .Y(men_men_n145_));
  OR4        u135(.A(men_men_n145_), .B(men_men_n110_), .C(men_men_n82_), .D(men_men_n70_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule