//Benchmark atmr_max1024_476_0.0625

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n444_, mai_mai_n445_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO4        o012(.A(ori_ori_n28_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  AN2        o021(.A(x8), .B(x7), .Y(ori_ori_n38_));
  NA3        o022(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o023(.A(x4), .B(x3), .Y(ori_ori_n40_));
  AOI210     o024(.A0(ori_ori_n39_), .A1(ori_ori_n23_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o025(.A(x2), .B(x0), .Y(ori_ori_n42_));
  INV        o026(.A(x3), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  INV        o028(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n42_), .Y(ori_ori_n47_));
  INV        o031(.A(x4), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(x2), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n50_), .A1(ori_ori_n20_), .B0(ori_ori_n47_), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n52_));
  AOI220     o036(.A0(ori_ori_n52_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n53_));
  INV        o037(.A(x2), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  OAI210     o041(.A0(ori_ori_n53_), .A1(ori_ori_n32_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  NO3        o042(.A(ori_ori_n58_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori01));
  NA2        o043(.A(x8), .B(x7), .Y(ori_ori_n60_));
  NA2        o044(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n61_));
  INV        o045(.A(x9), .Y(ori_ori_n62_));
  NO2        o046(.A(x7), .B(x6), .Y(ori_ori_n63_));
  NO2        o047(.A(ori_ori_n61_), .B(x5), .Y(ori_ori_n64_));
  NO2        o048(.A(x8), .B(x2), .Y(ori_ori_n65_));
  INV        o049(.A(ori_ori_n65_), .Y(ori_ori_n66_));
  NO2        o050(.A(ori_ori_n66_), .B(x1), .Y(ori_ori_n67_));
  OA210      o051(.A0(ori_ori_n67_), .A1(ori_ori_n64_), .B0(ori_ori_n63_), .Y(ori_ori_n68_));
  OAI210     o052(.A0(ori_ori_n44_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n56_), .A1(ori_ori_n20_), .B0(ori_ori_n69_), .Y(ori_ori_n70_));
  NO2        o054(.A(ori_ori_n70_), .B(ori_ori_n68_), .Y(ori_ori_n71_));
  NA2        o055(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n73_));
  OAI210     o057(.A0(ori_ori_n73_), .A1(ori_ori_n56_), .B0(x0), .Y(ori_ori_n74_));
  NA2        o058(.A(x5), .B(x3), .Y(ori_ori_n75_));
  NO2        o059(.A(x8), .B(x6), .Y(ori_ori_n76_));
  NO4        o060(.A(ori_ori_n76_), .B(ori_ori_n75_), .C(ori_ori_n63_), .D(ori_ori_n54_), .Y(ori_ori_n77_));
  NAi21      o061(.An(x4), .B(x3), .Y(ori_ori_n78_));
  INV        o062(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NO2        o063(.A(ori_ori_n79_), .B(ori_ori_n22_), .Y(ori_ori_n80_));
  NO2        o064(.A(x4), .B(x2), .Y(ori_ori_n81_));
  NO2        o065(.A(ori_ori_n81_), .B(x3), .Y(ori_ori_n82_));
  NO3        o066(.A(ori_ori_n82_), .B(ori_ori_n80_), .C(ori_ori_n18_), .Y(ori_ori_n83_));
  NO3        o067(.A(ori_ori_n83_), .B(ori_ori_n77_), .C(ori_ori_n74_), .Y(ori_ori_n84_));
  NA2        o068(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n85_));
  NO2        o069(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n86_));
  INV        o070(.A(x8), .Y(ori_ori_n87_));
  NA2        o071(.A(x2), .B(x1), .Y(ori_ori_n88_));
  INV        o072(.A(ori_ori_n86_), .Y(ori_ori_n89_));
  NO2        o073(.A(ori_ori_n89_), .B(ori_ori_n26_), .Y(ori_ori_n90_));
  AOI210     o074(.A0(ori_ori_n56_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n91_));
  OAI210     o075(.A0(ori_ori_n45_), .A1(ori_ori_n37_), .B0(ori_ori_n48_), .Y(ori_ori_n92_));
  NO3        o076(.A(ori_ori_n92_), .B(ori_ori_n91_), .C(ori_ori_n90_), .Y(ori_ori_n93_));
  NA2        o077(.A(x4), .B(ori_ori_n43_), .Y(ori_ori_n94_));
  NO2        o078(.A(ori_ori_n48_), .B(ori_ori_n54_), .Y(ori_ori_n95_));
  OAI210     o079(.A0(ori_ori_n95_), .A1(ori_ori_n43_), .B0(ori_ori_n18_), .Y(ori_ori_n96_));
  AOI210     o080(.A0(ori_ori_n94_), .A1(ori_ori_n52_), .B0(ori_ori_n96_), .Y(ori_ori_n97_));
  NO2        o081(.A(x3), .B(x2), .Y(ori_ori_n98_));
  NA3        o082(.A(ori_ori_n98_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n99_));
  INV        o083(.A(ori_ori_n99_), .Y(ori_ori_n100_));
  NA2        o084(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n101_));
  OAI210     o085(.A0(ori_ori_n101_), .A1(ori_ori_n40_), .B0(ori_ori_n17_), .Y(ori_ori_n102_));
  NO4        o086(.A(ori_ori_n102_), .B(ori_ori_n100_), .C(ori_ori_n97_), .D(ori_ori_n93_), .Y(ori_ori_n103_));
  AO210      o087(.A0(ori_ori_n84_), .A1(ori_ori_n72_), .B0(ori_ori_n103_), .Y(ori02));
  NO2        o088(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n105_));
  NO2        o089(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n106_));
  NA2        o090(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n107_));
  INV        o091(.A(ori_ori_n107_), .Y(ori_ori_n108_));
  AOI220     o092(.A0(ori_ori_n108_), .A1(ori_ori_n106_), .B0(ori_ori_n105_), .B1(x4), .Y(ori_ori_n109_));
  NO3        o093(.A(ori_ori_n109_), .B(x7), .C(x5), .Y(ori_ori_n110_));
  OR2        o094(.A(x8), .B(x0), .Y(ori_ori_n111_));
  INV        o095(.A(ori_ori_n111_), .Y(ori_ori_n112_));
  NAi21      o096(.An(x2), .B(x8), .Y(ori_ori_n113_));
  NO2        o097(.A(x4), .B(x1), .Y(ori_ori_n114_));
  NA3        o098(.A(ori_ori_n114_), .B(x2), .C(ori_ori_n60_), .Y(ori_ori_n115_));
  NOi21      o099(.An(x0), .B(x1), .Y(ori_ori_n116_));
  NO3        o100(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n117_));
  NOi21      o101(.An(x0), .B(x4), .Y(ori_ori_n118_));
  NAi21      o102(.An(x8), .B(x7), .Y(ori_ori_n119_));
  NO2        o103(.A(ori_ori_n119_), .B(ori_ori_n62_), .Y(ori_ori_n120_));
  AOI220     o104(.A0(ori_ori_n120_), .A1(ori_ori_n118_), .B0(ori_ori_n117_), .B1(ori_ori_n116_), .Y(ori_ori_n121_));
  AOI210     o105(.A0(ori_ori_n121_), .A1(ori_ori_n115_), .B0(ori_ori_n75_), .Y(ori_ori_n122_));
  NO2        o106(.A(x5), .B(ori_ori_n48_), .Y(ori_ori_n123_));
  NA2        o107(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n124_));
  AOI210     o108(.A0(ori_ori_n124_), .A1(ori_ori_n101_), .B0(ori_ori_n107_), .Y(ori_ori_n125_));
  OAI210     o109(.A0(ori_ori_n125_), .A1(ori_ori_n35_), .B0(ori_ori_n123_), .Y(ori_ori_n126_));
  NAi21      o110(.An(x0), .B(x4), .Y(ori_ori_n127_));
  NO2        o111(.A(ori_ori_n127_), .B(x1), .Y(ori_ori_n128_));
  NO2        o112(.A(x7), .B(x0), .Y(ori_ori_n129_));
  NO2        o113(.A(ori_ori_n81_), .B(ori_ori_n95_), .Y(ori_ori_n130_));
  NO2        o114(.A(ori_ori_n130_), .B(x3), .Y(ori_ori_n131_));
  OAI210     o115(.A0(ori_ori_n129_), .A1(ori_ori_n128_), .B0(ori_ori_n131_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n133_));
  NA2        o117(.A(x5), .B(x0), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n135_));
  NA3        o119(.A(ori_ori_n135_), .B(ori_ori_n134_), .C(ori_ori_n133_), .Y(ori_ori_n136_));
  NA4        o120(.A(ori_ori_n136_), .B(ori_ori_n132_), .C(ori_ori_n126_), .D(ori_ori_n36_), .Y(ori_ori_n137_));
  NO3        o121(.A(ori_ori_n137_), .B(ori_ori_n122_), .C(ori_ori_n110_), .Y(ori_ori_n138_));
  NO3        o122(.A(ori_ori_n75_), .B(ori_ori_n73_), .C(ori_ori_n24_), .Y(ori_ori_n139_));
  NO2        o123(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n140_));
  NA2        o124(.A(x7), .B(x3), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n94_), .B(x5), .Y(ori_ori_n142_));
  NO2        o126(.A(x9), .B(x7), .Y(ori_ori_n143_));
  NOi21      o127(.An(x8), .B(x0), .Y(ori_ori_n144_));
  NO2        o128(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n145_));
  INV        o129(.A(x7), .Y(ori_ori_n146_));
  NA2        o130(.A(ori_ori_n146_), .B(ori_ori_n18_), .Y(ori_ori_n147_));
  AOI220     o131(.A0(ori_ori_n147_), .A1(ori_ori_n145_), .B0(ori_ori_n105_), .B1(ori_ori_n38_), .Y(ori_ori_n148_));
  NO2        o132(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n149_));
  NO2        o133(.A(ori_ori_n149_), .B(ori_ori_n118_), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n150_), .B(ori_ori_n148_), .Y(ori_ori_n151_));
  INV        o135(.A(ori_ori_n151_), .Y(ori_ori_n152_));
  OAI210     o136(.A0(ori_ori_n141_), .A1(ori_ori_n50_), .B0(ori_ori_n152_), .Y(ori_ori_n153_));
  NA2        o137(.A(x5), .B(x1), .Y(ori_ori_n154_));
  INV        o138(.A(ori_ori_n154_), .Y(ori_ori_n155_));
  AOI210     o139(.A0(ori_ori_n155_), .A1(ori_ori_n118_), .B0(ori_ori_n36_), .Y(ori_ori_n156_));
  NAi21      o140(.An(x2), .B(x7), .Y(ori_ori_n157_));
  NO2        o141(.A(ori_ori_n157_), .B(ori_ori_n48_), .Y(ori_ori_n158_));
  NA2        o142(.A(ori_ori_n158_), .B(ori_ori_n64_), .Y(ori_ori_n159_));
  NAi31      o143(.An(ori_ori_n75_), .B(ori_ori_n38_), .C(ori_ori_n35_), .Y(ori_ori_n160_));
  NA3        o144(.A(ori_ori_n160_), .B(ori_ori_n159_), .C(ori_ori_n156_), .Y(ori_ori_n161_));
  NO3        o145(.A(ori_ori_n161_), .B(ori_ori_n153_), .C(ori_ori_n139_), .Y(ori_ori_n162_));
  NO2        o146(.A(ori_ori_n162_), .B(ori_ori_n138_), .Y(ori_ori_n163_));
  NO2        o147(.A(ori_ori_n134_), .B(ori_ori_n130_), .Y(ori_ori_n164_));
  NA2        o148(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n165_));
  NA2        o149(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n166_));
  NA3        o150(.A(ori_ori_n166_), .B(ori_ori_n165_), .C(ori_ori_n24_), .Y(ori_ori_n167_));
  AN2        o151(.A(ori_ori_n167_), .B(ori_ori_n135_), .Y(ori_ori_n168_));
  NA2        o152(.A(x8), .B(x0), .Y(ori_ori_n169_));
  NO2        o153(.A(ori_ori_n146_), .B(ori_ori_n25_), .Y(ori_ori_n170_));
  NA2        o154(.A(x2), .B(x0), .Y(ori_ori_n171_));
  NA2        o155(.A(x4), .B(x1), .Y(ori_ori_n172_));
  NAi21      o156(.An(ori_ori_n114_), .B(ori_ori_n172_), .Y(ori_ori_n173_));
  NOi31      o157(.An(ori_ori_n173_), .B(ori_ori_n149_), .C(ori_ori_n171_), .Y(ori_ori_n174_));
  NO3        o158(.A(ori_ori_n174_), .B(ori_ori_n168_), .C(ori_ori_n164_), .Y(ori_ori_n175_));
  NO2        o159(.A(ori_ori_n175_), .B(ori_ori_n43_), .Y(ori_ori_n176_));
  NO2        o160(.A(ori_ori_n167_), .B(ori_ori_n73_), .Y(ori_ori_n177_));
  INV        o161(.A(ori_ori_n123_), .Y(ori_ori_n178_));
  NO2        o162(.A(ori_ori_n101_), .B(ori_ori_n17_), .Y(ori_ori_n179_));
  AOI210     o163(.A0(ori_ori_n35_), .A1(ori_ori_n87_), .B0(ori_ori_n179_), .Y(ori_ori_n180_));
  NO3        o164(.A(ori_ori_n180_), .B(ori_ori_n178_), .C(x7), .Y(ori_ori_n181_));
  NA3        o165(.A(ori_ori_n173_), .B(ori_ori_n178_), .C(ori_ori_n42_), .Y(ori_ori_n182_));
  OAI210     o166(.A0(ori_ori_n166_), .A1(ori_ori_n130_), .B0(ori_ori_n182_), .Y(ori_ori_n183_));
  NO3        o167(.A(ori_ori_n183_), .B(ori_ori_n181_), .C(ori_ori_n177_), .Y(ori_ori_n184_));
  NO2        o168(.A(ori_ori_n184_), .B(x3), .Y(ori_ori_n185_));
  NO3        o169(.A(ori_ori_n185_), .B(ori_ori_n176_), .C(ori_ori_n163_), .Y(ori03));
  NO2        o170(.A(ori_ori_n48_), .B(x3), .Y(ori_ori_n187_));
  NO2        o171(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n188_));
  NO2        o172(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n189_));
  NO2        o173(.A(ori_ori_n75_), .B(x6), .Y(ori_ori_n190_));
  NA2        o174(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n191_));
  NO2        o175(.A(ori_ori_n191_), .B(x4), .Y(ori_ori_n192_));
  NO2        o176(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n193_));
  AO220      o177(.A0(ori_ori_n193_), .A1(ori_ori_n192_), .B0(ori_ori_n190_), .B1(ori_ori_n55_), .Y(ori_ori_n194_));
  NA2        o178(.A(ori_ori_n194_), .B(ori_ori_n62_), .Y(ori_ori_n195_));
  NA2        o179(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n196_));
  NO2        o180(.A(ori_ori_n196_), .B(ori_ori_n191_), .Y(ori_ori_n197_));
  NA2        o181(.A(ori_ori_n191_), .B(ori_ori_n78_), .Y(ori_ori_n198_));
  AOI210     o182(.A0(ori_ori_n25_), .A1(x3), .B0(ori_ori_n171_), .Y(ori_ori_n199_));
  AOI220     o183(.A0(ori_ori_n199_), .A1(ori_ori_n198_), .B0(x9), .B1(ori_ori_n197_), .Y(ori_ori_n200_));
  NO3        o184(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n201_));
  NO2        o185(.A(x5), .B(x1), .Y(ori_ori_n202_));
  NO2        o186(.A(ori_ori_n196_), .B(ori_ori_n165_), .Y(ori_ori_n203_));
  NO3        o187(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n204_));
  NO2        o188(.A(ori_ori_n204_), .B(ori_ori_n203_), .Y(ori_ori_n205_));
  INV        o189(.A(ori_ori_n205_), .Y(ori_ori_n206_));
  NA2        o190(.A(ori_ori_n206_), .B(ori_ori_n48_), .Y(ori_ori_n207_));
  NA3        o191(.A(ori_ori_n207_), .B(ori_ori_n200_), .C(ori_ori_n195_), .Y(ori_ori_n208_));
  NO2        o192(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n209_));
  NA2        o193(.A(ori_ori_n209_), .B(ori_ori_n19_), .Y(ori_ori_n210_));
  NO2        o194(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n211_));
  NO2        o195(.A(ori_ori_n211_), .B(x6), .Y(ori_ori_n212_));
  NOi21      o196(.An(ori_ori_n81_), .B(ori_ori_n212_), .Y(ori_ori_n213_));
  NA2        o197(.A(ori_ori_n211_), .B(x6), .Y(ori_ori_n214_));
  AOI210     o198(.A0(ori_ori_n214_), .A1(ori_ori_n213_), .B0(ori_ori_n146_), .Y(ori_ori_n215_));
  AO210      o199(.A0(ori_ori_n215_), .A1(ori_ori_n210_), .B0(ori_ori_n170_), .Y(ori_ori_n216_));
  NA2        o200(.A(ori_ori_n43_), .B(ori_ori_n54_), .Y(ori_ori_n217_));
  OAI210     o201(.A0(ori_ori_n217_), .A1(ori_ori_n25_), .B0(ori_ori_n166_), .Y(ori_ori_n218_));
  NO2        o202(.A(ori_ori_n172_), .B(x6), .Y(ori_ori_n219_));
  AOI220     o203(.A0(ori_ori_n219_), .A1(ori_ori_n218_), .B0(ori_ori_n135_), .B1(ori_ori_n86_), .Y(ori_ori_n220_));
  NA2        o204(.A(x6), .B(ori_ori_n48_), .Y(ori_ori_n221_));
  OAI210     o205(.A0(ori_ori_n112_), .A1(ori_ori_n76_), .B0(x4), .Y(ori_ori_n222_));
  AOI210     o206(.A0(ori_ori_n222_), .A1(ori_ori_n221_), .B0(ori_ori_n75_), .Y(ori_ori_n223_));
  NO2        o207(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n224_));
  NO2        o208(.A(ori_ori_n154_), .B(ori_ori_n43_), .Y(ori_ori_n225_));
  OAI210     o209(.A0(ori_ori_n225_), .A1(ori_ori_n203_), .B0(ori_ori_n224_), .Y(ori_ori_n226_));
  NA2        o210(.A(ori_ori_n188_), .B(ori_ori_n128_), .Y(ori_ori_n227_));
  NA3        o211(.A(ori_ori_n196_), .B(ori_ori_n123_), .C(x6), .Y(ori_ori_n228_));
  OAI210     o212(.A0(ori_ori_n87_), .A1(ori_ori_n36_), .B0(ori_ori_n64_), .Y(ori_ori_n229_));
  NA4        o213(.A(ori_ori_n229_), .B(ori_ori_n228_), .C(ori_ori_n227_), .D(ori_ori_n226_), .Y(ori_ori_n230_));
  OAI210     o214(.A0(ori_ori_n230_), .A1(ori_ori_n223_), .B0(x2), .Y(ori_ori_n231_));
  NA3        o215(.A(ori_ori_n231_), .B(ori_ori_n220_), .C(ori_ori_n216_), .Y(ori_ori_n232_));
  AOI210     o216(.A0(ori_ori_n208_), .A1(x8), .B0(ori_ori_n232_), .Y(ori_ori_n233_));
  NO2        o217(.A(ori_ori_n87_), .B(x3), .Y(ori_ori_n234_));
  NA2        o218(.A(ori_ori_n234_), .B(ori_ori_n192_), .Y(ori_ori_n235_));
  NO3        o219(.A(ori_ori_n85_), .B(ori_ori_n76_), .C(ori_ori_n25_), .Y(ori_ori_n236_));
  AOI210     o220(.A0(ori_ori_n212_), .A1(ori_ori_n149_), .B0(ori_ori_n236_), .Y(ori_ori_n237_));
  AOI210     o221(.A0(ori_ori_n237_), .A1(ori_ori_n235_), .B0(x2), .Y(ori_ori_n238_));
  NO2        o222(.A(x4), .B(ori_ori_n54_), .Y(ori_ori_n239_));
  AOI220     o223(.A0(ori_ori_n192_), .A1(ori_ori_n179_), .B0(ori_ori_n239_), .B1(ori_ori_n64_), .Y(ori_ori_n240_));
  NA2        o224(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n241_));
  NA2        o225(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n242_));
  NO2        o226(.A(ori_ori_n242_), .B(ori_ori_n25_), .Y(ori_ori_n243_));
  NA2        o227(.A(ori_ori_n243_), .B(ori_ori_n114_), .Y(ori_ori_n244_));
  NA2        o228(.A(ori_ori_n196_), .B(x6), .Y(ori_ori_n245_));
  NO2        o229(.A(ori_ori_n196_), .B(x6), .Y(ori_ori_n246_));
  INV        o230(.A(ori_ori_n246_), .Y(ori_ori_n247_));
  NA3        o231(.A(ori_ori_n247_), .B(ori_ori_n245_), .C(ori_ori_n140_), .Y(ori_ori_n248_));
  NA4        o232(.A(ori_ori_n248_), .B(ori_ori_n244_), .C(ori_ori_n240_), .D(ori_ori_n146_), .Y(ori_ori_n249_));
  NA2        o233(.A(ori_ori_n188_), .B(ori_ori_n211_), .Y(ori_ori_n250_));
  NO2        o234(.A(ori_ori_n134_), .B(ori_ori_n18_), .Y(ori_ori_n251_));
  NAi21      o235(.An(x1), .B(x4), .Y(ori_ori_n252_));
  AOI210     o236(.A0(x3), .A1(x2), .B0(ori_ori_n48_), .Y(ori_ori_n253_));
  OAI210     o237(.A0(ori_ori_n134_), .A1(x3), .B0(ori_ori_n253_), .Y(ori_ori_n254_));
  NA2        o238(.A(ori_ori_n254_), .B(ori_ori_n252_), .Y(ori_ori_n255_));
  NA2        o239(.A(ori_ori_n255_), .B(ori_ori_n250_), .Y(ori_ori_n256_));
  NA2        o240(.A(ori_ori_n62_), .B(x2), .Y(ori_ori_n257_));
  NA2        o241(.A(x6), .B(x2), .Y(ori_ori_n258_));
  NA2        o242(.A(x4), .B(ori_ori_n256_), .Y(ori_ori_n259_));
  NA2        o243(.A(x9), .B(ori_ori_n43_), .Y(ori_ori_n260_));
  NO2        o244(.A(ori_ori_n260_), .B(ori_ori_n191_), .Y(ori_ori_n261_));
  OR3        o245(.A(ori_ori_n261_), .B(ori_ori_n190_), .C(ori_ori_n142_), .Y(ori_ori_n262_));
  NA2        o246(.A(x4), .B(x0), .Y(ori_ori_n263_));
  NA2        o247(.A(ori_ori_n262_), .B(ori_ori_n42_), .Y(ori_ori_n264_));
  AOI210     o248(.A0(ori_ori_n264_), .A1(ori_ori_n259_), .B0(x8), .Y(ori_ori_n265_));
  INV        o249(.A(ori_ori_n241_), .Y(ori_ori_n266_));
  OAI210     o250(.A0(ori_ori_n251_), .A1(ori_ori_n202_), .B0(ori_ori_n266_), .Y(ori_ori_n267_));
  INV        o251(.A(ori_ori_n169_), .Y(ori_ori_n268_));
  OAI210     o252(.A0(ori_ori_n268_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n269_));
  AOI210     o253(.A0(ori_ori_n269_), .A1(ori_ori_n267_), .B0(ori_ori_n217_), .Y(ori_ori_n270_));
  NO4        o254(.A(ori_ori_n270_), .B(ori_ori_n265_), .C(ori_ori_n249_), .D(ori_ori_n238_), .Y(ori_ori_n271_));
  INV        o255(.A(x1), .Y(ori_ori_n272_));
  NO3        o256(.A(ori_ori_n272_), .B(x3), .C(ori_ori_n36_), .Y(ori_ori_n273_));
  OAI210     o257(.A0(ori_ori_n273_), .A1(ori_ori_n246_), .B0(x2), .Y(ori_ori_n274_));
  OAI210     o258(.A0(ori_ori_n268_), .A1(x6), .B0(ori_ori_n44_), .Y(ori_ori_n275_));
  AOI210     o259(.A0(ori_ori_n275_), .A1(ori_ori_n274_), .B0(ori_ori_n178_), .Y(ori_ori_n276_));
  NOi21      o260(.An(ori_ori_n258_), .B(ori_ori_n17_), .Y(ori_ori_n277_));
  NA3        o261(.A(ori_ori_n277_), .B(ori_ori_n202_), .C(ori_ori_n40_), .Y(ori_ori_n278_));
  AOI210     o262(.A0(ori_ori_n36_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n279_));
  NA3        o263(.A(ori_ori_n279_), .B(ori_ori_n155_), .C(ori_ori_n32_), .Y(ori_ori_n280_));
  NA2        o264(.A(x3), .B(x2), .Y(ori_ori_n281_));
  AOI220     o265(.A0(ori_ori_n281_), .A1(ori_ori_n217_), .B0(ori_ori_n280_), .B1(ori_ori_n278_), .Y(ori_ori_n282_));
  NAi21      o266(.An(x4), .B(x0), .Y(ori_ori_n283_));
  NO3        o267(.A(ori_ori_n283_), .B(ori_ori_n44_), .C(x2), .Y(ori_ori_n284_));
  OAI210     o268(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n284_), .Y(ori_ori_n285_));
  OAI220     o269(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n286_));
  NO2        o270(.A(ori_ori_n279_), .B(ori_ori_n277_), .Y(ori_ori_n287_));
  AOI220     o271(.A0(ori_ori_n287_), .A1(ori_ori_n79_), .B0(ori_ori_n286_), .B1(ori_ori_n31_), .Y(ori_ori_n288_));
  AOI210     o272(.A0(ori_ori_n288_), .A1(ori_ori_n285_), .B0(ori_ori_n25_), .Y(ori_ori_n289_));
  NA3        o273(.A(ori_ori_n36_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n290_));
  OAI210     o274(.A0(ori_ori_n279_), .A1(ori_ori_n277_), .B0(ori_ori_n290_), .Y(ori_ori_n291_));
  INV        o275(.A(ori_ori_n203_), .Y(ori_ori_n292_));
  NA2        o276(.A(ori_ori_n36_), .B(ori_ori_n43_), .Y(ori_ori_n293_));
  OR2        o277(.A(ori_ori_n293_), .B(ori_ori_n263_), .Y(ori_ori_n294_));
  OAI220     o278(.A0(ori_ori_n294_), .A1(ori_ori_n154_), .B0(ori_ori_n221_), .B1(ori_ori_n292_), .Y(ori_ori_n295_));
  AO210      o279(.A0(ori_ori_n291_), .A1(ori_ori_n142_), .B0(ori_ori_n295_), .Y(ori_ori_n296_));
  NO4        o280(.A(ori_ori_n296_), .B(ori_ori_n289_), .C(ori_ori_n282_), .D(ori_ori_n276_), .Y(ori_ori_n297_));
  OAI210     o281(.A0(ori_ori_n271_), .A1(ori_ori_n233_), .B0(ori_ori_n297_), .Y(ori04));
  NO2        o282(.A(x2), .B(x1), .Y(ori_ori_n299_));
  OAI210     o283(.A0(ori_ori_n242_), .A1(ori_ori_n299_), .B0(ori_ori_n36_), .Y(ori_ori_n300_));
  INV        o284(.A(ori_ori_n283_), .Y(ori_ori_n301_));
  OAI210     o285(.A0(ori_ori_n54_), .A1(ori_ori_n301_), .B0(ori_ori_n234_), .Y(ori_ori_n302_));
  NO2        o286(.A(ori_ori_n281_), .B(ori_ori_n193_), .Y(ori_ori_n303_));
  NA2        o287(.A(x9), .B(x0), .Y(ori_ori_n304_));
  AOI210     o288(.A0(ori_ori_n85_), .A1(ori_ori_n73_), .B0(ori_ori_n304_), .Y(ori_ori_n305_));
  OAI210     o289(.A0(ori_ori_n305_), .A1(ori_ori_n303_), .B0(ori_ori_n87_), .Y(ori_ori_n306_));
  NA3        o290(.A(ori_ori_n306_), .B(x6), .C(ori_ori_n302_), .Y(ori_ori_n307_));
  NA2        o291(.A(ori_ori_n307_), .B(ori_ori_n300_), .Y(ori_ori_n308_));
  OAI210     o292(.A0(ori_ori_n111_), .A1(ori_ori_n101_), .B0(ori_ori_n169_), .Y(ori_ori_n309_));
  NA3        o293(.A(ori_ori_n309_), .B(x6), .C(x3), .Y(ori_ori_n310_));
  NOi21      o294(.An(ori_ori_n144_), .B(ori_ori_n124_), .Y(ori_ori_n311_));
  AOI210     o295(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n312_));
  NO2        o296(.A(ori_ori_n312_), .B(ori_ori_n293_), .Y(ori_ori_n313_));
  AOI210     o297(.A0(ori_ori_n311_), .A1(x6), .B0(ori_ori_n313_), .Y(ori_ori_n314_));
  NA2        o298(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n315_));
  OAI210     o299(.A0(ori_ori_n101_), .A1(ori_ori_n17_), .B0(ori_ori_n315_), .Y(ori_ori_n316_));
  NA2        o300(.A(ori_ori_n316_), .B(ori_ori_n76_), .Y(ori_ori_n317_));
  NA3        o301(.A(ori_ori_n317_), .B(ori_ori_n314_), .C(ori_ori_n310_), .Y(ori_ori_n318_));
  OAI210     o302(.A0(ori_ori_n106_), .A1(x3), .B0(ori_ori_n284_), .Y(ori_ori_n319_));
  NA2        o303(.A(ori_ori_n201_), .B(ori_ori_n81_), .Y(ori_ori_n320_));
  NA3        o304(.A(ori_ori_n320_), .B(ori_ori_n319_), .C(ori_ori_n146_), .Y(ori_ori_n321_));
  AOI210     o305(.A0(ori_ori_n318_), .A1(x4), .B0(ori_ori_n321_), .Y(ori_ori_n322_));
  NOi21      o306(.An(x4), .B(x0), .Y(ori_ori_n323_));
  XO2        o307(.A(x4), .B(x0), .Y(ori_ori_n324_));
  INV        o308(.A(ori_ori_n252_), .Y(ori_ori_n325_));
  AOI220     o309(.A0(ori_ori_n325_), .A1(x8), .B0(ori_ori_n323_), .B1(ori_ori_n88_), .Y(ori_ori_n326_));
  NO2        o310(.A(ori_ori_n326_), .B(x3), .Y(ori_ori_n327_));
  INV        o311(.A(ori_ori_n88_), .Y(ori_ori_n328_));
  NO2        o312(.A(ori_ori_n87_), .B(x4), .Y(ori_ori_n329_));
  AOI220     o313(.A0(ori_ori_n329_), .A1(ori_ori_n44_), .B0(ori_ori_n118_), .B1(ori_ori_n328_), .Y(ori_ori_n330_));
  NO2        o314(.A(ori_ori_n324_), .B(x2), .Y(ori_ori_n331_));
  INV        o315(.A(ori_ori_n331_), .Y(ori_ori_n332_));
  NA4        o316(.A(ori_ori_n332_), .B(ori_ori_n330_), .C(ori_ori_n210_), .D(x6), .Y(ori_ori_n333_));
  OAI220     o317(.A0(ori_ori_n283_), .A1(ori_ori_n85_), .B0(ori_ori_n171_), .B1(ori_ori_n87_), .Y(ori_ori_n334_));
  NO2        o318(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n335_));
  NA2        o319(.A(ori_ori_n334_), .B(ori_ori_n61_), .Y(ori_ori_n336_));
  NO2        o320(.A(ori_ori_n144_), .B(ori_ori_n78_), .Y(ori_ori_n337_));
  NO2        o321(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n338_));
  NOi21      o322(.An(ori_ori_n114_), .B(ori_ori_n27_), .Y(ori_ori_n339_));
  AOI210     o323(.A0(ori_ori_n338_), .A1(ori_ori_n337_), .B0(ori_ori_n339_), .Y(ori_ori_n340_));
  OAI210     o324(.A0(ori_ori_n336_), .A1(ori_ori_n62_), .B0(ori_ori_n340_), .Y(ori_ori_n341_));
  OAI220     o325(.A0(ori_ori_n341_), .A1(x6), .B0(ori_ori_n333_), .B1(ori_ori_n327_), .Y(ori_ori_n342_));
  OAI210     o326(.A0(x6), .A1(ori_ori_n48_), .B0(ori_ori_n42_), .Y(ori_ori_n343_));
  OAI210     o327(.A0(ori_ori_n343_), .A1(ori_ori_n87_), .B0(ori_ori_n294_), .Y(ori_ori_n344_));
  AOI210     o328(.A0(ori_ori_n344_), .A1(ori_ori_n18_), .B0(ori_ori_n146_), .Y(ori_ori_n345_));
  AO220      o329(.A0(ori_ori_n345_), .A1(ori_ori_n342_), .B0(ori_ori_n322_), .B1(ori_ori_n308_), .Y(ori_ori_n346_));
  NA2        o330(.A(ori_ori_n338_), .B(x6), .Y(ori_ori_n347_));
  AOI210     o331(.A0(x6), .A1(x1), .B0(ori_ori_n145_), .Y(ori_ori_n348_));
  NA2        o332(.A(ori_ori_n329_), .B(x0), .Y(ori_ori_n349_));
  NA2        o333(.A(ori_ori_n81_), .B(x6), .Y(ori_ori_n350_));
  OAI210     o334(.A0(ori_ori_n349_), .A1(ori_ori_n348_), .B0(ori_ori_n350_), .Y(ori_ori_n351_));
  AOI220     o335(.A0(ori_ori_n351_), .A1(ori_ori_n347_), .B0(ori_ori_n204_), .B1(ori_ori_n49_), .Y(ori_ori_n352_));
  NA2        o336(.A(ori_ori_n352_), .B(ori_ori_n346_), .Y(ori_ori_n353_));
  AOI210     o337(.A0(ori_ori_n189_), .A1(x8), .B0(ori_ori_n106_), .Y(ori_ori_n354_));
  NA2        o338(.A(ori_ori_n354_), .B(ori_ori_n315_), .Y(ori_ori_n355_));
  NA3        o339(.A(ori_ori_n355_), .B(ori_ori_n187_), .C(ori_ori_n146_), .Y(ori_ori_n356_));
  OAI210     o340(.A0(ori_ori_n28_), .A1(x1), .B0(ori_ori_n217_), .Y(ori_ori_n357_));
  AO220      o341(.A0(ori_ori_n357_), .A1(ori_ori_n143_), .B0(ori_ori_n105_), .B1(x4), .Y(ori_ori_n358_));
  NA3        o342(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n359_));
  NA2        o343(.A(ori_ori_n209_), .B(x0), .Y(ori_ori_n360_));
  OAI220     o344(.A0(ori_ori_n360_), .A1(x2), .B0(ori_ori_n359_), .B1(ori_ori_n328_), .Y(ori_ori_n361_));
  AOI210     o345(.A0(ori_ori_n358_), .A1(ori_ori_n112_), .B0(ori_ori_n361_), .Y(ori_ori_n362_));
  AOI210     o346(.A0(ori_ori_n362_), .A1(ori_ori_n356_), .B0(ori_ori_n25_), .Y(ori_ori_n363_));
  AOI210     o347(.A0(ori_ori_n113_), .A1(ori_ori_n111_), .B0(ori_ori_n42_), .Y(ori_ori_n364_));
  NOi31      o348(.An(ori_ori_n364_), .B(ori_ori_n335_), .C(ori_ori_n172_), .Y(ori_ori_n365_));
  NA2        o349(.A(ori_ori_n365_), .B(ori_ori_n143_), .Y(ori_ori_n366_));
  NAi31      o350(.An(ori_ori_n50_), .B(ori_ori_n272_), .C(ori_ori_n170_), .Y(ori_ori_n367_));
  NA2        o351(.A(ori_ori_n367_), .B(ori_ori_n366_), .Y(ori_ori_n368_));
  OAI210     o352(.A0(ori_ori_n368_), .A1(ori_ori_n363_), .B0(x6), .Y(ori_ori_n369_));
  NA3        o353(.A(ori_ori_n55_), .B(ori_ori_n38_), .C(ori_ori_n31_), .Y(ori_ori_n370_));
  AOI210     o354(.A0(ori_ori_n370_), .A1(x0), .B0(ori_ori_n32_), .Y(ori_ori_n371_));
  NA2        o355(.A(ori_ori_n187_), .B(ori_ori_n146_), .Y(ori_ori_n372_));
  AOI210     o356(.A0(ori_ori_n120_), .A1(ori_ori_n239_), .B0(x1), .Y(ori_ori_n373_));
  OAI210     o357(.A0(ori_ori_n372_), .A1(x8), .B0(ori_ori_n373_), .Y(ori_ori_n374_));
  NAi31      o358(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n375_));
  OAI210     o359(.A0(ori_ori_n375_), .A1(x4), .B0(ori_ori_n157_), .Y(ori_ori_n376_));
  NA3        o360(.A(ori_ori_n376_), .B(ori_ori_n141_), .C(x9), .Y(ori_ori_n377_));
  NA2        o361(.A(ori_ori_n337_), .B(ori_ori_n146_), .Y(ori_ori_n378_));
  NA4        o362(.A(ori_ori_n378_), .B(x1), .C(ori_ori_n377_), .D(ori_ori_n50_), .Y(ori_ori_n379_));
  OAI210     o363(.A0(ori_ori_n374_), .A1(ori_ori_n371_), .B0(ori_ori_n379_), .Y(ori_ori_n380_));
  AOI210     o364(.A0(ori_ori_n38_), .A1(x9), .B0(ori_ori_n127_), .Y(ori_ori_n381_));
  NO3        o365(.A(ori_ori_n381_), .B(ori_ori_n117_), .C(ori_ori_n43_), .Y(ori_ori_n382_));
  NOi31      o366(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n383_));
  AOI220     o367(.A0(ori_ori_n383_), .A1(ori_ori_n323_), .B0(ori_ori_n118_), .B1(x3), .Y(ori_ori_n384_));
  AOI210     o368(.A0(ori_ori_n252_), .A1(ori_ori_n60_), .B0(ori_ori_n116_), .Y(ori_ori_n385_));
  OAI210     o369(.A0(ori_ori_n385_), .A1(x3), .B0(ori_ori_n384_), .Y(ori_ori_n386_));
  NO3        o370(.A(ori_ori_n386_), .B(ori_ori_n382_), .C(x2), .Y(ori_ori_n387_));
  OAI210     o371(.A0(ori_ori_n283_), .A1(ori_ori_n43_), .B0(ori_ori_n324_), .Y(ori_ori_n388_));
  AOI210     o372(.A0(x9), .A1(ori_ori_n48_), .B0(ori_ori_n359_), .Y(ori_ori_n389_));
  AOI220     o373(.A0(ori_ori_n389_), .A1(ori_ori_n87_), .B0(ori_ori_n388_), .B1(ori_ori_n146_), .Y(ori_ori_n390_));
  NO2        o374(.A(ori_ori_n390_), .B(ori_ori_n54_), .Y(ori_ori_n391_));
  NO2        o375(.A(ori_ori_n391_), .B(ori_ori_n387_), .Y(ori_ori_n392_));
  AOI210     o376(.A0(ori_ori_n392_), .A1(ori_ori_n380_), .B0(ori_ori_n25_), .Y(ori_ori_n393_));
  NA4        o377(.A(ori_ori_n31_), .B(ori_ori_n87_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n394_));
  NO3        o378(.A(ori_ori_n62_), .B(x4), .C(x1), .Y(ori_ori_n395_));
  NO2        o379(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n396_));
  AOI220     o380(.A0(ori_ori_n396_), .A1(ori_ori_n253_), .B0(ori_ori_n395_), .B1(ori_ori_n364_), .Y(ori_ori_n397_));
  NO2        o381(.A(ori_ori_n397_), .B(ori_ori_n98_), .Y(ori_ori_n398_));
  NO3        o382(.A(ori_ori_n257_), .B(ori_ori_n169_), .C(ori_ori_n40_), .Y(ori_ori_n399_));
  OAI210     o383(.A0(ori_ori_n399_), .A1(ori_ori_n398_), .B0(x7), .Y(ori_ori_n400_));
  INV        o384(.A(x7), .Y(ori_ori_n401_));
  NA3        o385(.A(ori_ori_n401_), .B(ori_ori_n145_), .C(ori_ori_n128_), .Y(ori_ori_n402_));
  NA3        o386(.A(ori_ori_n402_), .B(ori_ori_n400_), .C(ori_ori_n394_), .Y(ori_ori_n403_));
  OAI210     o387(.A0(ori_ori_n403_), .A1(ori_ori_n393_), .B0(ori_ori_n36_), .Y(ori_ori_n404_));
  INV        o388(.A(ori_ori_n193_), .Y(ori_ori_n405_));
  NO4        o389(.A(ori_ori_n405_), .B(ori_ori_n75_), .C(x4), .D(ori_ori_n54_), .Y(ori_ori_n406_));
  NA2        o390(.A(ori_ori_n242_), .B(ori_ori_n21_), .Y(ori_ori_n407_));
  NO2        o391(.A(ori_ori_n154_), .B(ori_ori_n129_), .Y(ori_ori_n408_));
  NA2        o392(.A(ori_ori_n408_), .B(ori_ori_n407_), .Y(ori_ori_n409_));
  AOI210     o393(.A0(ori_ori_n409_), .A1(ori_ori_n160_), .B0(ori_ori_n28_), .Y(ori_ori_n410_));
  AOI220     o394(.A0(ori_ori_n335_), .A1(ori_ori_n87_), .B0(ori_ori_n144_), .B1(ori_ori_n189_), .Y(ori_ori_n411_));
  NA3        o395(.A(ori_ori_n411_), .B(ori_ori_n375_), .C(ori_ori_n85_), .Y(ori_ori_n412_));
  NA2        o396(.A(ori_ori_n412_), .B(ori_ori_n170_), .Y(ori_ori_n413_));
  OAI220     o397(.A0(ori_ori_n260_), .A1(ori_ori_n66_), .B0(ori_ori_n154_), .B1(ori_ori_n43_), .Y(ori_ori_n414_));
  NA2        o398(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n415_));
  OAI210     o399(.A0(ori_ori_n143_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n416_));
  NO3        o400(.A(ori_ori_n383_), .B(x3), .C(ori_ori_n54_), .Y(ori_ori_n417_));
  NA2        o401(.A(ori_ori_n417_), .B(ori_ori_n416_), .Y(ori_ori_n418_));
  OAI210     o402(.A0(ori_ori_n147_), .A1(ori_ori_n415_), .B0(ori_ori_n418_), .Y(ori_ori_n419_));
  AOI220     o403(.A0(ori_ori_n419_), .A1(x0), .B0(ori_ori_n414_), .B1(ori_ori_n129_), .Y(ori_ori_n420_));
  AOI210     o404(.A0(ori_ori_n420_), .A1(ori_ori_n413_), .B0(ori_ori_n221_), .Y(ori_ori_n421_));
  NO3        o405(.A(ori_ori_n421_), .B(ori_ori_n410_), .C(ori_ori_n406_), .Y(ori_ori_n422_));
  NA3        o406(.A(ori_ori_n422_), .B(ori_ori_n404_), .C(ori_ori_n369_), .Y(ori_ori_n423_));
  AOI210     o407(.A0(ori_ori_n353_), .A1(ori_ori_n25_), .B0(ori_ori_n423_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  INV        m012(.A(mai_mai_n24_), .Y(mai_mai_n29_));
  NO2        m013(.A(x4), .B(x3), .Y(mai_mai_n30_));
  INV        m014(.A(mai_mai_n30_), .Y(mai_mai_n31_));
  OA210      m015(.A0(mai_mai_n31_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n32_));
  NOi31      m016(.An(mai_mai_n23_), .B(mai_mai_n32_), .C(mai_mai_n29_), .Y(mai00));
  NO2        m017(.A(x1), .B(x0), .Y(mai_mai_n34_));
  INV        m018(.A(x6), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n35_), .B(mai_mai_n25_), .Y(mai_mai_n36_));
  NA2        m020(.A(x4), .B(x3), .Y(mai_mai_n37_));
  NO2        m021(.A(mai_mai_n23_), .B(mai_mai_n37_), .Y(mai_mai_n38_));
  NO2        m022(.A(x2), .B(x0), .Y(mai_mai_n39_));
  INV        m023(.A(x3), .Y(mai_mai_n40_));
  NO2        m024(.A(mai_mai_n40_), .B(mai_mai_n18_), .Y(mai_mai_n41_));
  INV        m025(.A(mai_mai_n41_), .Y(mai_mai_n42_));
  NO2        m026(.A(mai_mai_n36_), .B(x4), .Y(mai_mai_n43_));
  OAI210     m027(.A0(mai_mai_n43_), .A1(mai_mai_n42_), .B0(mai_mai_n39_), .Y(mai_mai_n44_));
  INV        m028(.A(x4), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n45_), .B(mai_mai_n17_), .Y(mai_mai_n46_));
  NA2        m030(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n47_));
  OAI210     m031(.A0(mai_mai_n47_), .A1(mai_mai_n20_), .B0(mai_mai_n44_), .Y(mai_mai_n48_));
  AOI210     m032(.A0(mai_mai_n22_), .A1(mai_mai_n19_), .B0(mai_mai_n34_), .Y(mai_mai_n49_));
  INV        m033(.A(x2), .Y(mai_mai_n50_));
  NO2        m034(.A(mai_mai_n50_), .B(mai_mai_n17_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n40_), .B(mai_mai_n18_), .Y(mai_mai_n52_));
  NA2        m036(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  OAI210     m037(.A0(mai_mai_n49_), .A1(mai_mai_n31_), .B0(mai_mai_n53_), .Y(mai_mai_n54_));
  NO3        m038(.A(mai_mai_n54_), .B(mai_mai_n48_), .C(mai_mai_n38_), .Y(mai01));
  NA2        m039(.A(x8), .B(x7), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n40_), .B(x1), .Y(mai_mai_n57_));
  INV        m041(.A(x9), .Y(mai_mai_n58_));
  INV        m042(.A(x6), .Y(mai_mai_n59_));
  NO3        m043(.A(mai_mai_n59_), .B(mai_mai_n57_), .C(mai_mai_n56_), .Y(mai_mai_n60_));
  NO2        m044(.A(x7), .B(x6), .Y(mai_mai_n61_));
  NO2        m045(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n62_));
  NO2        m046(.A(x8), .B(x2), .Y(mai_mai_n63_));
  AN2        m047(.A(mai_mai_n62_), .B(mai_mai_n61_), .Y(mai_mai_n64_));
  OAI210     m048(.A0(mai_mai_n41_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n65_));
  OAI210     m049(.A0(mai_mai_n52_), .A1(mai_mai_n20_), .B0(mai_mai_n65_), .Y(mai_mai_n66_));
  NAi31      m050(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n67_));
  NO2        m051(.A(mai_mai_n66_), .B(mai_mai_n64_), .Y(mai_mai_n68_));
  OAI210     m052(.A0(mai_mai_n68_), .A1(mai_mai_n60_), .B0(x4), .Y(mai_mai_n69_));
  NA2        m053(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n70_), .A1(mai_mai_n52_), .B0(x0), .Y(mai_mai_n71_));
  NA2        m055(.A(x5), .B(x3), .Y(mai_mai_n72_));
  NO2        m056(.A(x8), .B(x6), .Y(mai_mai_n73_));
  NO4        m057(.A(mai_mai_n73_), .B(mai_mai_n72_), .C(mai_mai_n61_), .D(mai_mai_n50_), .Y(mai_mai_n74_));
  NAi21      m058(.An(x4), .B(x3), .Y(mai_mai_n75_));
  INV        m059(.A(mai_mai_n75_), .Y(mai_mai_n76_));
  NO2        m060(.A(mai_mai_n76_), .B(mai_mai_n22_), .Y(mai_mai_n77_));
  NO2        m061(.A(x4), .B(x2), .Y(mai_mai_n78_));
  NO2        m062(.A(mai_mai_n78_), .B(x3), .Y(mai_mai_n79_));
  NO3        m063(.A(mai_mai_n79_), .B(mai_mai_n77_), .C(mai_mai_n18_), .Y(mai_mai_n80_));
  NO3        m064(.A(mai_mai_n80_), .B(mai_mai_n74_), .C(mai_mai_n71_), .Y(mai_mai_n81_));
  NO4        m065(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n40_), .D(x1), .Y(mai_mai_n82_));
  NA2        m066(.A(mai_mai_n58_), .B(mai_mai_n45_), .Y(mai_mai_n83_));
  INV        m067(.A(mai_mai_n83_), .Y(mai_mai_n84_));
  OAI210     m068(.A0(mai_mai_n82_), .A1(mai_mai_n62_), .B0(mai_mai_n84_), .Y(mai_mai_n85_));
  NA2        m069(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n86_));
  NO2        m070(.A(mai_mai_n86_), .B(mai_mai_n25_), .Y(mai_mai_n87_));
  INV        m071(.A(x8), .Y(mai_mai_n88_));
  NA2        m072(.A(x2), .B(x1), .Y(mai_mai_n89_));
  NO2        m073(.A(mai_mai_n89_), .B(mai_mai_n88_), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n90_), .B(mai_mai_n87_), .Y(mai_mai_n91_));
  NO2        m075(.A(mai_mai_n91_), .B(mai_mai_n26_), .Y(mai_mai_n92_));
  AOI210     m076(.A0(mai_mai_n52_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n93_));
  OAI210     m077(.A0(mai_mai_n42_), .A1(mai_mai_n36_), .B0(mai_mai_n45_), .Y(mai_mai_n94_));
  NO3        m078(.A(mai_mai_n94_), .B(mai_mai_n93_), .C(mai_mai_n92_), .Y(mai_mai_n95_));
  NA2        m079(.A(x4), .B(mai_mai_n40_), .Y(mai_mai_n96_));
  NO2        m080(.A(mai_mai_n45_), .B(mai_mai_n50_), .Y(mai_mai_n97_));
  NO2        m081(.A(mai_mai_n96_), .B(x1), .Y(mai_mai_n98_));
  NO2        m082(.A(x3), .B(x2), .Y(mai_mai_n99_));
  NA2        m083(.A(mai_mai_n99_), .B(mai_mai_n25_), .Y(mai_mai_n100_));
  AOI210     m084(.A0(x8), .A1(x6), .B0(mai_mai_n100_), .Y(mai_mai_n101_));
  NA2        m085(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n102_));
  OAI210     m086(.A0(mai_mai_n102_), .A1(mai_mai_n37_), .B0(mai_mai_n17_), .Y(mai_mai_n103_));
  NO4        m087(.A(mai_mai_n103_), .B(mai_mai_n101_), .C(mai_mai_n98_), .D(mai_mai_n95_), .Y(mai_mai_n104_));
  AO220      m088(.A0(mai_mai_n104_), .A1(mai_mai_n85_), .B0(mai_mai_n81_), .B1(mai_mai_n69_), .Y(mai02));
  NO2        m089(.A(x3), .B(mai_mai_n50_), .Y(mai_mai_n106_));
  NO2        m090(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n107_));
  NA2        m091(.A(mai_mai_n50_), .B(mai_mai_n17_), .Y(mai_mai_n108_));
  NA2        m092(.A(mai_mai_n40_), .B(x0), .Y(mai_mai_n109_));
  OAI210     m093(.A0(mai_mai_n83_), .A1(mai_mai_n108_), .B0(mai_mai_n109_), .Y(mai_mai_n110_));
  AOI220     m094(.A0(mai_mai_n110_), .A1(mai_mai_n107_), .B0(mai_mai_n106_), .B1(x4), .Y(mai_mai_n111_));
  NO3        m095(.A(mai_mai_n111_), .B(x7), .C(x5), .Y(mai_mai_n112_));
  NA2        m096(.A(x9), .B(x2), .Y(mai_mai_n113_));
  OR2        m097(.A(x8), .B(x0), .Y(mai_mai_n114_));
  INV        m098(.A(mai_mai_n114_), .Y(mai_mai_n115_));
  NAi21      m099(.An(x2), .B(x8), .Y(mai_mai_n116_));
  INV        m100(.A(mai_mai_n116_), .Y(mai_mai_n117_));
  OAI220     m101(.A0(mai_mai_n117_), .A1(mai_mai_n115_), .B0(mai_mai_n113_), .B1(x7), .Y(mai_mai_n118_));
  NO2        m102(.A(x4), .B(x1), .Y(mai_mai_n119_));
  NA3        m103(.A(mai_mai_n119_), .B(mai_mai_n118_), .C(mai_mai_n56_), .Y(mai_mai_n120_));
  NOi21      m104(.An(x0), .B(x1), .Y(mai_mai_n121_));
  NO3        m105(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n122_));
  NOi21      m106(.An(x0), .B(x4), .Y(mai_mai_n123_));
  NAi21      m107(.An(x8), .B(x7), .Y(mai_mai_n124_));
  NO2        m108(.A(mai_mai_n120_), .B(mai_mai_n72_), .Y(mai_mai_n125_));
  NO2        m109(.A(x5), .B(mai_mai_n45_), .Y(mai_mai_n126_));
  NA2        m110(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n127_));
  AOI210     m111(.A0(mai_mai_n127_), .A1(mai_mai_n102_), .B0(mai_mai_n109_), .Y(mai_mai_n128_));
  OAI210     m112(.A0(mai_mai_n128_), .A1(mai_mai_n34_), .B0(mai_mai_n126_), .Y(mai_mai_n129_));
  NAi21      m113(.An(x0), .B(x4), .Y(mai_mai_n130_));
  NO2        m114(.A(mai_mai_n130_), .B(x1), .Y(mai_mai_n131_));
  NO2        m115(.A(x7), .B(x0), .Y(mai_mai_n132_));
  NO2        m116(.A(mai_mai_n78_), .B(mai_mai_n97_), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n133_), .B(x3), .Y(mai_mai_n134_));
  OAI210     m118(.A0(mai_mai_n132_), .A1(mai_mai_n131_), .B0(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m119(.A(mai_mai_n21_), .B(mai_mai_n40_), .Y(mai_mai_n136_));
  NA2        m120(.A(x5), .B(x0), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n138_));
  NA3        m122(.A(mai_mai_n138_), .B(mai_mai_n137_), .C(mai_mai_n136_), .Y(mai_mai_n139_));
  NA4        m123(.A(mai_mai_n139_), .B(mai_mai_n135_), .C(mai_mai_n129_), .D(mai_mai_n35_), .Y(mai_mai_n140_));
  NO3        m124(.A(mai_mai_n140_), .B(mai_mai_n125_), .C(mai_mai_n112_), .Y(mai_mai_n141_));
  NO3        m125(.A(mai_mai_n72_), .B(mai_mai_n70_), .C(mai_mai_n24_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n143_));
  AOI220     m127(.A0(mai_mai_n121_), .A1(mai_mai_n143_), .B0(mai_mai_n62_), .B1(mai_mai_n17_), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n144_), .B(mai_mai_n56_), .Y(mai_mai_n145_));
  NA2        m129(.A(x7), .B(x3), .Y(mai_mai_n146_));
  NO2        m130(.A(mai_mai_n96_), .B(x5), .Y(mai_mai_n147_));
  NO2        m131(.A(x9), .B(x7), .Y(mai_mai_n148_));
  NOi21      m132(.An(x8), .B(x0), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n40_), .B(x2), .Y(mai_mai_n150_));
  INV        m134(.A(x7), .Y(mai_mai_n151_));
  NA2        m135(.A(mai_mai_n151_), .B(mai_mai_n18_), .Y(mai_mai_n152_));
  NA2        m136(.A(mai_mai_n152_), .B(mai_mai_n150_), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n154_));
  NO2        m138(.A(mai_mai_n154_), .B(mai_mai_n123_), .Y(mai_mai_n155_));
  NO2        m139(.A(mai_mai_n155_), .B(mai_mai_n153_), .Y(mai_mai_n156_));
  AOI210     m140(.A0(mai_mai_n149_), .A1(mai_mai_n147_), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  OAI210     m141(.A0(mai_mai_n146_), .A1(mai_mai_n47_), .B0(mai_mai_n157_), .Y(mai_mai_n158_));
  NA2        m142(.A(x5), .B(x1), .Y(mai_mai_n159_));
  INV        m143(.A(mai_mai_n159_), .Y(mai_mai_n160_));
  AOI210     m144(.A0(mai_mai_n160_), .A1(mai_mai_n123_), .B0(mai_mai_n35_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n58_), .B(mai_mai_n88_), .Y(mai_mai_n162_));
  NAi21      m146(.An(x2), .B(x7), .Y(mai_mai_n163_));
  INV        m147(.A(mai_mai_n161_), .Y(mai_mai_n164_));
  NO4        m148(.A(mai_mai_n164_), .B(mai_mai_n158_), .C(mai_mai_n145_), .D(mai_mai_n142_), .Y(mai_mai_n165_));
  NO2        m149(.A(mai_mai_n165_), .B(mai_mai_n141_), .Y(mai_mai_n166_));
  NO2        m150(.A(mai_mai_n137_), .B(mai_mai_n133_), .Y(mai_mai_n167_));
  NA2        m151(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n168_));
  NA2        m152(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n169_));
  NA3        m153(.A(mai_mai_n169_), .B(mai_mai_n168_), .C(mai_mai_n24_), .Y(mai_mai_n170_));
  AN2        m154(.A(mai_mai_n170_), .B(mai_mai_n138_), .Y(mai_mai_n171_));
  NA2        m155(.A(x8), .B(x0), .Y(mai_mai_n172_));
  NO2        m156(.A(mai_mai_n151_), .B(mai_mai_n25_), .Y(mai_mai_n173_));
  NO2        m157(.A(mai_mai_n121_), .B(x4), .Y(mai_mai_n174_));
  NA2        m158(.A(mai_mai_n174_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  AOI210     m159(.A0(mai_mai_n172_), .A1(mai_mai_n127_), .B0(mai_mai_n175_), .Y(mai_mai_n176_));
  NA2        m160(.A(x2), .B(x0), .Y(mai_mai_n177_));
  NA2        m161(.A(x4), .B(x1), .Y(mai_mai_n178_));
  NAi21      m162(.An(mai_mai_n119_), .B(mai_mai_n178_), .Y(mai_mai_n179_));
  NOi31      m163(.An(mai_mai_n179_), .B(mai_mai_n154_), .C(mai_mai_n177_), .Y(mai_mai_n180_));
  NO4        m164(.A(mai_mai_n180_), .B(mai_mai_n176_), .C(mai_mai_n171_), .D(mai_mai_n167_), .Y(mai_mai_n181_));
  NO2        m165(.A(mai_mai_n181_), .B(mai_mai_n40_), .Y(mai_mai_n182_));
  NO2        m166(.A(mai_mai_n170_), .B(mai_mai_n70_), .Y(mai_mai_n183_));
  INV        m167(.A(mai_mai_n126_), .Y(mai_mai_n184_));
  NO2        m168(.A(mai_mai_n102_), .B(mai_mai_n17_), .Y(mai_mai_n185_));
  AOI210     m169(.A0(mai_mai_n34_), .A1(mai_mai_n88_), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  NO3        m170(.A(mai_mai_n186_), .B(mai_mai_n184_), .C(x7), .Y(mai_mai_n187_));
  NA3        m171(.A(mai_mai_n179_), .B(mai_mai_n184_), .C(mai_mai_n39_), .Y(mai_mai_n188_));
  OAI210     m172(.A0(mai_mai_n169_), .A1(mai_mai_n133_), .B0(mai_mai_n188_), .Y(mai_mai_n189_));
  NO3        m173(.A(mai_mai_n189_), .B(mai_mai_n187_), .C(mai_mai_n183_), .Y(mai_mai_n190_));
  NO2        m174(.A(mai_mai_n190_), .B(x3), .Y(mai_mai_n191_));
  NO3        m175(.A(mai_mai_n191_), .B(mai_mai_n182_), .C(mai_mai_n166_), .Y(mai03));
  NO2        m176(.A(mai_mai_n45_), .B(x3), .Y(mai_mai_n193_));
  NO2        m177(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n194_));
  INV        m178(.A(mai_mai_n194_), .Y(mai_mai_n195_));
  NO2        m179(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n196_));
  OAI210     m180(.A0(mai_mai_n196_), .A1(mai_mai_n25_), .B0(x6), .Y(mai_mai_n197_));
  OAI220     m181(.A0(mai_mai_n197_), .A1(mai_mai_n17_), .B0(mai_mai_n195_), .B1(mai_mai_n102_), .Y(mai_mai_n198_));
  NA2        m182(.A(mai_mai_n198_), .B(mai_mai_n193_), .Y(mai_mai_n199_));
  NO2        m183(.A(mai_mai_n72_), .B(x6), .Y(mai_mai_n200_));
  NA2        m184(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n201_), .B(x4), .Y(mai_mai_n202_));
  NO2        m186(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n203_));
  AO220      m187(.A0(mai_mai_n203_), .A1(mai_mai_n202_), .B0(mai_mai_n200_), .B1(mai_mai_n51_), .Y(mai_mai_n204_));
  INV        m188(.A(mai_mai_n204_), .Y(mai_mai_n205_));
  NA2        m189(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n206_));
  NA2        m190(.A(x9), .B(mai_mai_n50_), .Y(mai_mai_n207_));
  NO3        m191(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n208_));
  NO2        m192(.A(x5), .B(x1), .Y(mai_mai_n209_));
  AOI220     m193(.A0(mai_mai_n209_), .A1(mai_mai_n17_), .B0(mai_mai_n99_), .B1(x5), .Y(mai_mai_n210_));
  NO2        m194(.A(mai_mai_n206_), .B(mai_mai_n168_), .Y(mai_mai_n211_));
  INV        m195(.A(mai_mai_n211_), .Y(mai_mai_n212_));
  OAI210     m196(.A0(mai_mai_n210_), .A1(mai_mai_n59_), .B0(mai_mai_n212_), .Y(mai_mai_n213_));
  AOI220     m197(.A0(mai_mai_n213_), .A1(mai_mai_n45_), .B0(mai_mai_n208_), .B1(mai_mai_n126_), .Y(mai_mai_n214_));
  NA3        m198(.A(mai_mai_n214_), .B(mai_mai_n205_), .C(mai_mai_n199_), .Y(mai_mai_n215_));
  NO2        m199(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n216_));
  NA2        m200(.A(mai_mai_n216_), .B(mai_mai_n19_), .Y(mai_mai_n217_));
  NO2        m201(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n218_));
  NO2        m202(.A(mai_mai_n218_), .B(x6), .Y(mai_mai_n219_));
  NOi21      m203(.An(mai_mai_n78_), .B(mai_mai_n219_), .Y(mai_mai_n220_));
  NA2        m204(.A(mai_mai_n58_), .B(mai_mai_n88_), .Y(mai_mai_n221_));
  NA3        m205(.A(mai_mai_n221_), .B(mai_mai_n218_), .C(x6), .Y(mai_mai_n222_));
  AOI210     m206(.A0(mai_mai_n222_), .A1(mai_mai_n220_), .B0(mai_mai_n151_), .Y(mai_mai_n223_));
  AO210      m207(.A0(mai_mai_n223_), .A1(mai_mai_n217_), .B0(mai_mai_n173_), .Y(mai_mai_n224_));
  NA2        m208(.A(mai_mai_n40_), .B(mai_mai_n50_), .Y(mai_mai_n225_));
  NA2        m209(.A(mai_mai_n138_), .B(mai_mai_n87_), .Y(mai_mai_n226_));
  NA2        m210(.A(x6), .B(mai_mai_n45_), .Y(mai_mai_n227_));
  OAI210     m211(.A0(mai_mai_n115_), .A1(mai_mai_n73_), .B0(x4), .Y(mai_mai_n228_));
  AOI210     m212(.A0(mai_mai_n228_), .A1(mai_mai_n227_), .B0(mai_mai_n72_), .Y(mai_mai_n229_));
  NA2        m213(.A(mai_mai_n194_), .B(mai_mai_n131_), .Y(mai_mai_n230_));
  NA3        m214(.A(mai_mai_n206_), .B(mai_mai_n126_), .C(x6), .Y(mai_mai_n231_));
  OAI210     m215(.A0(mai_mai_n88_), .A1(mai_mai_n35_), .B0(mai_mai_n62_), .Y(mai_mai_n232_));
  NA3        m216(.A(mai_mai_n232_), .B(mai_mai_n231_), .C(mai_mai_n230_), .Y(mai_mai_n233_));
  OAI210     m217(.A0(mai_mai_n233_), .A1(mai_mai_n229_), .B0(x2), .Y(mai_mai_n234_));
  NA3        m218(.A(mai_mai_n234_), .B(mai_mai_n226_), .C(mai_mai_n224_), .Y(mai_mai_n235_));
  AOI210     m219(.A0(mai_mai_n215_), .A1(x8), .B0(mai_mai_n235_), .Y(mai_mai_n236_));
  NO2        m220(.A(mai_mai_n88_), .B(x3), .Y(mai_mai_n237_));
  NA2        m221(.A(mai_mai_n237_), .B(mai_mai_n202_), .Y(mai_mai_n238_));
  NO2        m222(.A(mai_mai_n86_), .B(mai_mai_n25_), .Y(mai_mai_n239_));
  AOI210     m223(.A0(mai_mai_n219_), .A1(mai_mai_n154_), .B0(mai_mai_n239_), .Y(mai_mai_n240_));
  AOI210     m224(.A0(mai_mai_n240_), .A1(mai_mai_n238_), .B0(x2), .Y(mai_mai_n241_));
  NO2        m225(.A(x4), .B(mai_mai_n50_), .Y(mai_mai_n242_));
  AOI220     m226(.A0(mai_mai_n202_), .A1(mai_mai_n185_), .B0(mai_mai_n242_), .B1(mai_mai_n62_), .Y(mai_mai_n243_));
  NA2        m227(.A(mai_mai_n58_), .B(x6), .Y(mai_mai_n244_));
  NA3        m228(.A(mai_mai_n25_), .B(x3), .C(x2), .Y(mai_mai_n245_));
  AOI210     m229(.A0(mai_mai_n245_), .A1(mai_mai_n137_), .B0(mai_mai_n244_), .Y(mai_mai_n246_));
  NA2        m230(.A(mai_mai_n40_), .B(mai_mai_n17_), .Y(mai_mai_n247_));
  NO2        m231(.A(mai_mai_n247_), .B(mai_mai_n25_), .Y(mai_mai_n248_));
  OAI210     m232(.A0(mai_mai_n248_), .A1(mai_mai_n246_), .B0(mai_mai_n119_), .Y(mai_mai_n249_));
  NA2        m233(.A(mai_mai_n206_), .B(x6), .Y(mai_mai_n250_));
  NO2        m234(.A(mai_mai_n206_), .B(x6), .Y(mai_mai_n251_));
  NAi21      m235(.An(mai_mai_n162_), .B(mai_mai_n251_), .Y(mai_mai_n252_));
  NA3        m236(.A(mai_mai_n252_), .B(mai_mai_n250_), .C(mai_mai_n143_), .Y(mai_mai_n253_));
  NA4        m237(.A(mai_mai_n253_), .B(mai_mai_n249_), .C(mai_mai_n243_), .D(mai_mai_n151_), .Y(mai_mai_n254_));
  NA2        m238(.A(mai_mai_n194_), .B(mai_mai_n218_), .Y(mai_mai_n255_));
  NO2        m239(.A(x9), .B(x6), .Y(mai_mai_n256_));
  NO2        m240(.A(mai_mai_n137_), .B(mai_mai_n18_), .Y(mai_mai_n257_));
  NAi21      m241(.An(mai_mai_n257_), .B(mai_mai_n245_), .Y(mai_mai_n258_));
  NAi21      m242(.An(x1), .B(x4), .Y(mai_mai_n259_));
  AOI210     m243(.A0(x3), .A1(x2), .B0(mai_mai_n45_), .Y(mai_mai_n260_));
  OAI210     m244(.A0(mai_mai_n137_), .A1(x3), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  AOI220     m245(.A0(mai_mai_n261_), .A1(mai_mai_n259_), .B0(mai_mai_n258_), .B1(mai_mai_n256_), .Y(mai_mai_n262_));
  NA2        m246(.A(mai_mai_n262_), .B(mai_mai_n255_), .Y(mai_mai_n263_));
  NA2        m247(.A(mai_mai_n58_), .B(x2), .Y(mai_mai_n264_));
  NO2        m248(.A(mai_mai_n264_), .B(mai_mai_n255_), .Y(mai_mai_n265_));
  NO3        m249(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n266_));
  NA2        m250(.A(mai_mai_n102_), .B(mai_mai_n25_), .Y(mai_mai_n267_));
  NA2        m251(.A(x6), .B(x2), .Y(mai_mai_n268_));
  NO2        m252(.A(mai_mai_n268_), .B(mai_mai_n168_), .Y(mai_mai_n269_));
  AOI210     m253(.A0(mai_mai_n267_), .A1(mai_mai_n266_), .B0(mai_mai_n269_), .Y(mai_mai_n270_));
  OAI220     m254(.A0(mai_mai_n270_), .A1(mai_mai_n40_), .B0(mai_mai_n174_), .B1(mai_mai_n43_), .Y(mai_mai_n271_));
  OAI210     m255(.A0(mai_mai_n271_), .A1(mai_mai_n265_), .B0(mai_mai_n263_), .Y(mai_mai_n272_));
  NA2        m256(.A(x4), .B(x0), .Y(mai_mai_n273_));
  NA2        m257(.A(mai_mai_n200_), .B(mai_mai_n39_), .Y(mai_mai_n274_));
  AOI210     m258(.A0(mai_mai_n274_), .A1(mai_mai_n272_), .B0(x8), .Y(mai_mai_n275_));
  NA2        m259(.A(mai_mai_n209_), .B(x6), .Y(mai_mai_n276_));
  INV        m260(.A(mai_mai_n172_), .Y(mai_mai_n277_));
  OAI210     m261(.A0(mai_mai_n277_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n278_));
  AOI210     m262(.A0(mai_mai_n278_), .A1(mai_mai_n276_), .B0(mai_mai_n225_), .Y(mai_mai_n279_));
  NO4        m263(.A(mai_mai_n279_), .B(mai_mai_n275_), .C(mai_mai_n254_), .D(mai_mai_n241_), .Y(mai_mai_n280_));
  NO2        m264(.A(mai_mai_n162_), .B(x1), .Y(mai_mai_n281_));
  NO3        m265(.A(mai_mai_n281_), .B(x3), .C(mai_mai_n35_), .Y(mai_mai_n282_));
  OAI210     m266(.A0(mai_mai_n282_), .A1(mai_mai_n251_), .B0(x2), .Y(mai_mai_n283_));
  OAI210     m267(.A0(mai_mai_n277_), .A1(x6), .B0(mai_mai_n41_), .Y(mai_mai_n284_));
  AOI210     m268(.A0(mai_mai_n284_), .A1(mai_mai_n283_), .B0(mai_mai_n184_), .Y(mai_mai_n285_));
  NOi21      m269(.An(mai_mai_n268_), .B(mai_mai_n17_), .Y(mai_mai_n286_));
  NA3        m270(.A(mai_mai_n286_), .B(mai_mai_n209_), .C(mai_mai_n37_), .Y(mai_mai_n287_));
  AOI210     m271(.A0(mai_mai_n35_), .A1(mai_mai_n50_), .B0(x0), .Y(mai_mai_n288_));
  NA3        m272(.A(mai_mai_n288_), .B(mai_mai_n160_), .C(mai_mai_n31_), .Y(mai_mai_n289_));
  NA2        m273(.A(x3), .B(x2), .Y(mai_mai_n290_));
  AOI220     m274(.A0(mai_mai_n290_), .A1(mai_mai_n225_), .B0(mai_mai_n289_), .B1(mai_mai_n287_), .Y(mai_mai_n291_));
  NAi21      m275(.An(x4), .B(x0), .Y(mai_mai_n292_));
  NO3        m276(.A(mai_mai_n292_), .B(mai_mai_n41_), .C(x2), .Y(mai_mai_n293_));
  OAI210     m277(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n293_), .Y(mai_mai_n294_));
  OAI220     m278(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n295_));
  NO2        m279(.A(x9), .B(x8), .Y(mai_mai_n296_));
  NA3        m280(.A(mai_mai_n296_), .B(mai_mai_n35_), .C(mai_mai_n50_), .Y(mai_mai_n297_));
  OAI210     m281(.A0(mai_mai_n288_), .A1(mai_mai_n286_), .B0(mai_mai_n297_), .Y(mai_mai_n298_));
  AOI220     m282(.A0(mai_mai_n298_), .A1(mai_mai_n76_), .B0(mai_mai_n295_), .B1(mai_mai_n30_), .Y(mai_mai_n299_));
  AOI210     m283(.A0(mai_mai_n299_), .A1(mai_mai_n294_), .B0(mai_mai_n25_), .Y(mai_mai_n300_));
  NA3        m284(.A(mai_mai_n35_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n301_));
  OAI210     m285(.A0(mai_mai_n288_), .A1(mai_mai_n286_), .B0(mai_mai_n301_), .Y(mai_mai_n302_));
  INV        m286(.A(mai_mai_n211_), .Y(mai_mai_n303_));
  NA2        m287(.A(mai_mai_n35_), .B(mai_mai_n40_), .Y(mai_mai_n304_));
  OR2        m288(.A(mai_mai_n304_), .B(mai_mai_n273_), .Y(mai_mai_n305_));
  OAI220     m289(.A0(mai_mai_n305_), .A1(mai_mai_n159_), .B0(mai_mai_n227_), .B1(mai_mai_n303_), .Y(mai_mai_n306_));
  AO210      m290(.A0(mai_mai_n302_), .A1(mai_mai_n147_), .B0(mai_mai_n306_), .Y(mai_mai_n307_));
  NO4        m291(.A(mai_mai_n307_), .B(mai_mai_n300_), .C(mai_mai_n291_), .D(mai_mai_n285_), .Y(mai_mai_n308_));
  OAI210     m292(.A0(mai_mai_n280_), .A1(mai_mai_n236_), .B0(mai_mai_n308_), .Y(mai04));
  OAI210     m293(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n310_));
  NA3        m294(.A(mai_mai_n310_), .B(mai_mai_n266_), .C(mai_mai_n79_), .Y(mai_mai_n311_));
  NO2        m295(.A(x2), .B(x1), .Y(mai_mai_n312_));
  OAI210     m296(.A0(mai_mai_n247_), .A1(mai_mai_n312_), .B0(mai_mai_n35_), .Y(mai_mai_n313_));
  NO2        m297(.A(mai_mai_n312_), .B(mai_mai_n292_), .Y(mai_mai_n314_));
  AOI210     m298(.A0(mai_mai_n58_), .A1(x4), .B0(mai_mai_n108_), .Y(mai_mai_n315_));
  OAI210     m299(.A0(mai_mai_n315_), .A1(mai_mai_n314_), .B0(mai_mai_n237_), .Y(mai_mai_n316_));
  NO2        m300(.A(mai_mai_n264_), .B(mai_mai_n86_), .Y(mai_mai_n317_));
  NO2        m301(.A(mai_mai_n317_), .B(mai_mai_n35_), .Y(mai_mai_n318_));
  NO2        m302(.A(mai_mai_n290_), .B(mai_mai_n203_), .Y(mai_mai_n319_));
  NA2        m303(.A(mai_mai_n319_), .B(mai_mai_n88_), .Y(mai_mai_n320_));
  NA3        m304(.A(mai_mai_n320_), .B(mai_mai_n318_), .C(mai_mai_n316_), .Y(mai_mai_n321_));
  NA2        m305(.A(mai_mai_n321_), .B(mai_mai_n313_), .Y(mai_mai_n322_));
  NO2        m306(.A(mai_mai_n207_), .B(mai_mai_n109_), .Y(mai_mai_n323_));
  NO3        m307(.A(mai_mai_n244_), .B(mai_mai_n116_), .C(mai_mai_n18_), .Y(mai_mai_n324_));
  NO2        m308(.A(mai_mai_n324_), .B(mai_mai_n323_), .Y(mai_mai_n325_));
  OAI210     m309(.A0(mai_mai_n114_), .A1(mai_mai_n102_), .B0(mai_mai_n172_), .Y(mai_mai_n326_));
  NA3        m310(.A(mai_mai_n326_), .B(x6), .C(x3), .Y(mai_mai_n327_));
  AOI210     m311(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n328_));
  OAI220     m312(.A0(mai_mai_n328_), .A1(mai_mai_n304_), .B0(mai_mai_n264_), .B1(mai_mai_n301_), .Y(mai_mai_n329_));
  INV        m313(.A(mai_mai_n329_), .Y(mai_mai_n330_));
  NA2        m314(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n331_));
  OAI210     m315(.A0(mai_mai_n102_), .A1(mai_mai_n17_), .B0(mai_mai_n331_), .Y(mai_mai_n332_));
  AOI220     m316(.A0(mai_mai_n332_), .A1(mai_mai_n73_), .B0(mai_mai_n317_), .B1(mai_mai_n88_), .Y(mai_mai_n333_));
  NA4        m317(.A(mai_mai_n333_), .B(mai_mai_n330_), .C(mai_mai_n327_), .D(mai_mai_n325_), .Y(mai_mai_n334_));
  OAI210     m318(.A0(mai_mai_n107_), .A1(x3), .B0(mai_mai_n293_), .Y(mai_mai_n335_));
  NA3        m319(.A(mai_mai_n221_), .B(mai_mai_n208_), .C(mai_mai_n78_), .Y(mai_mai_n336_));
  NA3        m320(.A(mai_mai_n336_), .B(mai_mai_n335_), .C(mai_mai_n151_), .Y(mai_mai_n337_));
  AOI210     m321(.A0(mai_mai_n334_), .A1(x4), .B0(mai_mai_n337_), .Y(mai_mai_n338_));
  NA3        m322(.A(mai_mai_n314_), .B(mai_mai_n207_), .C(mai_mai_n88_), .Y(mai_mai_n339_));
  NOi21      m323(.An(x4), .B(x0), .Y(mai_mai_n340_));
  XO2        m324(.A(x4), .B(x0), .Y(mai_mai_n341_));
  OAI210     m325(.A0(mai_mai_n341_), .A1(mai_mai_n113_), .B0(mai_mai_n259_), .Y(mai_mai_n342_));
  AOI220     m326(.A0(mai_mai_n342_), .A1(x8), .B0(mai_mai_n340_), .B1(mai_mai_n89_), .Y(mai_mai_n343_));
  AOI210     m327(.A0(mai_mai_n343_), .A1(mai_mai_n339_), .B0(x3), .Y(mai_mai_n344_));
  INV        m328(.A(mai_mai_n89_), .Y(mai_mai_n345_));
  NO2        m329(.A(mai_mai_n88_), .B(x4), .Y(mai_mai_n346_));
  AOI220     m330(.A0(mai_mai_n346_), .A1(mai_mai_n41_), .B0(mai_mai_n123_), .B1(mai_mai_n345_), .Y(mai_mai_n347_));
  NO3        m331(.A(mai_mai_n341_), .B(mai_mai_n162_), .C(x2), .Y(mai_mai_n348_));
  NO3        m332(.A(mai_mai_n221_), .B(mai_mai_n28_), .C(mai_mai_n24_), .Y(mai_mai_n349_));
  NO2        m333(.A(mai_mai_n349_), .B(mai_mai_n348_), .Y(mai_mai_n350_));
  NA4        m334(.A(mai_mai_n350_), .B(mai_mai_n347_), .C(mai_mai_n217_), .D(x6), .Y(mai_mai_n351_));
  OAI220     m335(.A0(mai_mai_n292_), .A1(mai_mai_n86_), .B0(mai_mai_n177_), .B1(mai_mai_n88_), .Y(mai_mai_n352_));
  BUFFER     m336(.A(mai_mai_n346_), .Y(mai_mai_n353_));
  NO2        m337(.A(mai_mai_n149_), .B(mai_mai_n102_), .Y(mai_mai_n354_));
  AOI220     m338(.A0(mai_mai_n354_), .A1(mai_mai_n353_), .B0(mai_mai_n352_), .B1(mai_mai_n57_), .Y(mai_mai_n355_));
  NO2        m339(.A(mai_mai_n149_), .B(mai_mai_n75_), .Y(mai_mai_n356_));
  NO2        m340(.A(mai_mai_n34_), .B(x2), .Y(mai_mai_n357_));
  NOi21      m341(.An(mai_mai_n119_), .B(mai_mai_n27_), .Y(mai_mai_n358_));
  AOI210     m342(.A0(mai_mai_n357_), .A1(mai_mai_n356_), .B0(mai_mai_n358_), .Y(mai_mai_n359_));
  OAI210     m343(.A0(mai_mai_n355_), .A1(mai_mai_n58_), .B0(mai_mai_n359_), .Y(mai_mai_n360_));
  OAI220     m344(.A0(mai_mai_n360_), .A1(x6), .B0(mai_mai_n351_), .B1(mai_mai_n344_), .Y(mai_mai_n361_));
  INV        m345(.A(mai_mai_n305_), .Y(mai_mai_n362_));
  AOI210     m346(.A0(mai_mai_n362_), .A1(mai_mai_n18_), .B0(mai_mai_n151_), .Y(mai_mai_n363_));
  AO220      m347(.A0(mai_mai_n363_), .A1(mai_mai_n361_), .B0(mai_mai_n338_), .B1(mai_mai_n322_), .Y(mai_mai_n364_));
  NA2        m348(.A(mai_mai_n357_), .B(x6), .Y(mai_mai_n365_));
  AOI210     m349(.A0(x6), .A1(x1), .B0(mai_mai_n150_), .Y(mai_mai_n366_));
  NA2        m350(.A(mai_mai_n346_), .B(x0), .Y(mai_mai_n367_));
  NA2        m351(.A(mai_mai_n78_), .B(x6), .Y(mai_mai_n368_));
  OAI210     m352(.A0(mai_mai_n367_), .A1(mai_mai_n366_), .B0(mai_mai_n368_), .Y(mai_mai_n369_));
  NA2        m353(.A(mai_mai_n369_), .B(mai_mai_n365_), .Y(mai_mai_n370_));
  NA3        m354(.A(mai_mai_n370_), .B(mai_mai_n364_), .C(mai_mai_n311_), .Y(mai_mai_n371_));
  AOI210     m355(.A0(mai_mai_n196_), .A1(x8), .B0(mai_mai_n107_), .Y(mai_mai_n372_));
  NA2        m356(.A(mai_mai_n372_), .B(mai_mai_n331_), .Y(mai_mai_n373_));
  NA3        m357(.A(mai_mai_n373_), .B(mai_mai_n193_), .C(mai_mai_n151_), .Y(mai_mai_n374_));
  OAI210     m358(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n225_), .Y(mai_mai_n375_));
  AO220      m359(.A0(mai_mai_n375_), .A1(mai_mai_n148_), .B0(mai_mai_n106_), .B1(x4), .Y(mai_mai_n376_));
  NA3        m360(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n377_));
  NA2        m361(.A(mai_mai_n216_), .B(x0), .Y(mai_mai_n378_));
  OAI220     m362(.A0(mai_mai_n378_), .A1(mai_mai_n207_), .B0(mai_mai_n377_), .B1(mai_mai_n345_), .Y(mai_mai_n379_));
  AOI210     m363(.A0(mai_mai_n376_), .A1(mai_mai_n115_), .B0(mai_mai_n379_), .Y(mai_mai_n380_));
  AOI210     m364(.A0(mai_mai_n380_), .A1(mai_mai_n374_), .B0(mai_mai_n25_), .Y(mai_mai_n381_));
  NA3        m365(.A(mai_mai_n117_), .B(mai_mai_n216_), .C(x0), .Y(mai_mai_n382_));
  OAI210     m366(.A0(mai_mai_n193_), .A1(mai_mai_n63_), .B0(mai_mai_n203_), .Y(mai_mai_n383_));
  NA3        m367(.A(mai_mai_n196_), .B(mai_mai_n218_), .C(x8), .Y(mai_mai_n384_));
  AOI210     m368(.A0(mai_mai_n384_), .A1(mai_mai_n383_), .B0(mai_mai_n25_), .Y(mai_mai_n385_));
  NA2        m369(.A(mai_mai_n385_), .B(mai_mai_n148_), .Y(mai_mai_n386_));
  NA2        m370(.A(mai_mai_n386_), .B(mai_mai_n382_), .Y(mai_mai_n387_));
  OAI210     m371(.A0(mai_mai_n387_), .A1(mai_mai_n381_), .B0(x6), .Y(mai_mai_n388_));
  OAI210     m372(.A0(mai_mai_n162_), .A1(mai_mai_n45_), .B0(mai_mai_n132_), .Y(mai_mai_n389_));
  AOI210     m373(.A0(mai_mai_n37_), .A1(mai_mai_n31_), .B0(mai_mai_n389_), .Y(mai_mai_n390_));
  NO2        m374(.A(mai_mai_n151_), .B(x0), .Y(mai_mai_n391_));
  AOI220     m375(.A0(mai_mai_n391_), .A1(mai_mai_n216_), .B0(mai_mai_n193_), .B1(mai_mai_n151_), .Y(mai_mai_n392_));
  OAI210     m376(.A0(mai_mai_n392_), .A1(x8), .B0(mai_mai_n445_), .Y(mai_mai_n393_));
  NO3        m377(.A(mai_mai_n124_), .B(mai_mai_n292_), .C(x2), .Y(mai_mai_n394_));
  NOi21      m378(.An(mai_mai_n122_), .B(mai_mai_n177_), .Y(mai_mai_n395_));
  NO3        m379(.A(mai_mai_n395_), .B(mai_mai_n394_), .C(mai_mai_n18_), .Y(mai_mai_n396_));
  NO3        m380(.A(x9), .B(mai_mai_n151_), .C(x0), .Y(mai_mai_n397_));
  AOI220     m381(.A0(mai_mai_n397_), .A1(mai_mai_n237_), .B0(mai_mai_n356_), .B1(mai_mai_n151_), .Y(mai_mai_n398_));
  NA3        m382(.A(mai_mai_n398_), .B(mai_mai_n396_), .C(mai_mai_n47_), .Y(mai_mai_n399_));
  OAI210     m383(.A0(mai_mai_n393_), .A1(mai_mai_n390_), .B0(mai_mai_n399_), .Y(mai_mai_n400_));
  NOi31      m384(.An(mai_mai_n391_), .B(mai_mai_n31_), .C(x8), .Y(mai_mai_n401_));
  INV        m385(.A(mai_mai_n130_), .Y(mai_mai_n402_));
  NO3        m386(.A(mai_mai_n402_), .B(mai_mai_n122_), .C(mai_mai_n40_), .Y(mai_mai_n403_));
  NOi31      m387(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n404_));
  AOI220     m388(.A0(mai_mai_n404_), .A1(mai_mai_n340_), .B0(mai_mai_n123_), .B1(x3), .Y(mai_mai_n405_));
  AOI210     m389(.A0(mai_mai_n259_), .A1(mai_mai_n56_), .B0(mai_mai_n121_), .Y(mai_mai_n406_));
  OAI210     m390(.A0(mai_mai_n406_), .A1(x3), .B0(mai_mai_n405_), .Y(mai_mai_n407_));
  NO3        m391(.A(mai_mai_n407_), .B(mai_mai_n403_), .C(x2), .Y(mai_mai_n408_));
  OAI220     m392(.A0(mai_mai_n341_), .A1(mai_mai_n296_), .B0(mai_mai_n292_), .B1(mai_mai_n40_), .Y(mai_mai_n409_));
  INV        m393(.A(mai_mai_n377_), .Y(mai_mai_n410_));
  AOI220     m394(.A0(mai_mai_n410_), .A1(mai_mai_n88_), .B0(mai_mai_n409_), .B1(mai_mai_n151_), .Y(mai_mai_n411_));
  NO2        m395(.A(mai_mai_n411_), .B(mai_mai_n50_), .Y(mai_mai_n412_));
  NO3        m396(.A(mai_mai_n412_), .B(mai_mai_n408_), .C(mai_mai_n401_), .Y(mai_mai_n413_));
  AOI210     m397(.A0(mai_mai_n413_), .A1(mai_mai_n400_), .B0(mai_mai_n25_), .Y(mai_mai_n414_));
  NA4        m398(.A(mai_mai_n30_), .B(mai_mai_n88_), .C(x2), .D(mai_mai_n17_), .Y(mai_mai_n415_));
  NO3        m399(.A(mai_mai_n63_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n416_));
  NA2        m400(.A(mai_mai_n416_), .B(mai_mai_n260_), .Y(mai_mai_n417_));
  NO2        m401(.A(mai_mai_n417_), .B(mai_mai_n99_), .Y(mai_mai_n418_));
  NO3        m402(.A(mai_mai_n264_), .B(mai_mai_n172_), .C(mai_mai_n37_), .Y(mai_mai_n419_));
  OAI210     m403(.A0(mai_mai_n419_), .A1(mai_mai_n418_), .B0(x7), .Y(mai_mai_n420_));
  NA2        m404(.A(mai_mai_n221_), .B(x7), .Y(mai_mai_n421_));
  NA3        m405(.A(mai_mai_n421_), .B(mai_mai_n150_), .C(mai_mai_n131_), .Y(mai_mai_n422_));
  NA3        m406(.A(mai_mai_n422_), .B(mai_mai_n420_), .C(mai_mai_n415_), .Y(mai_mai_n423_));
  OAI210     m407(.A0(mai_mai_n423_), .A1(mai_mai_n414_), .B0(mai_mai_n35_), .Y(mai_mai_n424_));
  NO2        m408(.A(mai_mai_n397_), .B(mai_mai_n203_), .Y(mai_mai_n425_));
  NO4        m409(.A(mai_mai_n425_), .B(mai_mai_n72_), .C(x4), .D(mai_mai_n50_), .Y(mai_mai_n426_));
  NA2        m410(.A(mai_mai_n444_), .B(mai_mai_n173_), .Y(mai_mai_n427_));
  NO2        m411(.A(mai_mai_n159_), .B(mai_mai_n40_), .Y(mai_mai_n428_));
  NA2        m412(.A(x3), .B(mai_mai_n50_), .Y(mai_mai_n429_));
  AOI210     m413(.A0(mai_mai_n163_), .A1(mai_mai_n27_), .B0(mai_mai_n67_), .Y(mai_mai_n430_));
  OAI210     m414(.A0(mai_mai_n148_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n431_));
  NO3        m415(.A(mai_mai_n404_), .B(x3), .C(mai_mai_n50_), .Y(mai_mai_n432_));
  AOI210     m416(.A0(mai_mai_n432_), .A1(mai_mai_n431_), .B0(mai_mai_n430_), .Y(mai_mai_n433_));
  OAI210     m417(.A0(mai_mai_n152_), .A1(mai_mai_n429_), .B0(mai_mai_n433_), .Y(mai_mai_n434_));
  AOI220     m418(.A0(mai_mai_n434_), .A1(x0), .B0(mai_mai_n428_), .B1(mai_mai_n132_), .Y(mai_mai_n435_));
  AOI210     m419(.A0(mai_mai_n435_), .A1(mai_mai_n427_), .B0(mai_mai_n227_), .Y(mai_mai_n436_));
  INV        m420(.A(x5), .Y(mai_mai_n437_));
  NO4        m421(.A(mai_mai_n102_), .B(mai_mai_n437_), .C(mai_mai_n56_), .D(mai_mai_n31_), .Y(mai_mai_n438_));
  NO3        m422(.A(mai_mai_n438_), .B(mai_mai_n436_), .C(mai_mai_n426_), .Y(mai_mai_n439_));
  NA3        m423(.A(mai_mai_n439_), .B(mai_mai_n424_), .C(mai_mai_n388_), .Y(mai_mai_n440_));
  AOI210     m424(.A0(mai_mai_n371_), .A1(mai_mai_n25_), .B0(mai_mai_n440_), .Y(mai05));
  INV        m425(.A(mai_mai_n86_), .Y(mai_mai_n444_));
  INV        m426(.A(x1), .Y(mai_mai_n445_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  INV        u005(.A(men_men_n19_), .Y(men_men_n22_));
  NA2        u006(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n23_));
  INV        u007(.A(x5), .Y(men_men_n24_));
  NA2        u008(.A(x7), .B(x6), .Y(men_men_n25_));
  NA2        u009(.A(x8), .B(x3), .Y(men_men_n26_));
  NA2        u010(.A(x4), .B(x2), .Y(men_men_n27_));
  NO4        u011(.A(men_men_n27_), .B(men_men_n26_), .C(men_men_n25_), .D(men_men_n24_), .Y(men_men_n28_));
  NO2        u012(.A(men_men_n28_), .B(men_men_n23_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  NOi21      u015(.An(men_men_n22_), .B(men_men_n29_), .Y(men00));
  NO2        u016(.A(x1), .B(x0), .Y(men_men_n33_));
  INV        u017(.A(x6), .Y(men_men_n34_));
  NO2        u018(.A(men_men_n34_), .B(men_men_n24_), .Y(men_men_n35_));
  AN2        u019(.A(x8), .B(x7), .Y(men_men_n36_));
  NA3        u020(.A(men_men_n36_), .B(men_men_n35_), .C(men_men_n33_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  AOI210     u022(.A0(men_men_n37_), .A1(men_men_n22_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n35_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n50_));
  NA2        u034(.A(men_men_n50_), .B(men_men_n33_), .Y(men_men_n51_));
  INV        u035(.A(x2), .Y(men_men_n52_));
  NO2        u036(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  OAI210     u039(.A0(men_men_n51_), .A1(men_men_n31_), .B0(men_men_n55_), .Y(men_men_n56_));
  NO3        u040(.A(men_men_n56_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u041(.A(x8), .B(x7), .Y(men_men_n58_));
  NA2        u042(.A(men_men_n41_), .B(x1), .Y(men_men_n59_));
  INV        u043(.A(x9), .Y(men_men_n60_));
  NO2        u044(.A(men_men_n60_), .B(men_men_n34_), .Y(men_men_n61_));
  INV        u045(.A(men_men_n61_), .Y(men_men_n62_));
  NO3        u046(.A(men_men_n62_), .B(men_men_n59_), .C(men_men_n58_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n59_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  NO2        u051(.A(men_men_n67_), .B(x1), .Y(men_men_n68_));
  OA210      u052(.A0(men_men_n68_), .A1(men_men_n65_), .B0(men_men_n64_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n42_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n54_), .A1(men_men_n20_), .B0(men_men_n70_), .Y(men_men_n71_));
  NAi31      u055(.An(x1), .B(x9), .C(x5), .Y(men_men_n72_));
  OAI220     u056(.A0(men_men_n72_), .A1(men_men_n41_), .B0(men_men_n71_), .B1(men_men_n69_), .Y(men_men_n73_));
  OAI210     u057(.A0(men_men_n73_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n74_));
  NA2        u058(.A(men_men_n46_), .B(x2), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n76_));
  NA2        u060(.A(x5), .B(x3), .Y(men_men_n77_));
  NO2        u061(.A(x8), .B(x6), .Y(men_men_n78_));
  NO4        u062(.A(men_men_n78_), .B(men_men_n77_), .C(men_men_n64_), .D(men_men_n52_), .Y(men_men_n79_));
  NAi21      u063(.An(x4), .B(x3), .Y(men_men_n80_));
  INV        u064(.A(men_men_n80_), .Y(men_men_n81_));
  NO2        u065(.A(x4), .B(x2), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(x3), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n80_), .B(men_men_n18_), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n79_), .C(men_men_n76_), .Y(men_men_n85_));
  NO4        u069(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .D(x1), .Y(men_men_n86_));
  INV        u070(.A(x4), .Y(men_men_n87_));
  NA2        u071(.A(men_men_n86_), .B(men_men_n87_), .Y(men_men_n88_));
  NA2        u072(.A(x3), .B(men_men_n18_), .Y(men_men_n89_));
  NO2        u073(.A(men_men_n89_), .B(men_men_n24_), .Y(men_men_n90_));
  INV        u074(.A(x8), .Y(men_men_n91_));
  NA2        u075(.A(x2), .B(x1), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n91_), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n90_), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n94_), .B(men_men_n25_), .Y(men_men_n95_));
  AOI210     u079(.A0(men_men_n54_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n96_));
  OAI210     u080(.A0(men_men_n43_), .A1(men_men_n35_), .B0(men_men_n46_), .Y(men_men_n97_));
  NO3        u081(.A(men_men_n97_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n98_));
  NA2        u082(.A(x4), .B(men_men_n41_), .Y(men_men_n99_));
  NO2        u083(.A(men_men_n46_), .B(men_men_n52_), .Y(men_men_n100_));
  OAI210     u084(.A0(men_men_n100_), .A1(men_men_n41_), .B0(men_men_n18_), .Y(men_men_n101_));
  AOI210     u085(.A0(men_men_n99_), .A1(men_men_n50_), .B0(men_men_n101_), .Y(men_men_n102_));
  NO2        u086(.A(x3), .B(x2), .Y(men_men_n103_));
  NA3        u087(.A(men_men_n103_), .B(men_men_n25_), .C(men_men_n24_), .Y(men_men_n104_));
  AOI210     u088(.A0(x8), .A1(x6), .B0(men_men_n104_), .Y(men_men_n105_));
  NA2        u089(.A(men_men_n52_), .B(x1), .Y(men_men_n106_));
  OAI210     u090(.A0(men_men_n106_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n107_));
  NO4        u091(.A(men_men_n107_), .B(men_men_n105_), .C(men_men_n102_), .D(men_men_n98_), .Y(men_men_n108_));
  AO220      u092(.A0(men_men_n108_), .A1(men_men_n88_), .B0(men_men_n85_), .B1(men_men_n74_), .Y(men02));
  NO2        u093(.A(x3), .B(men_men_n52_), .Y(men_men_n110_));
  NO2        u094(.A(x8), .B(men_men_n18_), .Y(men_men_n111_));
  NA2        u095(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n41_), .B(x0), .Y(men_men_n113_));
  OAI210     u097(.A0(x4), .A1(men_men_n112_), .B0(men_men_n113_), .Y(men_men_n114_));
  AOI220     u098(.A0(men_men_n114_), .A1(men_men_n111_), .B0(men_men_n110_), .B1(x4), .Y(men_men_n115_));
  NO3        u099(.A(men_men_n115_), .B(x7), .C(x5), .Y(men_men_n116_));
  NA2        u100(.A(x9), .B(x2), .Y(men_men_n117_));
  OR2        u101(.A(x8), .B(x0), .Y(men_men_n118_));
  INV        u102(.A(men_men_n118_), .Y(men_men_n119_));
  NAi21      u103(.An(x2), .B(x8), .Y(men_men_n120_));
  INV        u104(.A(men_men_n120_), .Y(men_men_n121_));
  NO2        u105(.A(x4), .B(x1), .Y(men_men_n122_));
  NA3        u106(.A(men_men_n122_), .B(x0), .C(men_men_n58_), .Y(men_men_n123_));
  NOi21      u107(.An(x0), .B(x1), .Y(men_men_n124_));
  NO3        u108(.A(x9), .B(x8), .C(x7), .Y(men_men_n125_));
  NOi21      u109(.An(x0), .B(x4), .Y(men_men_n126_));
  NAi21      u110(.An(x8), .B(x7), .Y(men_men_n127_));
  NO2        u111(.A(men_men_n127_), .B(men_men_n60_), .Y(men_men_n128_));
  AOI220     u112(.A0(men_men_n128_), .A1(men_men_n126_), .B0(men_men_n125_), .B1(men_men_n124_), .Y(men_men_n129_));
  AOI210     u113(.A0(men_men_n129_), .A1(men_men_n123_), .B0(men_men_n77_), .Y(men_men_n130_));
  NO2        u114(.A(x5), .B(men_men_n46_), .Y(men_men_n131_));
  NA2        u115(.A(x2), .B(men_men_n18_), .Y(men_men_n132_));
  AOI210     u116(.A0(men_men_n132_), .A1(men_men_n106_), .B0(men_men_n113_), .Y(men_men_n133_));
  OAI210     u117(.A0(men_men_n133_), .A1(men_men_n33_), .B0(men_men_n131_), .Y(men_men_n134_));
  NAi21      u118(.An(x0), .B(x4), .Y(men_men_n135_));
  NO2        u119(.A(men_men_n135_), .B(x1), .Y(men_men_n136_));
  NO2        u120(.A(x7), .B(x0), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n82_), .B(men_men_n100_), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n138_), .B(x3), .Y(men_men_n139_));
  OAI210     u123(.A0(men_men_n137_), .A1(men_men_n136_), .B0(men_men_n139_), .Y(men_men_n140_));
  NA2        u124(.A(x5), .B(x0), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n46_), .B(x2), .Y(men_men_n142_));
  NA3        u126(.A(men_men_n140_), .B(men_men_n134_), .C(men_men_n34_), .Y(men_men_n143_));
  NO3        u127(.A(men_men_n143_), .B(men_men_n130_), .C(men_men_n116_), .Y(men_men_n144_));
  NO3        u128(.A(men_men_n77_), .B(men_men_n75_), .C(men_men_n23_), .Y(men_men_n145_));
  NO2        u129(.A(men_men_n27_), .B(men_men_n24_), .Y(men_men_n146_));
  AOI220     u130(.A0(men_men_n124_), .A1(men_men_n146_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n147_), .B(men_men_n58_), .C(men_men_n60_), .Y(men_men_n148_));
  NA2        u132(.A(x7), .B(x3), .Y(men_men_n149_));
  NO2        u133(.A(men_men_n99_), .B(x5), .Y(men_men_n150_));
  NO2        u134(.A(x9), .B(x7), .Y(men_men_n151_));
  NOi21      u135(.An(x8), .B(x0), .Y(men_men_n152_));
  OA210      u136(.A0(men_men_n151_), .A1(x1), .B0(men_men_n152_), .Y(men_men_n153_));
  NO2        u137(.A(men_men_n41_), .B(x2), .Y(men_men_n154_));
  INV        u138(.A(x7), .Y(men_men_n155_));
  NA2        u139(.A(men_men_n155_), .B(men_men_n18_), .Y(men_men_n156_));
  AOI220     u140(.A0(men_men_n156_), .A1(men_men_n154_), .B0(men_men_n110_), .B1(men_men_n36_), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n24_), .B(x4), .Y(men_men_n158_));
  NO2        u142(.A(men_men_n158_), .B(men_men_n126_), .Y(men_men_n159_));
  NO2        u143(.A(men_men_n159_), .B(men_men_n157_), .Y(men_men_n160_));
  AOI210     u144(.A0(men_men_n153_), .A1(men_men_n150_), .B0(men_men_n160_), .Y(men_men_n161_));
  OAI210     u145(.A0(men_men_n149_), .A1(men_men_n48_), .B0(men_men_n161_), .Y(men_men_n162_));
  NA2        u146(.A(x5), .B(x1), .Y(men_men_n163_));
  INV        u147(.A(men_men_n163_), .Y(men_men_n164_));
  AOI210     u148(.A0(men_men_n164_), .A1(men_men_n126_), .B0(men_men_n34_), .Y(men_men_n165_));
  NO2        u149(.A(men_men_n60_), .B(men_men_n91_), .Y(men_men_n166_));
  NAi21      u150(.An(x2), .B(x7), .Y(men_men_n167_));
  NO3        u151(.A(men_men_n167_), .B(men_men_n166_), .C(men_men_n46_), .Y(men_men_n168_));
  NA2        u152(.A(men_men_n168_), .B(men_men_n65_), .Y(men_men_n169_));
  NAi31      u153(.An(men_men_n77_), .B(men_men_n36_), .C(men_men_n33_), .Y(men_men_n170_));
  NA3        u154(.A(men_men_n170_), .B(men_men_n169_), .C(men_men_n165_), .Y(men_men_n171_));
  NO4        u155(.A(men_men_n171_), .B(men_men_n162_), .C(men_men_n148_), .D(men_men_n145_), .Y(men_men_n172_));
  NO2        u156(.A(men_men_n172_), .B(men_men_n144_), .Y(men_men_n173_));
  NO2        u157(.A(men_men_n141_), .B(men_men_n138_), .Y(men_men_n174_));
  NA2        u158(.A(men_men_n24_), .B(men_men_n18_), .Y(men_men_n175_));
  NA2        u159(.A(men_men_n24_), .B(men_men_n17_), .Y(men_men_n176_));
  NA3        u160(.A(men_men_n176_), .B(men_men_n175_), .C(men_men_n23_), .Y(men_men_n177_));
  AN2        u161(.A(men_men_n177_), .B(men_men_n142_), .Y(men_men_n178_));
  NA2        u162(.A(x8), .B(x0), .Y(men_men_n179_));
  NO2        u163(.A(men_men_n155_), .B(men_men_n24_), .Y(men_men_n180_));
  NO2        u164(.A(men_men_n124_), .B(x4), .Y(men_men_n181_));
  NA2        u165(.A(men_men_n181_), .B(men_men_n180_), .Y(men_men_n182_));
  AOI210     u166(.A0(men_men_n179_), .A1(men_men_n132_), .B0(men_men_n182_), .Y(men_men_n183_));
  NA2        u167(.A(x2), .B(x0), .Y(men_men_n184_));
  NA2        u168(.A(x4), .B(x1), .Y(men_men_n185_));
  NAi21      u169(.An(men_men_n122_), .B(men_men_n185_), .Y(men_men_n186_));
  NOi31      u170(.An(men_men_n186_), .B(men_men_n158_), .C(men_men_n184_), .Y(men_men_n187_));
  NO4        u171(.A(men_men_n187_), .B(men_men_n183_), .C(men_men_n178_), .D(men_men_n174_), .Y(men_men_n188_));
  NO2        u172(.A(men_men_n188_), .B(men_men_n41_), .Y(men_men_n189_));
  NO2        u173(.A(men_men_n177_), .B(men_men_n75_), .Y(men_men_n190_));
  INV        u174(.A(men_men_n131_), .Y(men_men_n191_));
  NO2        u175(.A(men_men_n106_), .B(men_men_n17_), .Y(men_men_n192_));
  AOI210     u176(.A0(men_men_n33_), .A1(men_men_n91_), .B0(men_men_n192_), .Y(men_men_n193_));
  NO3        u177(.A(men_men_n193_), .B(men_men_n191_), .C(x7), .Y(men_men_n194_));
  NA3        u178(.A(men_men_n186_), .B(men_men_n191_), .C(men_men_n40_), .Y(men_men_n195_));
  OAI210     u179(.A0(men_men_n176_), .A1(men_men_n138_), .B0(men_men_n195_), .Y(men_men_n196_));
  NO3        u180(.A(men_men_n196_), .B(men_men_n194_), .C(men_men_n190_), .Y(men_men_n197_));
  NO2        u181(.A(men_men_n197_), .B(x3), .Y(men_men_n198_));
  NO3        u182(.A(men_men_n198_), .B(men_men_n189_), .C(men_men_n173_), .Y(men03));
  NO2        u183(.A(men_men_n46_), .B(x3), .Y(men_men_n200_));
  NO2        u184(.A(x6), .B(men_men_n24_), .Y(men_men_n201_));
  NO2        u185(.A(men_men_n52_), .B(x1), .Y(men_men_n202_));
  OAI210     u186(.A0(men_men_n202_), .A1(men_men_n24_), .B0(men_men_n61_), .Y(men_men_n203_));
  NO2        u187(.A(men_men_n203_), .B(men_men_n17_), .Y(men_men_n204_));
  NA2        u188(.A(men_men_n204_), .B(men_men_n200_), .Y(men_men_n205_));
  NA2        u189(.A(x6), .B(men_men_n24_), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n206_), .B(x4), .Y(men_men_n207_));
  NO2        u191(.A(men_men_n18_), .B(x0), .Y(men_men_n208_));
  NA2        u192(.A(x3), .B(men_men_n17_), .Y(men_men_n209_));
  NO2        u193(.A(men_men_n209_), .B(men_men_n206_), .Y(men_men_n210_));
  NA2        u194(.A(x9), .B(men_men_n52_), .Y(men_men_n211_));
  NA2        u195(.A(men_men_n211_), .B(x4), .Y(men_men_n212_));
  NA2        u196(.A(men_men_n206_), .B(men_men_n80_), .Y(men_men_n213_));
  AOI210     u197(.A0(men_men_n24_), .A1(x3), .B0(men_men_n184_), .Y(men_men_n214_));
  AOI220     u198(.A0(men_men_n214_), .A1(men_men_n213_), .B0(men_men_n212_), .B1(men_men_n210_), .Y(men_men_n215_));
  NO2        u199(.A(x5), .B(x1), .Y(men_men_n216_));
  AOI220     u200(.A0(men_men_n216_), .A1(men_men_n17_), .B0(men_men_n103_), .B1(x5), .Y(men_men_n217_));
  NO2        u201(.A(men_men_n209_), .B(men_men_n175_), .Y(men_men_n218_));
  NO3        u202(.A(x3), .B(x2), .C(x1), .Y(men_men_n219_));
  NO2        u203(.A(men_men_n219_), .B(men_men_n218_), .Y(men_men_n220_));
  OAI210     u204(.A0(men_men_n217_), .A1(men_men_n62_), .B0(men_men_n220_), .Y(men_men_n221_));
  NA2        u205(.A(men_men_n221_), .B(men_men_n46_), .Y(men_men_n222_));
  NA3        u206(.A(men_men_n222_), .B(men_men_n215_), .C(men_men_n205_), .Y(men_men_n223_));
  NO2        u207(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n224_));
  NA2        u208(.A(men_men_n224_), .B(men_men_n19_), .Y(men_men_n225_));
  NO2        u209(.A(x3), .B(men_men_n17_), .Y(men_men_n226_));
  NO2        u210(.A(men_men_n226_), .B(x6), .Y(men_men_n227_));
  NOi21      u211(.An(men_men_n82_), .B(men_men_n227_), .Y(men_men_n228_));
  NA2        u212(.A(men_men_n60_), .B(men_men_n91_), .Y(men_men_n229_));
  NO2        u213(.A(men_men_n228_), .B(men_men_n155_), .Y(men_men_n230_));
  OR2        u214(.A(men_men_n230_), .B(men_men_n180_), .Y(men_men_n231_));
  NA2        u215(.A(men_men_n41_), .B(men_men_n52_), .Y(men_men_n232_));
  OAI210     u216(.A0(men_men_n232_), .A1(men_men_n24_), .B0(men_men_n176_), .Y(men_men_n233_));
  NO3        u217(.A(men_men_n185_), .B(men_men_n60_), .C(x6), .Y(men_men_n234_));
  AOI220     u218(.A0(men_men_n234_), .A1(men_men_n233_), .B0(men_men_n142_), .B1(men_men_n90_), .Y(men_men_n235_));
  NA2        u219(.A(x6), .B(men_men_n46_), .Y(men_men_n236_));
  OAI210     u220(.A0(men_men_n119_), .A1(men_men_n78_), .B0(x4), .Y(men_men_n237_));
  AOI210     u221(.A0(men_men_n237_), .A1(men_men_n236_), .B0(men_men_n77_), .Y(men_men_n238_));
  NO2        u222(.A(men_men_n60_), .B(x6), .Y(men_men_n239_));
  NO2        u223(.A(men_men_n163_), .B(men_men_n41_), .Y(men_men_n240_));
  OAI210     u224(.A0(men_men_n240_), .A1(men_men_n218_), .B0(men_men_n239_), .Y(men_men_n241_));
  NA2        u225(.A(men_men_n201_), .B(men_men_n136_), .Y(men_men_n242_));
  NA3        u226(.A(men_men_n209_), .B(men_men_n131_), .C(x6), .Y(men_men_n243_));
  OAI210     u227(.A0(men_men_n91_), .A1(men_men_n34_), .B0(men_men_n65_), .Y(men_men_n244_));
  NA4        u228(.A(men_men_n244_), .B(men_men_n243_), .C(men_men_n242_), .D(men_men_n241_), .Y(men_men_n245_));
  OAI210     u229(.A0(men_men_n245_), .A1(men_men_n238_), .B0(x2), .Y(men_men_n246_));
  NA3        u230(.A(men_men_n246_), .B(men_men_n235_), .C(men_men_n231_), .Y(men_men_n247_));
  AOI210     u231(.A0(men_men_n223_), .A1(x8), .B0(men_men_n247_), .Y(men_men_n248_));
  NO2        u232(.A(men_men_n91_), .B(x3), .Y(men_men_n249_));
  NA2        u233(.A(men_men_n249_), .B(men_men_n207_), .Y(men_men_n250_));
  NO3        u234(.A(men_men_n89_), .B(men_men_n78_), .C(men_men_n24_), .Y(men_men_n251_));
  AOI210     u235(.A0(men_men_n227_), .A1(men_men_n158_), .B0(men_men_n251_), .Y(men_men_n252_));
  AOI210     u236(.A0(men_men_n252_), .A1(men_men_n250_), .B0(x2), .Y(men_men_n253_));
  NO2        u237(.A(x4), .B(men_men_n52_), .Y(men_men_n254_));
  AOI220     u238(.A0(men_men_n207_), .A1(men_men_n192_), .B0(men_men_n254_), .B1(men_men_n65_), .Y(men_men_n255_));
  NA2        u239(.A(men_men_n60_), .B(x6), .Y(men_men_n256_));
  NA3        u240(.A(men_men_n24_), .B(x3), .C(x2), .Y(men_men_n257_));
  AOI210     u241(.A0(men_men_n257_), .A1(men_men_n141_), .B0(men_men_n256_), .Y(men_men_n258_));
  NA2        u242(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n259_));
  NO2        u243(.A(men_men_n259_), .B(men_men_n24_), .Y(men_men_n260_));
  OAI210     u244(.A0(men_men_n260_), .A1(men_men_n258_), .B0(men_men_n122_), .Y(men_men_n261_));
  NA2        u245(.A(men_men_n209_), .B(x6), .Y(men_men_n262_));
  NO2        u246(.A(men_men_n209_), .B(x6), .Y(men_men_n263_));
  NA2        u247(.A(men_men_n262_), .B(men_men_n146_), .Y(men_men_n264_));
  NA4        u248(.A(men_men_n264_), .B(men_men_n261_), .C(men_men_n255_), .D(men_men_n155_), .Y(men_men_n265_));
  NA2        u249(.A(men_men_n201_), .B(men_men_n226_), .Y(men_men_n266_));
  NO2        u250(.A(x9), .B(x6), .Y(men_men_n267_));
  NO2        u251(.A(men_men_n141_), .B(men_men_n18_), .Y(men_men_n268_));
  NAi21      u252(.An(men_men_n268_), .B(men_men_n257_), .Y(men_men_n269_));
  NAi21      u253(.An(x1), .B(x4), .Y(men_men_n270_));
  AOI210     u254(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n271_));
  OAI210     u255(.A0(men_men_n141_), .A1(x3), .B0(men_men_n271_), .Y(men_men_n272_));
  AOI220     u256(.A0(men_men_n272_), .A1(men_men_n270_), .B0(men_men_n269_), .B1(men_men_n267_), .Y(men_men_n273_));
  NA2        u257(.A(men_men_n273_), .B(men_men_n266_), .Y(men_men_n274_));
  NA2        u258(.A(men_men_n60_), .B(x2), .Y(men_men_n275_));
  NO2        u259(.A(men_men_n275_), .B(men_men_n266_), .Y(men_men_n276_));
  NO3        u260(.A(x9), .B(x6), .C(x0), .Y(men_men_n277_));
  NA2        u261(.A(men_men_n106_), .B(men_men_n24_), .Y(men_men_n278_));
  NA2        u262(.A(x6), .B(x2), .Y(men_men_n279_));
  NO2        u263(.A(men_men_n279_), .B(men_men_n175_), .Y(men_men_n280_));
  AOI210     u264(.A0(men_men_n278_), .A1(men_men_n277_), .B0(men_men_n280_), .Y(men_men_n281_));
  OAI220     u265(.A0(men_men_n281_), .A1(men_men_n41_), .B0(men_men_n181_), .B1(men_men_n44_), .Y(men_men_n282_));
  OAI210     u266(.A0(men_men_n282_), .A1(men_men_n276_), .B0(men_men_n274_), .Y(men_men_n283_));
  NO2        u267(.A(x3), .B(men_men_n206_), .Y(men_men_n284_));
  NA2        u268(.A(x4), .B(x0), .Y(men_men_n285_));
  NO3        u269(.A(men_men_n72_), .B(men_men_n285_), .C(x6), .Y(men_men_n286_));
  AOI210     u270(.A0(men_men_n284_), .A1(men_men_n40_), .B0(men_men_n286_), .Y(men_men_n287_));
  AOI210     u271(.A0(men_men_n287_), .A1(men_men_n283_), .B0(x8), .Y(men_men_n288_));
  INV        u272(.A(men_men_n256_), .Y(men_men_n289_));
  OAI210     u273(.A0(men_men_n268_), .A1(men_men_n216_), .B0(men_men_n289_), .Y(men_men_n290_));
  OAI210     u274(.A0(x0), .A1(x4), .B0(men_men_n20_), .Y(men_men_n291_));
  AOI210     u275(.A0(men_men_n291_), .A1(men_men_n290_), .B0(men_men_n232_), .Y(men_men_n292_));
  NO4        u276(.A(men_men_n292_), .B(men_men_n288_), .C(men_men_n265_), .D(men_men_n253_), .Y(men_men_n293_));
  NO2        u277(.A(men_men_n166_), .B(x1), .Y(men_men_n294_));
  NO3        u278(.A(men_men_n294_), .B(x3), .C(men_men_n34_), .Y(men_men_n295_));
  OAI210     u279(.A0(men_men_n295_), .A1(men_men_n263_), .B0(x2), .Y(men_men_n296_));
  OAI210     u280(.A0(x0), .A1(x6), .B0(men_men_n42_), .Y(men_men_n297_));
  AOI210     u281(.A0(men_men_n297_), .A1(men_men_n296_), .B0(men_men_n191_), .Y(men_men_n298_));
  NOi21      u282(.An(men_men_n279_), .B(men_men_n17_), .Y(men_men_n299_));
  NA3        u283(.A(men_men_n299_), .B(men_men_n216_), .C(men_men_n38_), .Y(men_men_n300_));
  AOI210     u284(.A0(men_men_n34_), .A1(men_men_n52_), .B0(x0), .Y(men_men_n301_));
  NA3        u285(.A(men_men_n301_), .B(men_men_n164_), .C(men_men_n31_), .Y(men_men_n302_));
  NA2        u286(.A(x3), .B(x2), .Y(men_men_n303_));
  AOI220     u287(.A0(men_men_n303_), .A1(men_men_n232_), .B0(men_men_n302_), .B1(men_men_n300_), .Y(men_men_n304_));
  NAi21      u288(.An(x4), .B(x0), .Y(men_men_n305_));
  NO3        u289(.A(men_men_n305_), .B(men_men_n42_), .C(x2), .Y(men_men_n306_));
  OAI210     u290(.A0(x6), .A1(men_men_n18_), .B0(men_men_n306_), .Y(men_men_n307_));
  OAI220     u291(.A0(men_men_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n308_));
  NO2        u292(.A(x9), .B(x8), .Y(men_men_n309_));
  NA3        u293(.A(men_men_n309_), .B(men_men_n34_), .C(men_men_n52_), .Y(men_men_n310_));
  OAI210     u294(.A0(men_men_n301_), .A1(men_men_n299_), .B0(men_men_n310_), .Y(men_men_n311_));
  AOI220     u295(.A0(men_men_n311_), .A1(men_men_n81_), .B0(men_men_n308_), .B1(men_men_n30_), .Y(men_men_n312_));
  AOI210     u296(.A0(men_men_n312_), .A1(men_men_n307_), .B0(men_men_n24_), .Y(men_men_n313_));
  NA3        u297(.A(men_men_n34_), .B(x1), .C(men_men_n17_), .Y(men_men_n314_));
  OAI210     u298(.A0(men_men_n301_), .A1(men_men_n299_), .B0(men_men_n314_), .Y(men_men_n315_));
  INV        u299(.A(men_men_n218_), .Y(men_men_n316_));
  NA2        u300(.A(men_men_n34_), .B(men_men_n41_), .Y(men_men_n317_));
  OR2        u301(.A(men_men_n317_), .B(men_men_n285_), .Y(men_men_n318_));
  OAI220     u302(.A0(men_men_n318_), .A1(men_men_n163_), .B0(men_men_n236_), .B1(men_men_n316_), .Y(men_men_n319_));
  AO210      u303(.A0(men_men_n315_), .A1(men_men_n150_), .B0(men_men_n319_), .Y(men_men_n320_));
  NO4        u304(.A(men_men_n320_), .B(men_men_n313_), .C(men_men_n304_), .D(men_men_n298_), .Y(men_men_n321_));
  OAI210     u305(.A0(men_men_n293_), .A1(men_men_n248_), .B0(men_men_n321_), .Y(men04));
  OAI210     u306(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n323_));
  NA3        u307(.A(men_men_n323_), .B(men_men_n277_), .C(men_men_n83_), .Y(men_men_n324_));
  NO2        u308(.A(x2), .B(x1), .Y(men_men_n325_));
  OAI210     u309(.A0(men_men_n259_), .A1(men_men_n325_), .B0(men_men_n34_), .Y(men_men_n326_));
  NO2        u310(.A(men_men_n325_), .B(men_men_n305_), .Y(men_men_n327_));
  AOI210     u311(.A0(men_men_n60_), .A1(x4), .B0(men_men_n112_), .Y(men_men_n328_));
  OAI210     u312(.A0(men_men_n328_), .A1(men_men_n327_), .B0(men_men_n249_), .Y(men_men_n329_));
  NO2        u313(.A(men_men_n275_), .B(men_men_n89_), .Y(men_men_n330_));
  NO2        u314(.A(men_men_n330_), .B(men_men_n34_), .Y(men_men_n331_));
  NO2        u315(.A(men_men_n303_), .B(men_men_n208_), .Y(men_men_n332_));
  NA2        u316(.A(x9), .B(x0), .Y(men_men_n333_));
  AOI210     u317(.A0(men_men_n89_), .A1(men_men_n75_), .B0(men_men_n333_), .Y(men_men_n334_));
  OAI210     u318(.A0(men_men_n334_), .A1(men_men_n332_), .B0(men_men_n91_), .Y(men_men_n335_));
  NA3        u319(.A(men_men_n335_), .B(men_men_n331_), .C(men_men_n329_), .Y(men_men_n336_));
  NA2        u320(.A(men_men_n336_), .B(men_men_n326_), .Y(men_men_n337_));
  NO2        u321(.A(men_men_n211_), .B(men_men_n113_), .Y(men_men_n338_));
  NO3        u322(.A(men_men_n256_), .B(men_men_n120_), .C(men_men_n18_), .Y(men_men_n339_));
  NO2        u323(.A(men_men_n339_), .B(men_men_n338_), .Y(men_men_n340_));
  NOi21      u324(.An(men_men_n152_), .B(men_men_n132_), .Y(men_men_n341_));
  AOI210     u325(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n342_));
  OAI220     u326(.A0(men_men_n342_), .A1(men_men_n317_), .B0(men_men_n275_), .B1(men_men_n314_), .Y(men_men_n343_));
  AOI210     u327(.A0(men_men_n341_), .A1(men_men_n61_), .B0(men_men_n343_), .Y(men_men_n344_));
  NA2        u328(.A(x2), .B(men_men_n17_), .Y(men_men_n345_));
  NA2        u329(.A(men_men_n330_), .B(men_men_n91_), .Y(men_men_n346_));
  NA3        u330(.A(men_men_n346_), .B(men_men_n344_), .C(men_men_n340_), .Y(men_men_n347_));
  OAI210     u331(.A0(men_men_n111_), .A1(x3), .B0(men_men_n306_), .Y(men_men_n348_));
  NA2        u332(.A(men_men_n348_), .B(men_men_n155_), .Y(men_men_n349_));
  AOI210     u333(.A0(men_men_n347_), .A1(x4), .B0(men_men_n349_), .Y(men_men_n350_));
  NA3        u334(.A(men_men_n327_), .B(men_men_n211_), .C(men_men_n91_), .Y(men_men_n351_));
  NOi21      u335(.An(x4), .B(x0), .Y(men_men_n352_));
  XO2        u336(.A(x4), .B(x0), .Y(men_men_n353_));
  OAI210     u337(.A0(men_men_n353_), .A1(men_men_n117_), .B0(men_men_n270_), .Y(men_men_n354_));
  AOI220     u338(.A0(men_men_n354_), .A1(x8), .B0(men_men_n352_), .B1(men_men_n92_), .Y(men_men_n355_));
  AOI210     u339(.A0(men_men_n355_), .A1(men_men_n351_), .B0(x3), .Y(men_men_n356_));
  INV        u340(.A(men_men_n92_), .Y(men_men_n357_));
  NO2        u341(.A(men_men_n91_), .B(x4), .Y(men_men_n358_));
  AOI220     u342(.A0(men_men_n358_), .A1(men_men_n42_), .B0(men_men_n126_), .B1(men_men_n357_), .Y(men_men_n359_));
  NO3        u343(.A(men_men_n353_), .B(men_men_n166_), .C(x2), .Y(men_men_n360_));
  NO3        u344(.A(men_men_n229_), .B(men_men_n27_), .C(men_men_n23_), .Y(men_men_n361_));
  NO2        u345(.A(men_men_n361_), .B(men_men_n360_), .Y(men_men_n362_));
  NA4        u346(.A(men_men_n362_), .B(men_men_n359_), .C(men_men_n225_), .D(x6), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n184_), .B(men_men_n91_), .Y(men_men_n364_));
  NO2        u348(.A(men_men_n41_), .B(x0), .Y(men_men_n365_));
  OR2        u349(.A(men_men_n358_), .B(men_men_n365_), .Y(men_men_n366_));
  NO2        u350(.A(men_men_n152_), .B(men_men_n106_), .Y(men_men_n367_));
  AOI220     u351(.A0(men_men_n367_), .A1(men_men_n366_), .B0(men_men_n364_), .B1(men_men_n59_), .Y(men_men_n368_));
  NO2        u352(.A(men_men_n152_), .B(men_men_n80_), .Y(men_men_n369_));
  NO2        u353(.A(men_men_n33_), .B(x2), .Y(men_men_n370_));
  NOi21      u354(.An(men_men_n122_), .B(men_men_n26_), .Y(men_men_n371_));
  AOI210     u355(.A0(men_men_n370_), .A1(men_men_n369_), .B0(men_men_n371_), .Y(men_men_n372_));
  OAI210     u356(.A0(men_men_n368_), .A1(men_men_n60_), .B0(men_men_n372_), .Y(men_men_n373_));
  OAI220     u357(.A0(men_men_n373_), .A1(x6), .B0(men_men_n363_), .B1(men_men_n356_), .Y(men_men_n374_));
  OAI210     u358(.A0(men_men_n61_), .A1(men_men_n46_), .B0(men_men_n40_), .Y(men_men_n375_));
  OAI210     u359(.A0(men_men_n375_), .A1(men_men_n91_), .B0(men_men_n318_), .Y(men_men_n376_));
  AOI210     u360(.A0(men_men_n376_), .A1(men_men_n18_), .B0(men_men_n155_), .Y(men_men_n377_));
  AO220      u361(.A0(men_men_n377_), .A1(men_men_n374_), .B0(men_men_n350_), .B1(men_men_n337_), .Y(men_men_n378_));
  NA2        u362(.A(men_men_n219_), .B(men_men_n47_), .Y(men_men_n379_));
  NA3        u363(.A(men_men_n379_), .B(men_men_n378_), .C(men_men_n324_), .Y(men_men_n380_));
  AOI210     u364(.A0(men_men_n202_), .A1(x8), .B0(men_men_n111_), .Y(men_men_n381_));
  NA2        u365(.A(men_men_n381_), .B(men_men_n345_), .Y(men_men_n382_));
  NA3        u366(.A(men_men_n382_), .B(men_men_n200_), .C(men_men_n155_), .Y(men_men_n383_));
  NA3        u367(.A(x7), .B(x3), .C(x0), .Y(men_men_n384_));
  NO2        u368(.A(men_men_n384_), .B(men_men_n357_), .Y(men_men_n385_));
  INV        u369(.A(men_men_n385_), .Y(men_men_n386_));
  AOI210     u370(.A0(men_men_n386_), .A1(men_men_n383_), .B0(men_men_n24_), .Y(men_men_n387_));
  NA3        u371(.A(men_men_n121_), .B(men_men_n224_), .C(x0), .Y(men_men_n388_));
  OAI210     u372(.A0(men_men_n200_), .A1(men_men_n66_), .B0(men_men_n208_), .Y(men_men_n389_));
  NA3        u373(.A(men_men_n202_), .B(men_men_n226_), .C(x8), .Y(men_men_n390_));
  AOI210     u374(.A0(men_men_n390_), .A1(men_men_n389_), .B0(men_men_n24_), .Y(men_men_n391_));
  AOI210     u375(.A0(men_men_n120_), .A1(men_men_n118_), .B0(men_men_n40_), .Y(men_men_n392_));
  NOi31      u376(.An(men_men_n392_), .B(men_men_n365_), .C(men_men_n185_), .Y(men_men_n393_));
  OAI210     u377(.A0(men_men_n393_), .A1(men_men_n391_), .B0(men_men_n151_), .Y(men_men_n394_));
  NAi31      u378(.An(men_men_n48_), .B(men_men_n294_), .C(men_men_n180_), .Y(men_men_n395_));
  NA3        u379(.A(men_men_n395_), .B(men_men_n394_), .C(men_men_n388_), .Y(men_men_n396_));
  OAI210     u380(.A0(men_men_n396_), .A1(men_men_n387_), .B0(x6), .Y(men_men_n397_));
  INV        u381(.A(men_men_n137_), .Y(men_men_n398_));
  NA3        u382(.A(men_men_n53_), .B(men_men_n36_), .C(men_men_n30_), .Y(men_men_n399_));
  AOI220     u383(.A0(men_men_n399_), .A1(men_men_n398_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n400_));
  NO2        u384(.A(men_men_n155_), .B(x0), .Y(men_men_n401_));
  AOI220     u385(.A0(men_men_n401_), .A1(men_men_n224_), .B0(men_men_n200_), .B1(men_men_n155_), .Y(men_men_n402_));
  AOI210     u386(.A0(men_men_n128_), .A1(men_men_n254_), .B0(x1), .Y(men_men_n403_));
  OAI210     u387(.A0(men_men_n402_), .A1(x8), .B0(men_men_n403_), .Y(men_men_n404_));
  NAi31      u388(.An(x2), .B(x8), .C(x0), .Y(men_men_n405_));
  OAI210     u389(.A0(men_men_n405_), .A1(x4), .B0(men_men_n167_), .Y(men_men_n406_));
  NA3        u390(.A(men_men_n406_), .B(men_men_n149_), .C(x9), .Y(men_men_n407_));
  NO4        u391(.A(men_men_n127_), .B(men_men_n305_), .C(x9), .D(x2), .Y(men_men_n408_));
  NOi21      u392(.An(men_men_n125_), .B(men_men_n184_), .Y(men_men_n409_));
  NO3        u393(.A(men_men_n409_), .B(men_men_n408_), .C(men_men_n18_), .Y(men_men_n410_));
  NO3        u394(.A(x9), .B(men_men_n155_), .C(x0), .Y(men_men_n411_));
  AOI220     u395(.A0(men_men_n411_), .A1(men_men_n249_), .B0(men_men_n369_), .B1(men_men_n155_), .Y(men_men_n412_));
  NA4        u396(.A(men_men_n412_), .B(men_men_n410_), .C(men_men_n407_), .D(men_men_n48_), .Y(men_men_n413_));
  OAI210     u397(.A0(men_men_n404_), .A1(men_men_n400_), .B0(men_men_n413_), .Y(men_men_n414_));
  NOi31      u398(.An(men_men_n401_), .B(men_men_n31_), .C(x8), .Y(men_men_n415_));
  AOI210     u399(.A0(men_men_n36_), .A1(x9), .B0(men_men_n135_), .Y(men_men_n416_));
  NO3        u400(.A(men_men_n416_), .B(men_men_n125_), .C(men_men_n41_), .Y(men_men_n417_));
  AOI210     u401(.A0(men_men_n270_), .A1(men_men_n58_), .B0(men_men_n124_), .Y(men_men_n418_));
  NO2        u402(.A(men_men_n418_), .B(x3), .Y(men_men_n419_));
  NO3        u403(.A(men_men_n419_), .B(men_men_n417_), .C(x2), .Y(men_men_n420_));
  OAI220     u404(.A0(men_men_n353_), .A1(men_men_n309_), .B0(men_men_n305_), .B1(men_men_n41_), .Y(men_men_n421_));
  AOI210     u405(.A0(x9), .A1(men_men_n46_), .B0(men_men_n384_), .Y(men_men_n422_));
  AOI220     u406(.A0(men_men_n422_), .A1(men_men_n91_), .B0(men_men_n421_), .B1(men_men_n155_), .Y(men_men_n423_));
  NO2        u407(.A(men_men_n423_), .B(men_men_n52_), .Y(men_men_n424_));
  NO3        u408(.A(men_men_n424_), .B(men_men_n420_), .C(men_men_n415_), .Y(men_men_n425_));
  AOI210     u409(.A0(men_men_n425_), .A1(men_men_n414_), .B0(men_men_n24_), .Y(men_men_n426_));
  NO3        u410(.A(men_men_n60_), .B(x4), .C(x1), .Y(men_men_n427_));
  NO3        u411(.A(men_men_n66_), .B(men_men_n18_), .C(x0), .Y(men_men_n428_));
  AOI220     u412(.A0(men_men_n428_), .A1(men_men_n271_), .B0(men_men_n427_), .B1(men_men_n392_), .Y(men_men_n429_));
  NO2        u413(.A(men_men_n429_), .B(men_men_n103_), .Y(men_men_n430_));
  NA2        u414(.A(men_men_n430_), .B(x7), .Y(men_men_n431_));
  NA2        u415(.A(men_men_n229_), .B(x7), .Y(men_men_n432_));
  NA3        u416(.A(men_men_n432_), .B(men_men_n154_), .C(men_men_n136_), .Y(men_men_n433_));
  NA2        u417(.A(men_men_n433_), .B(men_men_n431_), .Y(men_men_n434_));
  OAI210     u418(.A0(men_men_n434_), .A1(men_men_n426_), .B0(men_men_n34_), .Y(men_men_n435_));
  NO2        u419(.A(men_men_n411_), .B(men_men_n208_), .Y(men_men_n436_));
  NO4        u420(.A(men_men_n436_), .B(men_men_n77_), .C(x4), .D(men_men_n52_), .Y(men_men_n437_));
  NA2        u421(.A(men_men_n259_), .B(men_men_n21_), .Y(men_men_n438_));
  NO2        u422(.A(men_men_n163_), .B(men_men_n137_), .Y(men_men_n439_));
  NA2        u423(.A(men_men_n439_), .B(men_men_n438_), .Y(men_men_n440_));
  AOI210     u424(.A0(men_men_n440_), .A1(men_men_n170_), .B0(men_men_n27_), .Y(men_men_n441_));
  AOI220     u425(.A0(men_men_n365_), .A1(men_men_n91_), .B0(men_men_n152_), .B1(men_men_n202_), .Y(men_men_n442_));
  NA3        u426(.A(men_men_n442_), .B(men_men_n405_), .C(men_men_n89_), .Y(men_men_n443_));
  NA2        u427(.A(men_men_n443_), .B(men_men_n180_), .Y(men_men_n444_));
  OAI220     u428(.A0(x3), .A1(men_men_n67_), .B0(men_men_n163_), .B1(men_men_n41_), .Y(men_men_n445_));
  AOI210     u429(.A0(men_men_n167_), .A1(men_men_n26_), .B0(men_men_n72_), .Y(men_men_n446_));
  AOI220     u430(.A0(men_men_n446_), .A1(x0), .B0(men_men_n445_), .B1(men_men_n137_), .Y(men_men_n447_));
  AOI210     u431(.A0(men_men_n447_), .A1(men_men_n444_), .B0(men_men_n236_), .Y(men_men_n448_));
  NA2        u432(.A(x9), .B(x5), .Y(men_men_n449_));
  NO4        u433(.A(men_men_n106_), .B(men_men_n449_), .C(men_men_n58_), .D(men_men_n31_), .Y(men_men_n450_));
  NO4        u434(.A(men_men_n450_), .B(men_men_n448_), .C(men_men_n441_), .D(men_men_n437_), .Y(men_men_n451_));
  NA3        u435(.A(men_men_n451_), .B(men_men_n435_), .C(men_men_n397_), .Y(men_men_n452_));
  AOI210     u436(.A0(men_men_n380_), .A1(men_men_n24_), .B0(men_men_n452_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule