// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n139_,
    new_new_n140_, new_new_n141_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1092_, new_new_n1093_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  NO2        g0065(.A(i_2_), .B(i_7_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  OAI210     g0067(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n89_), .Y(new_new_n90_));
  NAi21      g0068(.An(i_6_), .B(i_10_), .Y(new_new_n91_));
  NA2        g0069(.A(i_6_), .B(i_9_), .Y(new_new_n92_));
  AOI210     g0070(.A0(new_new_n92_), .A1(new_new_n91_), .B0(new_new_n64_), .Y(new_new_n93_));
  NA2        g0071(.A(i_2_), .B(i_6_), .Y(new_new_n94_));
  NO3        g0072(.A(new_new_n94_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n95_));
  NO2        g0073(.A(new_new_n95_), .B(new_new_n93_), .Y(new_new_n96_));
  AOI210     g0074(.A0(new_new_n96_), .A1(new_new_n90_), .B0(new_new_n81_), .Y(new_new_n97_));
  AN3        g0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n98_));
  NAi21      g0076(.An(i_6_), .B(i_11_), .Y(new_new_n99_));
  NO2        g0077(.A(i_5_), .B(i_8_), .Y(new_new_n100_));
  NOi21      g0078(.An(new_new_n100_), .B(new_new_n99_), .Y(new_new_n101_));
  AOI220     g0079(.A0(new_new_n101_), .A1(new_new_n63_), .B0(new_new_n98_), .B1(new_new_n32_), .Y(new_new_n102_));
  INV        g0080(.A(i_7_), .Y(new_new_n103_));
  NA2        g0081(.A(new_new_n47_), .B(new_new_n103_), .Y(new_new_n104_));
  NO2        g0082(.A(i_0_), .B(i_5_), .Y(new_new_n105_));
  NO2        g0083(.A(new_new_n105_), .B(new_new_n87_), .Y(new_new_n106_));
  NA2        g0084(.A(i_12_), .B(i_3_), .Y(new_new_n107_));
  INV        g0085(.A(new_new_n107_), .Y(new_new_n108_));
  NA3        g0086(.A(new_new_n108_), .B(new_new_n106_), .C(new_new_n104_), .Y(new_new_n109_));
  NAi21      g0087(.An(i_7_), .B(i_11_), .Y(new_new_n110_));
  NO3        g0088(.A(new_new_n110_), .B(new_new_n91_), .C(new_new_n54_), .Y(new_new_n111_));
  AN2        g0089(.A(i_2_), .B(i_10_), .Y(new_new_n112_));
  NO2        g0090(.A(new_new_n112_), .B(i_7_), .Y(new_new_n113_));
  OR2        g0091(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n114_));
  NO2        g0092(.A(i_8_), .B(new_new_n103_), .Y(new_new_n115_));
  NO3        g0093(.A(new_new_n115_), .B(new_new_n114_), .C(new_new_n113_), .Y(new_new_n116_));
  NA2        g0094(.A(i_12_), .B(i_7_), .Y(new_new_n117_));
  NO2        g0095(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n118_));
  NA2        g0096(.A(i_11_), .B(i_12_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n1093_), .B(new_new_n116_), .Y(new_new_n120_));
  NAi41      g0098(.An(new_new_n111_), .B(new_new_n120_), .C(new_new_n109_), .D(new_new_n102_), .Y(new_new_n121_));
  NOi21      g0099(.An(i_1_), .B(i_5_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(i_11_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n124_));
  NA2        g0102(.A(i_7_), .B(new_new_n25_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n125_), .B(new_new_n124_), .Y(new_new_n126_));
  NO2        g0104(.A(new_new_n126_), .B(new_new_n47_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n92_), .B(new_new_n91_), .Y(new_new_n128_));
  NAi21      g0106(.An(i_3_), .B(i_8_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n129_), .B(new_new_n63_), .Y(new_new_n130_));
  NOi31      g0108(.An(new_new_n130_), .B(new_new_n128_), .C(new_new_n127_), .Y(new_new_n131_));
  NO2        g0109(.A(i_1_), .B(new_new_n87_), .Y(new_new_n132_));
  NO2        g0110(.A(i_6_), .B(i_5_), .Y(new_new_n133_));
  NA2        g0111(.A(new_new_n133_), .B(i_3_), .Y(new_new_n134_));
  AO210      g0112(.A0(new_new_n134_), .A1(new_new_n48_), .B0(new_new_n132_), .Y(new_new_n135_));
  OAI220     g0113(.A0(new_new_n135_), .A1(new_new_n110_), .B0(new_new_n131_), .B1(new_new_n123_), .Y(new_new_n136_));
  NO3        g0114(.A(new_new_n136_), .B(new_new_n121_), .C(new_new_n97_), .Y(new_new_n137_));
  NA3        g0115(.A(new_new_n137_), .B(new_new_n80_), .C(new_new_n57_), .Y(men2));
  NO2        g0116(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n139_));
  NA2        g0117(.A(i_6_), .B(new_new_n25_), .Y(new_new_n140_));
  NA2        g0118(.A(new_new_n140_), .B(new_new_n139_), .Y(new_new_n141_));
  NA4        g0119(.A(new_new_n141_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(men0));
  AN2        g0120(.A(i_8_), .B(i_7_), .Y(new_new_n143_));
  NA2        g0121(.A(new_new_n143_), .B(i_6_), .Y(new_new_n144_));
  NO2        g0122(.A(i_12_), .B(i_13_), .Y(new_new_n145_));
  NAi21      g0123(.An(i_5_), .B(i_11_), .Y(new_new_n146_));
  NOi21      g0124(.An(new_new_n145_), .B(new_new_n146_), .Y(new_new_n147_));
  NO2        g0125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NA2        g0126(.A(i_2_), .B(i_3_), .Y(new_new_n149_));
  NO2        g0127(.A(new_new_n149_), .B(i_4_), .Y(new_new_n150_));
  NA3        g0128(.A(new_new_n150_), .B(new_new_n148_), .C(new_new_n147_), .Y(new_new_n151_));
  AN2        g0129(.A(new_new_n145_), .B(new_new_n84_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n152_), .B(new_new_n27_), .Y(new_new_n153_));
  NA2        g0131(.A(i_1_), .B(i_5_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n155_));
  NA2        g0133(.A(new_new_n155_), .B(new_new_n36_), .Y(new_new_n156_));
  NO3        g0134(.A(new_new_n156_), .B(new_new_n154_), .C(new_new_n153_), .Y(new_new_n157_));
  OR2        g0135(.A(i_0_), .B(i_1_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n159_));
  NAi32      g0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n160_));
  NAi21      g0138(.An(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  NOi21      g0139(.An(i_4_), .B(i_10_), .Y(new_new_n162_));
  NA2        g0140(.A(new_new_n162_), .B(new_new_n40_), .Y(new_new_n163_));
  NO2        g0141(.A(i_3_), .B(i_5_), .Y(new_new_n164_));
  NO3        g0142(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n165_));
  NA2        g0143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OAI210     g0144(.A0(new_new_n166_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n167_));
  NO2        g0145(.A(new_new_n167_), .B(new_new_n157_), .Y(new_new_n168_));
  AOI210     g0146(.A0(new_new_n168_), .A1(new_new_n151_), .B0(new_new_n144_), .Y(new_new_n169_));
  NA3        g0147(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n170_));
  NA2        g0148(.A(i_3_), .B(new_new_n49_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_4_), .B(i_9_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_11_), .B(i_13_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n173_), .B(new_new_n172_), .Y(new_new_n174_));
  OR2        g0152(.A(new_new_n174_), .B(new_new_n171_), .Y(new_new_n175_));
  NO2        g0153(.A(i_4_), .B(i_5_), .Y(new_new_n176_));
  NAi21      g0154(.An(i_12_), .B(i_11_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n177_), .B(i_13_), .Y(new_new_n178_));
  NA3        g0156(.A(new_new_n178_), .B(new_new_n176_), .C(new_new_n84_), .Y(new_new_n179_));
  AOI210     g0157(.A0(new_new_n179_), .A1(new_new_n175_), .B0(new_new_n170_), .Y(new_new_n180_));
  NO2        g0158(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n181_), .B(new_new_n47_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n36_), .B(i_5_), .Y(new_new_n183_));
  NAi31      g0161(.An(new_new_n183_), .B(new_new_n152_), .C(i_11_), .Y(new_new_n184_));
  NA2        g0162(.A(i_3_), .B(i_5_), .Y(new_new_n185_));
  OR2        g0163(.A(new_new_n185_), .B(new_new_n174_), .Y(new_new_n186_));
  AOI210     g0164(.A0(new_new_n186_), .A1(new_new_n184_), .B0(new_new_n182_), .Y(new_new_n187_));
  NO2        g0165(.A(new_new_n74_), .B(i_5_), .Y(new_new_n188_));
  NO2        g0166(.A(i_13_), .B(i_10_), .Y(new_new_n189_));
  NA3        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n45_), .Y(new_new_n190_));
  NO2        g0168(.A(i_2_), .B(i_1_), .Y(new_new_n191_));
  NA2        g0169(.A(new_new_n191_), .B(i_3_), .Y(new_new_n192_));
  NAi21      g0170(.An(i_4_), .B(i_12_), .Y(new_new_n193_));
  NO4        g0171(.A(new_new_n193_), .B(new_new_n192_), .C(new_new_n190_), .D(new_new_n25_), .Y(new_new_n194_));
  NO3        g0172(.A(new_new_n194_), .B(new_new_n187_), .C(new_new_n180_), .Y(new_new_n195_));
  INV        g0173(.A(i_8_), .Y(new_new_n196_));
  NO2        g0174(.A(new_new_n196_), .B(i_7_), .Y(new_new_n197_));
  NA2        g0175(.A(new_new_n197_), .B(i_6_), .Y(new_new_n198_));
  NO3        g0176(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n199_));
  NA2        g0177(.A(new_new_n199_), .B(new_new_n115_), .Y(new_new_n200_));
  NO3        g0178(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n201_));
  NA3        g0179(.A(new_new_n201_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n202_));
  NO3        g0180(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n203_));
  OAI210     g0181(.A0(new_new_n98_), .A1(i_12_), .B0(new_new_n203_), .Y(new_new_n204_));
  AOI210     g0182(.A0(new_new_n204_), .A1(new_new_n202_), .B0(new_new_n200_), .Y(new_new_n205_));
  NO2        g0183(.A(i_3_), .B(i_8_), .Y(new_new_n206_));
  NO3        g0184(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n207_));
  NO2        g0185(.A(new_new_n105_), .B(new_new_n59_), .Y(new_new_n208_));
  NO2        g0186(.A(i_13_), .B(i_9_), .Y(new_new_n209_));
  NA3        g0187(.A(new_new_n209_), .B(i_6_), .C(new_new_n196_), .Y(new_new_n210_));
  NAi21      g0188(.An(i_12_), .B(i_3_), .Y(new_new_n211_));
  NO2        g0189(.A(new_new_n45_), .B(i_5_), .Y(new_new_n212_));
  NO3        g0190(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n213_));
  NA3        g0191(.A(new_new_n213_), .B(new_new_n212_), .C(i_10_), .Y(new_new_n214_));
  NO2        g0192(.A(new_new_n214_), .B(new_new_n210_), .Y(new_new_n215_));
  AOI210     g0193(.A0(new_new_n215_), .A1(i_7_), .B0(new_new_n205_), .Y(new_new_n216_));
  OAI220     g0194(.A0(new_new_n216_), .A1(i_4_), .B0(new_new_n198_), .B1(new_new_n195_), .Y(new_new_n217_));
  NAi21      g0195(.An(i_12_), .B(i_7_), .Y(new_new_n218_));
  NA3        g0196(.A(i_13_), .B(new_new_n196_), .C(i_10_), .Y(new_new_n219_));
  NO2        g0197(.A(new_new_n219_), .B(new_new_n218_), .Y(new_new_n220_));
  NA2        g0198(.A(i_0_), .B(i_5_), .Y(new_new_n221_));
  NA2        g0199(.A(new_new_n221_), .B(new_new_n106_), .Y(new_new_n222_));
  OAI220     g0200(.A0(new_new_n222_), .A1(new_new_n192_), .B0(new_new_n182_), .B1(new_new_n134_), .Y(new_new_n223_));
  NAi31      g0201(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n36_), .B(i_13_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n226_));
  NO2        g0204(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n227_));
  NA3        g0205(.A(new_new_n227_), .B(new_new_n226_), .C(new_new_n225_), .Y(new_new_n228_));
  INV        g0206(.A(i_13_), .Y(new_new_n229_));
  NO2        g0207(.A(i_12_), .B(new_new_n229_), .Y(new_new_n230_));
  NA3        g0208(.A(new_new_n230_), .B(new_new_n201_), .C(new_new_n199_), .Y(new_new_n231_));
  OAI210     g0209(.A0(new_new_n228_), .A1(new_new_n224_), .B0(new_new_n231_), .Y(new_new_n232_));
  AOI220     g0210(.A0(new_new_n232_), .A1(new_new_n143_), .B0(new_new_n223_), .B1(new_new_n220_), .Y(new_new_n233_));
  NO2        g0211(.A(i_12_), .B(new_new_n37_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n185_), .B(i_4_), .Y(new_new_n235_));
  NA2        g0213(.A(new_new_n235_), .B(new_new_n234_), .Y(new_new_n236_));
  OR2        g0214(.A(i_8_), .B(i_7_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n237_), .B(new_new_n87_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n54_), .B(i_1_), .Y(new_new_n239_));
  NA2        g0217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  INV        g0218(.A(i_12_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n45_), .B(new_new_n241_), .Y(new_new_n242_));
  NO3        g0220(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n243_));
  NA2        g0221(.A(i_2_), .B(i_1_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n240_), .B(new_new_n236_), .Y(new_new_n245_));
  NO3        g0223(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n246_));
  NAi21      g0224(.An(i_4_), .B(i_3_), .Y(new_new_n247_));
  NO2        g0225(.A(new_new_n247_), .B(new_new_n76_), .Y(new_new_n248_));
  NO2        g0226(.A(i_0_), .B(i_6_), .Y(new_new_n249_));
  NOi41      g0227(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n250_));
  NA2        g0228(.A(new_new_n250_), .B(new_new_n249_), .Y(new_new_n251_));
  NO2        g0229(.A(new_new_n244_), .B(new_new_n185_), .Y(new_new_n252_));
  NAi21      g0230(.An(new_new_n251_), .B(new_new_n252_), .Y(new_new_n253_));
  INV        g0231(.A(new_new_n253_), .Y(new_new_n254_));
  AOI220     g0232(.A0(new_new_n254_), .A1(new_new_n40_), .B0(new_new_n245_), .B1(new_new_n209_), .Y(new_new_n255_));
  NO2        g0233(.A(i_11_), .B(new_new_n229_), .Y(new_new_n256_));
  NOi21      g0234(.An(i_1_), .B(i_6_), .Y(new_new_n257_));
  NAi21      g0235(.An(i_3_), .B(i_7_), .Y(new_new_n258_));
  NA2        g0236(.A(new_new_n241_), .B(i_9_), .Y(new_new_n259_));
  OR4        g0237(.A(new_new_n259_), .B(new_new_n258_), .C(new_new_n257_), .D(new_new_n188_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n261_));
  NO2        g0239(.A(i_12_), .B(i_3_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n74_), .B(i_5_), .Y(new_new_n263_));
  NA2        g0241(.A(i_3_), .B(i_9_), .Y(new_new_n264_));
  NAi21      g0242(.An(i_7_), .B(i_10_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n266_));
  NA3        g0244(.A(new_new_n266_), .B(new_new_n263_), .C(new_new_n65_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n267_), .B(new_new_n260_), .Y(new_new_n268_));
  NA3        g0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n269_));
  INV        g0247(.A(new_new_n144_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n241_), .B(i_13_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n271_), .B(new_new_n76_), .Y(new_new_n272_));
  AOI220     g0250(.A0(new_new_n272_), .A1(new_new_n270_), .B0(new_new_n268_), .B1(new_new_n256_), .Y(new_new_n273_));
  NO2        g0251(.A(new_new_n237_), .B(new_new_n37_), .Y(new_new_n274_));
  NA2        g0252(.A(i_12_), .B(i_6_), .Y(new_new_n275_));
  OR2        g0253(.A(i_13_), .B(i_9_), .Y(new_new_n276_));
  NO3        g0254(.A(new_new_n276_), .B(new_new_n275_), .C(new_new_n49_), .Y(new_new_n277_));
  NO2        g0255(.A(new_new_n247_), .B(i_2_), .Y(new_new_n278_));
  NA2        g0256(.A(new_new_n256_), .B(i_9_), .Y(new_new_n279_));
  NA2        g0257(.A(new_new_n155_), .B(new_new_n64_), .Y(new_new_n280_));
  NO3        g0258(.A(i_11_), .B(new_new_n229_), .C(new_new_n25_), .Y(new_new_n281_));
  NO2        g0259(.A(new_new_n258_), .B(i_8_), .Y(new_new_n282_));
  NO2        g0260(.A(i_6_), .B(new_new_n49_), .Y(new_new_n283_));
  NA3        g0261(.A(new_new_n283_), .B(new_new_n282_), .C(new_new_n281_), .Y(new_new_n284_));
  NO3        g0262(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n285_));
  NA3        g0263(.A(new_new_n285_), .B(new_new_n274_), .C(new_new_n230_), .Y(new_new_n286_));
  AOI210     g0264(.A0(new_new_n286_), .A1(new_new_n284_), .B0(new_new_n280_), .Y(new_new_n287_));
  INV        g0265(.A(new_new_n287_), .Y(new_new_n288_));
  NA4        g0266(.A(new_new_n288_), .B(new_new_n273_), .C(new_new_n255_), .D(new_new_n233_), .Y(new_new_n289_));
  NO3        g0267(.A(i_12_), .B(new_new_n229_), .C(new_new_n37_), .Y(new_new_n290_));
  INV        g0268(.A(new_new_n290_), .Y(new_new_n291_));
  NA2        g0269(.A(i_8_), .B(new_new_n103_), .Y(new_new_n292_));
  NOi21      g0270(.An(new_new_n164_), .B(new_new_n87_), .Y(new_new_n293_));
  NO3        g0271(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n294_));
  AOI220     g0272(.A0(new_new_n294_), .A1(new_new_n199_), .B0(new_new_n293_), .B1(new_new_n239_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n295_), .B(new_new_n292_), .Y(new_new_n296_));
  NO3        g0274(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n244_), .B(i_0_), .Y(new_new_n298_));
  AOI220     g0276(.A0(new_new_n298_), .A1(new_new_n197_), .B0(new_new_n297_), .B1(new_new_n143_), .Y(new_new_n299_));
  NA2        g0277(.A(new_new_n283_), .B(new_new_n26_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n300_), .B(new_new_n299_), .Y(new_new_n301_));
  NA2        g0279(.A(i_0_), .B(i_1_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n302_), .B(i_2_), .Y(new_new_n303_));
  NO2        g0281(.A(new_new_n60_), .B(i_6_), .Y(new_new_n304_));
  NA3        g0282(.A(new_new_n304_), .B(new_new_n303_), .C(new_new_n164_), .Y(new_new_n305_));
  OAI210     g0283(.A0(new_new_n166_), .A1(new_new_n144_), .B0(new_new_n305_), .Y(new_new_n306_));
  NO3        g0284(.A(new_new_n306_), .B(new_new_n301_), .C(new_new_n296_), .Y(new_new_n307_));
  NO2        g0285(.A(i_3_), .B(i_10_), .Y(new_new_n308_));
  NA3        g0286(.A(new_new_n308_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n309_));
  NO2        g0287(.A(i_2_), .B(new_new_n103_), .Y(new_new_n310_));
  NA2        g0288(.A(i_1_), .B(new_new_n36_), .Y(new_new_n311_));
  NO2        g0289(.A(new_new_n311_), .B(i_8_), .Y(new_new_n312_));
  NA2        g0290(.A(new_new_n312_), .B(new_new_n310_), .Y(new_new_n313_));
  AN2        g0291(.A(i_3_), .B(i_10_), .Y(new_new_n314_));
  NA4        g0292(.A(new_new_n314_), .B(new_new_n201_), .C(new_new_n178_), .D(new_new_n176_), .Y(new_new_n315_));
  NO2        g0293(.A(i_5_), .B(new_new_n37_), .Y(new_new_n316_));
  NO2        g0294(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n317_));
  OR2        g0295(.A(new_new_n313_), .B(new_new_n309_), .Y(new_new_n318_));
  OAI220     g0296(.A0(new_new_n318_), .A1(i_6_), .B0(new_new_n307_), .B1(new_new_n291_), .Y(new_new_n319_));
  NO4        g0297(.A(new_new_n319_), .B(new_new_n289_), .C(new_new_n217_), .D(new_new_n169_), .Y(new_new_n320_));
  NO3        g0298(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n321_));
  NO2        g0299(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n322_));
  NA2        g0300(.A(new_new_n298_), .B(new_new_n322_), .Y(new_new_n323_));
  NO3        g0301(.A(i_6_), .B(new_new_n196_), .C(i_7_), .Y(new_new_n324_));
  NA2        g0302(.A(new_new_n324_), .B(new_new_n201_), .Y(new_new_n325_));
  AOI210     g0303(.A0(new_new_n325_), .A1(new_new_n323_), .B0(new_new_n171_), .Y(new_new_n326_));
  NO2        g0304(.A(i_2_), .B(i_3_), .Y(new_new_n327_));
  OR2        g0305(.A(i_0_), .B(i_5_), .Y(new_new_n328_));
  NA2        g0306(.A(new_new_n221_), .B(new_new_n328_), .Y(new_new_n329_));
  NA4        g0307(.A(new_new_n329_), .B(new_new_n238_), .C(new_new_n327_), .D(i_1_), .Y(new_new_n330_));
  NA3        g0308(.A(new_new_n298_), .B(new_new_n293_), .C(new_new_n115_), .Y(new_new_n331_));
  NAi21      g0309(.An(i_8_), .B(i_7_), .Y(new_new_n332_));
  NO2        g0310(.A(new_new_n332_), .B(i_6_), .Y(new_new_n333_));
  NO2        g0311(.A(new_new_n158_), .B(new_new_n47_), .Y(new_new_n334_));
  NA3        g0312(.A(new_new_n334_), .B(new_new_n333_), .C(new_new_n164_), .Y(new_new_n335_));
  NA3        g0313(.A(new_new_n335_), .B(new_new_n331_), .C(new_new_n330_), .Y(new_new_n336_));
  OAI210     g0314(.A0(new_new_n336_), .A1(new_new_n326_), .B0(i_4_), .Y(new_new_n337_));
  NO2        g0315(.A(i_12_), .B(i_10_), .Y(new_new_n338_));
  NOi21      g0316(.An(i_5_), .B(i_0_), .Y(new_new_n339_));
  NO3        g0317(.A(new_new_n311_), .B(new_new_n339_), .C(new_new_n129_), .Y(new_new_n340_));
  NA4        g0318(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n341_));
  NA2        g0319(.A(new_new_n340_), .B(new_new_n338_), .Y(new_new_n342_));
  NO2        g0320(.A(i_6_), .B(i_8_), .Y(new_new_n343_));
  NOi21      g0321(.An(i_0_), .B(i_2_), .Y(new_new_n344_));
  AN2        g0322(.A(new_new_n344_), .B(new_new_n343_), .Y(new_new_n345_));
  NO2        g0323(.A(i_1_), .B(i_7_), .Y(new_new_n346_));
  AO220      g0324(.A0(new_new_n346_), .A1(new_new_n345_), .B0(new_new_n333_), .B1(new_new_n239_), .Y(new_new_n347_));
  NA3        g0325(.A(new_new_n347_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n348_));
  NA3        g0326(.A(new_new_n348_), .B(new_new_n342_), .C(new_new_n337_), .Y(new_new_n349_));
  NO3        g0327(.A(new_new_n237_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n350_));
  NO3        g0328(.A(new_new_n332_), .B(i_2_), .C(i_1_), .Y(new_new_n351_));
  OAI210     g0329(.A0(new_new_n351_), .A1(new_new_n350_), .B0(i_6_), .Y(new_new_n352_));
  NA3        g0330(.A(new_new_n257_), .B(new_new_n310_), .C(new_new_n196_), .Y(new_new_n353_));
  AOI210     g0331(.A0(new_new_n353_), .A1(new_new_n352_), .B0(new_new_n329_), .Y(new_new_n354_));
  NOi21      g0332(.An(new_new_n154_), .B(new_new_n106_), .Y(new_new_n355_));
  NO2        g0333(.A(new_new_n355_), .B(new_new_n125_), .Y(new_new_n356_));
  OAI210     g0334(.A0(new_new_n356_), .A1(new_new_n354_), .B0(i_3_), .Y(new_new_n357_));
  INV        g0335(.A(new_new_n85_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n302_), .B(new_new_n82_), .Y(new_new_n359_));
  NA2        g0337(.A(new_new_n359_), .B(new_new_n133_), .Y(new_new_n360_));
  NO2        g0338(.A(new_new_n94_), .B(new_new_n196_), .Y(new_new_n361_));
  NA2        g0339(.A(new_new_n361_), .B(new_new_n64_), .Y(new_new_n362_));
  AOI210     g0340(.A0(new_new_n362_), .A1(new_new_n360_), .B0(new_new_n358_), .Y(new_new_n363_));
  NO2        g0341(.A(new_new_n196_), .B(i_9_), .Y(new_new_n364_));
  NA2        g0342(.A(new_new_n364_), .B(new_new_n208_), .Y(new_new_n365_));
  NO2        g0343(.A(new_new_n365_), .B(new_new_n47_), .Y(new_new_n366_));
  NO3        g0344(.A(new_new_n366_), .B(new_new_n363_), .C(new_new_n301_), .Y(new_new_n367_));
  AOI210     g0345(.A0(new_new_n367_), .A1(new_new_n357_), .B0(new_new_n163_), .Y(new_new_n368_));
  AOI210     g0346(.A0(new_new_n349_), .A1(new_new_n321_), .B0(new_new_n368_), .Y(new_new_n369_));
  NOi32      g0347(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n370_));
  INV        g0348(.A(new_new_n370_), .Y(new_new_n371_));
  NAi21      g0349(.An(i_0_), .B(i_6_), .Y(new_new_n372_));
  NAi21      g0350(.An(i_1_), .B(i_5_), .Y(new_new_n373_));
  NA2        g0351(.A(new_new_n373_), .B(new_new_n372_), .Y(new_new_n374_));
  NA2        g0352(.A(new_new_n374_), .B(new_new_n25_), .Y(new_new_n375_));
  OAI210     g0353(.A0(new_new_n375_), .A1(new_new_n160_), .B0(new_new_n251_), .Y(new_new_n376_));
  NAi41      g0354(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n377_));
  AOI210     g0355(.A0(new_new_n377_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n378_));
  NOi32      g0356(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n379_));
  NAi21      g0357(.An(i_6_), .B(i_1_), .Y(new_new_n380_));
  NA3        g0358(.A(new_new_n380_), .B(new_new_n379_), .C(new_new_n47_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n381_), .B(i_0_), .Y(new_new_n382_));
  OR2        g0360(.A(new_new_n382_), .B(new_new_n378_), .Y(new_new_n383_));
  NO2        g0361(.A(i_1_), .B(new_new_n103_), .Y(new_new_n384_));
  NAi21      g0362(.An(i_3_), .B(i_4_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n385_), .B(i_9_), .Y(new_new_n386_));
  AN2        g0364(.A(i_6_), .B(i_7_), .Y(new_new_n387_));
  OAI210     g0365(.A0(new_new_n387_), .A1(new_new_n384_), .B0(new_new_n386_), .Y(new_new_n388_));
  NA2        g0366(.A(i_2_), .B(i_7_), .Y(new_new_n389_));
  NO2        g0367(.A(new_new_n385_), .B(i_10_), .Y(new_new_n390_));
  NA3        g0368(.A(new_new_n390_), .B(new_new_n389_), .C(new_new_n249_), .Y(new_new_n391_));
  AOI210     g0369(.A0(new_new_n391_), .A1(new_new_n388_), .B0(new_new_n188_), .Y(new_new_n392_));
  AOI210     g0370(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n393_));
  OAI210     g0371(.A0(new_new_n393_), .A1(new_new_n191_), .B0(new_new_n390_), .Y(new_new_n394_));
  AOI220     g0372(.A0(new_new_n390_), .A1(new_new_n346_), .B0(new_new_n243_), .B1(new_new_n191_), .Y(new_new_n395_));
  AOI210     g0373(.A0(new_new_n395_), .A1(new_new_n394_), .B0(i_5_), .Y(new_new_n396_));
  NO4        g0374(.A(new_new_n396_), .B(new_new_n392_), .C(new_new_n383_), .D(new_new_n376_), .Y(new_new_n397_));
  NO2        g0375(.A(new_new_n397_), .B(new_new_n371_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n399_));
  AN2        g0377(.A(i_12_), .B(i_5_), .Y(new_new_n400_));
  NO2        g0378(.A(i_4_), .B(new_new_n26_), .Y(new_new_n401_));
  NA2        g0379(.A(new_new_n401_), .B(new_new_n400_), .Y(new_new_n402_));
  NO2        g0380(.A(i_11_), .B(i_6_), .Y(new_new_n403_));
  NA3        g0381(.A(new_new_n403_), .B(new_new_n334_), .C(new_new_n229_), .Y(new_new_n404_));
  NO2        g0382(.A(new_new_n404_), .B(new_new_n402_), .Y(new_new_n405_));
  NO2        g0383(.A(new_new_n247_), .B(i_5_), .Y(new_new_n406_));
  NO2        g0384(.A(i_5_), .B(i_10_), .Y(new_new_n407_));
  AOI220     g0385(.A0(new_new_n407_), .A1(new_new_n278_), .B0(new_new_n406_), .B1(new_new_n201_), .Y(new_new_n408_));
  NA2        g0386(.A(new_new_n145_), .B(new_new_n46_), .Y(new_new_n409_));
  NO2        g0387(.A(new_new_n409_), .B(new_new_n408_), .Y(new_new_n410_));
  OAI210     g0388(.A0(new_new_n410_), .A1(new_new_n405_), .B0(new_new_n399_), .Y(new_new_n411_));
  NO2        g0389(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n151_), .B(new_new_n87_), .Y(new_new_n413_));
  OAI210     g0391(.A0(new_new_n413_), .A1(new_new_n405_), .B0(new_new_n412_), .Y(new_new_n414_));
  NO3        g0392(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n415_));
  NO2        g0393(.A(i_3_), .B(new_new_n103_), .Y(new_new_n416_));
  NO2        g0394(.A(i_11_), .B(i_12_), .Y(new_new_n417_));
  NA2        g0395(.A(new_new_n407_), .B(new_new_n241_), .Y(new_new_n418_));
  NA3        g0396(.A(new_new_n115_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n419_));
  OAI220     g0397(.A0(new_new_n419_), .A1(new_new_n224_), .B0(new_new_n418_), .B1(new_new_n341_), .Y(new_new_n420_));
  NAi21      g0398(.An(i_13_), .B(i_0_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n421_), .B(new_new_n244_), .Y(new_new_n422_));
  NA2        g0400(.A(new_new_n420_), .B(new_new_n422_), .Y(new_new_n423_));
  NA3        g0401(.A(new_new_n423_), .B(new_new_n414_), .C(new_new_n411_), .Y(new_new_n424_));
  NO3        g0402(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n425_));
  NO2        g0403(.A(i_0_), .B(i_11_), .Y(new_new_n426_));
  INV        g0404(.A(i_5_), .Y(new_new_n427_));
  AN2        g0405(.A(i_1_), .B(i_6_), .Y(new_new_n428_));
  NOi21      g0406(.An(i_2_), .B(i_12_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n429_), .B(new_new_n428_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n430_), .B(new_new_n427_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n143_), .B(i_9_), .Y(new_new_n432_));
  NO2        g0410(.A(new_new_n432_), .B(i_4_), .Y(new_new_n433_));
  NA2        g0411(.A(new_new_n431_), .B(new_new_n433_), .Y(new_new_n434_));
  NAi21      g0412(.An(i_9_), .B(i_4_), .Y(new_new_n435_));
  OR2        g0413(.A(i_13_), .B(i_10_), .Y(new_new_n436_));
  NO3        g0414(.A(new_new_n436_), .B(new_new_n119_), .C(new_new_n435_), .Y(new_new_n437_));
  NO2        g0415(.A(new_new_n174_), .B(new_new_n124_), .Y(new_new_n438_));
  OR2        g0416(.A(new_new_n219_), .B(new_new_n218_), .Y(new_new_n439_));
  NO2        g0417(.A(new_new_n103_), .B(new_new_n25_), .Y(new_new_n440_));
  NA2        g0418(.A(new_new_n290_), .B(new_new_n440_), .Y(new_new_n441_));
  NA2        g0419(.A(new_new_n283_), .B(new_new_n213_), .Y(new_new_n442_));
  OAI220     g0420(.A0(new_new_n442_), .A1(new_new_n439_), .B0(new_new_n441_), .B1(new_new_n355_), .Y(new_new_n443_));
  INV        g0421(.A(new_new_n443_), .Y(new_new_n444_));
  AOI210     g0422(.A0(new_new_n444_), .A1(new_new_n434_), .B0(new_new_n26_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n331_), .B(new_new_n330_), .Y(new_new_n446_));
  AOI220     g0424(.A0(new_new_n304_), .A1(new_new_n294_), .B0(new_new_n298_), .B1(new_new_n322_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n447_), .B(new_new_n171_), .Y(new_new_n448_));
  NO2        g0426(.A(new_new_n185_), .B(new_new_n87_), .Y(new_new_n449_));
  AOI220     g0427(.A0(new_new_n449_), .A1(new_new_n303_), .B0(new_new_n285_), .B1(new_new_n213_), .Y(new_new_n450_));
  NO2        g0428(.A(new_new_n450_), .B(new_new_n292_), .Y(new_new_n451_));
  NO3        g0429(.A(new_new_n451_), .B(new_new_n448_), .C(new_new_n446_), .Y(new_new_n452_));
  NA2        g0430(.A(new_new_n199_), .B(new_new_n98_), .Y(new_new_n453_));
  NA3        g0431(.A(new_new_n334_), .B(new_new_n164_), .C(new_new_n87_), .Y(new_new_n454_));
  AOI210     g0432(.A0(new_new_n454_), .A1(new_new_n453_), .B0(new_new_n332_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n196_), .B(i_10_), .Y(new_new_n456_));
  NA3        g0434(.A(new_new_n263_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n304_), .B(new_new_n239_), .Y(new_new_n458_));
  OAI220     g0436(.A0(new_new_n458_), .A1(new_new_n185_), .B0(new_new_n457_), .B1(new_new_n456_), .Y(new_new_n459_));
  NO2        g0437(.A(i_3_), .B(new_new_n49_), .Y(new_new_n460_));
  NA3        g0438(.A(new_new_n346_), .B(new_new_n345_), .C(new_new_n460_), .Y(new_new_n461_));
  NA2        g0439(.A(new_new_n324_), .B(new_new_n329_), .Y(new_new_n462_));
  OAI210     g0440(.A0(new_new_n462_), .A1(new_new_n192_), .B0(new_new_n461_), .Y(new_new_n463_));
  NO3        g0441(.A(new_new_n463_), .B(new_new_n459_), .C(new_new_n455_), .Y(new_new_n464_));
  AOI210     g0442(.A0(new_new_n464_), .A1(new_new_n452_), .B0(new_new_n279_), .Y(new_new_n465_));
  NO4        g0443(.A(new_new_n465_), .B(new_new_n445_), .C(new_new_n424_), .D(new_new_n398_), .Y(new_new_n466_));
  NO2        g0444(.A(new_new_n64_), .B(i_4_), .Y(new_new_n467_));
  NO2        g0445(.A(new_new_n74_), .B(i_13_), .Y(new_new_n468_));
  NO2        g0446(.A(i_10_), .B(i_9_), .Y(new_new_n469_));
  NAi21      g0447(.An(i_12_), .B(i_8_), .Y(new_new_n470_));
  NO2        g0448(.A(new_new_n470_), .B(i_3_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n47_), .B(i_4_), .Y(new_new_n472_));
  NA2        g0450(.A(new_new_n317_), .B(i_0_), .Y(new_new_n473_));
  NO3        g0451(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n275_), .B(new_new_n99_), .Y(new_new_n475_));
  NA2        g0453(.A(new_new_n475_), .B(new_new_n474_), .Y(new_new_n476_));
  NA2        g0454(.A(i_8_), .B(i_9_), .Y(new_new_n477_));
  AOI210     g0455(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n478_));
  OR2        g0456(.A(new_new_n478_), .B(new_new_n477_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n290_), .B(new_new_n208_), .Y(new_new_n480_));
  NO2        g0458(.A(new_new_n480_), .B(new_new_n479_), .Y(new_new_n481_));
  NA2        g0459(.A(new_new_n256_), .B(new_new_n316_), .Y(new_new_n482_));
  NO3        g0460(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n483_));
  INV        g0461(.A(new_new_n483_), .Y(new_new_n484_));
  NA3        g0462(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n485_));
  NA4        g0463(.A(new_new_n146_), .B(new_new_n118_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n486_));
  OAI220     g0464(.A0(new_new_n486_), .A1(new_new_n485_), .B0(new_new_n484_), .B1(new_new_n482_), .Y(new_new_n487_));
  NO2        g0465(.A(new_new_n487_), .B(new_new_n481_), .Y(new_new_n488_));
  INV        g0466(.A(new_new_n303_), .Y(new_new_n489_));
  OR2        g0467(.A(new_new_n489_), .B(new_new_n210_), .Y(new_new_n490_));
  OA210      g0468(.A0(new_new_n365_), .A1(new_new_n103_), .B0(new_new_n305_), .Y(new_new_n491_));
  OA220      g0469(.A0(new_new_n491_), .A1(new_new_n163_), .B0(new_new_n490_), .B1(new_new_n236_), .Y(new_new_n492_));
  NA2        g0470(.A(new_new_n98_), .B(i_13_), .Y(new_new_n493_));
  NA2        g0471(.A(new_new_n449_), .B(new_new_n399_), .Y(new_new_n494_));
  NO2        g0472(.A(i_2_), .B(i_13_), .Y(new_new_n495_));
  NO2        g0473(.A(new_new_n494_), .B(new_new_n493_), .Y(new_new_n496_));
  NO3        g0474(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n497_));
  NO2        g0475(.A(i_6_), .B(i_7_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n498_), .B(new_new_n497_), .Y(new_new_n499_));
  NO2        g0477(.A(i_11_), .B(i_1_), .Y(new_new_n500_));
  NO2        g0478(.A(new_new_n74_), .B(i_3_), .Y(new_new_n501_));
  OR2        g0479(.A(i_11_), .B(i_8_), .Y(new_new_n502_));
  NOi21      g0480(.An(i_2_), .B(i_7_), .Y(new_new_n503_));
  NAi31      g0481(.An(new_new_n502_), .B(new_new_n503_), .C(new_new_n501_), .Y(new_new_n504_));
  NO2        g0482(.A(new_new_n436_), .B(i_6_), .Y(new_new_n505_));
  NA2        g0483(.A(new_new_n505_), .B(new_new_n467_), .Y(new_new_n506_));
  NO2        g0484(.A(new_new_n506_), .B(new_new_n504_), .Y(new_new_n507_));
  NO2        g0485(.A(i_3_), .B(new_new_n196_), .Y(new_new_n508_));
  NO2        g0486(.A(i_6_), .B(i_10_), .Y(new_new_n509_));
  NA4        g0487(.A(new_new_n509_), .B(new_new_n321_), .C(new_new_n508_), .D(new_new_n241_), .Y(new_new_n510_));
  NO2        g0488(.A(new_new_n510_), .B(new_new_n156_), .Y(new_new_n511_));
  NA3        g0489(.A(new_new_n250_), .B(new_new_n173_), .C(new_new_n133_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n513_));
  NO2        g0491(.A(new_new_n158_), .B(i_3_), .Y(new_new_n514_));
  NAi31      g0492(.An(new_new_n513_), .B(new_new_n514_), .C(new_new_n230_), .Y(new_new_n515_));
  NA3        g0493(.A(new_new_n412_), .B(new_new_n181_), .C(new_new_n150_), .Y(new_new_n516_));
  NA3        g0494(.A(new_new_n516_), .B(new_new_n515_), .C(new_new_n512_), .Y(new_new_n517_));
  NO4        g0495(.A(new_new_n517_), .B(new_new_n511_), .C(new_new_n507_), .D(new_new_n496_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n474_), .B(new_new_n400_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n483_), .B(new_new_n407_), .Y(new_new_n520_));
  NO2        g0498(.A(new_new_n520_), .B(new_new_n228_), .Y(new_new_n521_));
  NAi21      g0499(.An(new_new_n219_), .B(new_new_n417_), .Y(new_new_n522_));
  NO2        g0500(.A(new_new_n26_), .B(i_5_), .Y(new_new_n523_));
  NO2        g0501(.A(i_0_), .B(new_new_n87_), .Y(new_new_n524_));
  NA3        g0502(.A(new_new_n524_), .B(new_new_n523_), .C(new_new_n143_), .Y(new_new_n525_));
  OR3        g0503(.A(new_new_n311_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n526_));
  NO2        g0504(.A(new_new_n526_), .B(new_new_n525_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n27_), .B(i_10_), .Y(new_new_n528_));
  NA2        g0506(.A(new_new_n321_), .B(new_new_n243_), .Y(new_new_n529_));
  OAI220     g0507(.A0(new_new_n529_), .A1(new_new_n457_), .B0(new_new_n528_), .B1(new_new_n493_), .Y(new_new_n530_));
  NA4        g0508(.A(new_new_n314_), .B(new_new_n227_), .C(new_new_n74_), .D(new_new_n241_), .Y(new_new_n531_));
  NO2        g0509(.A(new_new_n531_), .B(new_new_n499_), .Y(new_new_n532_));
  NO4        g0510(.A(new_new_n532_), .B(new_new_n530_), .C(new_new_n527_), .D(new_new_n521_), .Y(new_new_n533_));
  NA4        g0511(.A(new_new_n533_), .B(new_new_n518_), .C(new_new_n492_), .D(new_new_n488_), .Y(new_new_n534_));
  NA3        g0512(.A(new_new_n314_), .B(new_new_n178_), .C(new_new_n176_), .Y(new_new_n535_));
  OAI210     g0513(.A0(new_new_n309_), .A1(new_new_n183_), .B0(new_new_n535_), .Y(new_new_n536_));
  AN2        g0514(.A(new_new_n294_), .B(new_new_n238_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n537_), .B(new_new_n536_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n321_), .B(new_new_n165_), .Y(new_new_n539_));
  OAI210     g0517(.A0(new_new_n539_), .A1(new_new_n236_), .B0(new_new_n315_), .Y(new_new_n540_));
  NA2        g0518(.A(new_new_n540_), .B(new_new_n333_), .Y(new_new_n541_));
  NA2        g0519(.A(new_new_n400_), .B(new_new_n229_), .Y(new_new_n542_));
  NA2        g0520(.A(new_new_n370_), .B(new_new_n74_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n387_), .B(new_new_n379_), .Y(new_new_n544_));
  AO210      g0522(.A0(new_new_n543_), .A1(new_new_n542_), .B0(new_new_n544_), .Y(new_new_n545_));
  NO2        g0523(.A(new_new_n36_), .B(i_8_), .Y(new_new_n546_));
  NAi41      g0524(.An(new_new_n543_), .B(new_new_n509_), .C(new_new_n546_), .D(new_new_n47_), .Y(new_new_n547_));
  AOI210     g0525(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n437_), .Y(new_new_n548_));
  NA3        g0526(.A(new_new_n548_), .B(new_new_n547_), .C(new_new_n545_), .Y(new_new_n549_));
  INV        g0527(.A(new_new_n549_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n263_), .B(new_new_n65_), .Y(new_new_n551_));
  OAI210     g0529(.A0(i_8_), .A1(new_new_n551_), .B0(new_new_n135_), .Y(new_new_n552_));
  AOI210     g0530(.A0(new_new_n197_), .A1(i_9_), .B0(new_new_n274_), .Y(new_new_n553_));
  NO2        g0531(.A(new_new_n553_), .B(new_new_n202_), .Y(new_new_n554_));
  OR2        g0532(.A(new_new_n185_), .B(i_4_), .Y(new_new_n555_));
  NO2        g0533(.A(new_new_n555_), .B(new_new_n87_), .Y(new_new_n556_));
  AOI220     g0534(.A0(new_new_n556_), .A1(new_new_n554_), .B0(new_new_n552_), .B1(new_new_n438_), .Y(new_new_n557_));
  NA4        g0535(.A(new_new_n557_), .B(new_new_n550_), .C(new_new_n541_), .D(new_new_n538_), .Y(new_new_n558_));
  NA2        g0536(.A(new_new_n406_), .B(new_new_n303_), .Y(new_new_n559_));
  OAI210     g0537(.A0(new_new_n402_), .A1(new_new_n170_), .B0(new_new_n559_), .Y(new_new_n560_));
  NO2        g0538(.A(i_12_), .B(new_new_n196_), .Y(new_new_n561_));
  NA2        g0539(.A(new_new_n561_), .B(new_new_n229_), .Y(new_new_n562_));
  NA3        g0540(.A(new_new_n509_), .B(new_new_n176_), .C(new_new_n27_), .Y(new_new_n563_));
  NO2        g0541(.A(new_new_n563_), .B(new_new_n562_), .Y(new_new_n564_));
  NOi31      g0542(.An(new_new_n324_), .B(new_new_n436_), .C(new_new_n38_), .Y(new_new_n565_));
  OAI210     g0543(.A0(new_new_n565_), .A1(new_new_n564_), .B0(new_new_n560_), .Y(new_new_n566_));
  NO2        g0544(.A(i_8_), .B(i_7_), .Y(new_new_n567_));
  OAI210     g0545(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n568_));
  NA2        g0546(.A(new_new_n568_), .B(new_new_n227_), .Y(new_new_n569_));
  AOI220     g0547(.A0(new_new_n334_), .A1(new_new_n40_), .B0(new_new_n239_), .B1(new_new_n209_), .Y(new_new_n570_));
  OAI220     g0548(.A0(new_new_n570_), .A1(new_new_n555_), .B0(new_new_n569_), .B1(new_new_n247_), .Y(new_new_n571_));
  NA2        g0549(.A(new_new_n45_), .B(i_10_), .Y(new_new_n572_));
  NO2        g0550(.A(new_new_n572_), .B(i_6_), .Y(new_new_n573_));
  NA3        g0551(.A(new_new_n573_), .B(new_new_n571_), .C(new_new_n567_), .Y(new_new_n574_));
  NOi31      g0552(.An(new_new_n298_), .B(new_new_n309_), .C(new_new_n183_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n158_), .B(i_5_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n575_), .B(new_new_n483_), .Y(new_new_n577_));
  NA3        g0555(.A(new_new_n577_), .B(new_new_n574_), .C(new_new_n566_), .Y(new_new_n578_));
  NA3        g0556(.A(new_new_n221_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n579_));
  NA2        g0557(.A(new_new_n290_), .B(new_new_n85_), .Y(new_new_n580_));
  AOI210     g0558(.A0(new_new_n579_), .A1(new_new_n360_), .B0(new_new_n580_), .Y(new_new_n581_));
  NA2        g0559(.A(new_new_n304_), .B(new_new_n294_), .Y(new_new_n582_));
  NO2        g0560(.A(new_new_n582_), .B(new_new_n175_), .Y(new_new_n583_));
  NA2        g0561(.A(new_new_n227_), .B(new_new_n226_), .Y(new_new_n584_));
  NA2        g0562(.A(new_new_n469_), .B(new_new_n225_), .Y(new_new_n585_));
  NO2        g0563(.A(new_new_n584_), .B(new_new_n585_), .Y(new_new_n586_));
  AOI210     g0564(.A0(new_new_n380_), .A1(new_new_n47_), .B0(new_new_n384_), .Y(new_new_n587_));
  NA2        g0565(.A(i_0_), .B(new_new_n49_), .Y(new_new_n588_));
  NA3        g0566(.A(new_new_n561_), .B(new_new_n281_), .C(new_new_n588_), .Y(new_new_n589_));
  NO2        g0567(.A(new_new_n587_), .B(new_new_n589_), .Y(new_new_n590_));
  NO4        g0568(.A(new_new_n590_), .B(new_new_n586_), .C(new_new_n583_), .D(new_new_n581_), .Y(new_new_n591_));
  NO4        g0569(.A(new_new_n257_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n592_));
  NO3        g0570(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n237_), .B(new_new_n36_), .Y(new_new_n594_));
  AN2        g0572(.A(new_new_n594_), .B(new_new_n593_), .Y(new_new_n595_));
  OA210      g0573(.A0(new_new_n595_), .A1(new_new_n592_), .B0(new_new_n370_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n436_), .B(i_1_), .Y(new_new_n597_));
  NOi31      g0575(.An(new_new_n597_), .B(new_new_n475_), .C(new_new_n74_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n447_), .B(new_new_n179_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n599_), .B(new_new_n596_), .Y(new_new_n600_));
  NOi21      g0578(.An(i_10_), .B(i_6_), .Y(new_new_n601_));
  NO2        g0579(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n117_), .B(new_new_n23_), .Y(new_new_n603_));
  NA2        g0581(.A(new_new_n324_), .B(new_new_n165_), .Y(new_new_n604_));
  AOI220     g0582(.A0(new_new_n604_), .A1(new_new_n458_), .B0(new_new_n186_), .B1(new_new_n184_), .Y(new_new_n605_));
  NOi31      g0583(.An(new_new_n147_), .B(i_10_), .C(new_new_n341_), .Y(new_new_n606_));
  NO2        g0584(.A(new_new_n606_), .B(new_new_n605_), .Y(new_new_n607_));
  INV        g0585(.A(new_new_n327_), .Y(new_new_n608_));
  NO2        g0586(.A(i_12_), .B(new_new_n87_), .Y(new_new_n609_));
  NA3        g0587(.A(new_new_n609_), .B(new_new_n281_), .C(new_new_n588_), .Y(new_new_n610_));
  NA3        g0588(.A(new_new_n403_), .B(new_new_n290_), .C(new_new_n221_), .Y(new_new_n611_));
  AOI210     g0589(.A0(new_new_n611_), .A1(new_new_n610_), .B0(new_new_n608_), .Y(new_new_n612_));
  NA2        g0590(.A(new_new_n176_), .B(i_0_), .Y(new_new_n613_));
  NO3        g0591(.A(new_new_n613_), .B(new_new_n352_), .C(new_new_n309_), .Y(new_new_n614_));
  OR2        g0592(.A(i_2_), .B(i_5_), .Y(new_new_n615_));
  OR2        g0593(.A(new_new_n615_), .B(new_new_n428_), .Y(new_new_n616_));
  AOI210     g0594(.A0(new_new_n389_), .A1(new_new_n249_), .B0(new_new_n201_), .Y(new_new_n617_));
  AOI210     g0595(.A0(new_new_n617_), .A1(new_new_n616_), .B0(new_new_n522_), .Y(new_new_n618_));
  NO3        g0596(.A(new_new_n618_), .B(new_new_n614_), .C(new_new_n612_), .Y(new_new_n619_));
  NA4        g0597(.A(new_new_n619_), .B(new_new_n607_), .C(new_new_n600_), .D(new_new_n591_), .Y(new_new_n620_));
  NO4        g0598(.A(new_new_n620_), .B(new_new_n578_), .C(new_new_n558_), .D(new_new_n534_), .Y(new_new_n621_));
  NA4        g0599(.A(new_new_n621_), .B(new_new_n466_), .C(new_new_n369_), .D(new_new_n320_), .Y(men7));
  NO2        g0600(.A(new_new_n94_), .B(new_new_n55_), .Y(new_new_n623_));
  NO2        g0601(.A(new_new_n110_), .B(new_new_n91_), .Y(new_new_n624_));
  NA2        g0602(.A(new_new_n401_), .B(new_new_n624_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n509_), .B(new_new_n85_), .Y(new_new_n626_));
  NA2        g0604(.A(i_11_), .B(new_new_n196_), .Y(new_new_n627_));
  NA2        g0605(.A(new_new_n145_), .B(new_new_n627_), .Y(new_new_n628_));
  OAI210     g0606(.A0(new_new_n628_), .A1(new_new_n626_), .B0(new_new_n625_), .Y(new_new_n629_));
  NA3        g0607(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n241_), .B(i_4_), .Y(new_new_n631_));
  NA2        g0609(.A(new_new_n631_), .B(i_8_), .Y(new_new_n632_));
  NO2        g0610(.A(new_new_n107_), .B(new_new_n630_), .Y(new_new_n633_));
  NA2        g0611(.A(i_2_), .B(new_new_n87_), .Y(new_new_n634_));
  OAI210     g0612(.A0(new_new_n88_), .A1(new_new_n206_), .B0(new_new_n207_), .Y(new_new_n635_));
  NO2        g0613(.A(i_7_), .B(new_new_n37_), .Y(new_new_n636_));
  NA2        g0614(.A(i_4_), .B(i_8_), .Y(new_new_n637_));
  AOI210     g0615(.A0(new_new_n637_), .A1(new_new_n314_), .B0(new_new_n636_), .Y(new_new_n638_));
  OAI220     g0616(.A0(new_new_n638_), .A1(new_new_n634_), .B0(new_new_n635_), .B1(i_13_), .Y(new_new_n639_));
  NO4        g0617(.A(new_new_n639_), .B(new_new_n633_), .C(new_new_n629_), .D(new_new_n623_), .Y(new_new_n640_));
  AOI210     g0618(.A0(new_new_n129_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n641_));
  AOI210     g0619(.A0(new_new_n641_), .A1(new_new_n241_), .B0(new_new_n162_), .Y(new_new_n642_));
  OR2        g0620(.A(i_6_), .B(i_10_), .Y(new_new_n643_));
  NO2        g0621(.A(new_new_n643_), .B(new_new_n23_), .Y(new_new_n644_));
  OR3        g0622(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n645_));
  NO3        g0623(.A(new_new_n645_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n646_));
  INV        g0624(.A(new_new_n203_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n646_), .B(new_new_n644_), .Y(new_new_n648_));
  OA220      g0626(.A0(new_new_n648_), .A1(new_new_n608_), .B0(new_new_n642_), .B1(new_new_n276_), .Y(new_new_n649_));
  AOI210     g0627(.A0(new_new_n649_), .A1(new_new_n640_), .B0(new_new_n64_), .Y(new_new_n650_));
  NOi21      g0628(.An(i_11_), .B(i_7_), .Y(new_new_n651_));
  AO210      g0629(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n652_), .B(new_new_n651_), .Y(new_new_n653_));
  NA2        g0631(.A(new_new_n653_), .B(new_new_n209_), .Y(new_new_n654_));
  NA3        g0632(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n655_));
  NAi31      g0633(.An(new_new_n655_), .B(new_new_n218_), .C(i_11_), .Y(new_new_n656_));
  AOI210     g0634(.A0(new_new_n656_), .A1(new_new_n654_), .B0(new_new_n64_), .Y(new_new_n657_));
  OR2        g0635(.A(new_new_n395_), .B(new_new_n41_), .Y(new_new_n658_));
  NO3        g0636(.A(new_new_n265_), .B(new_new_n211_), .C(new_new_n627_), .Y(new_new_n659_));
  OAI210     g0637(.A0(new_new_n659_), .A1(new_new_n230_), .B0(new_new_n64_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n429_), .B(new_new_n31_), .Y(new_new_n661_));
  OR2        g0639(.A(new_new_n211_), .B(new_new_n110_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n662_), .B(new_new_n661_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n64_), .B(i_9_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n664_), .B(i_4_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n665_), .B(new_new_n663_), .Y(new_new_n666_));
  NO2        g0644(.A(i_1_), .B(i_12_), .Y(new_new_n667_));
  NA3        g0645(.A(new_new_n666_), .B(new_new_n660_), .C(new_new_n658_), .Y(new_new_n668_));
  OAI210     g0646(.A0(new_new_n668_), .A1(new_new_n657_), .B0(i_6_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n655_), .B(new_new_n110_), .Y(new_new_n670_));
  NA2        g0648(.A(new_new_n670_), .B(new_new_n609_), .Y(new_new_n671_));
  NO2        g0649(.A(new_new_n241_), .B(new_new_n87_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n672_), .B(i_11_), .Y(new_new_n673_));
  NA2        g0651(.A(new_new_n671_), .B(new_new_n476_), .Y(new_new_n674_));
  NO4        g0652(.A(new_new_n218_), .B(new_new_n129_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n675_), .B(new_new_n664_), .Y(new_new_n676_));
  NA2        g0654(.A(new_new_n241_), .B(i_6_), .Y(new_new_n677_));
  NO3        g0655(.A(new_new_n643_), .B(new_new_n237_), .C(new_new_n23_), .Y(new_new_n678_));
  AOI210     g0656(.A0(i_1_), .A1(new_new_n266_), .B0(new_new_n678_), .Y(new_new_n679_));
  OAI210     g0657(.A0(new_new_n679_), .A1(new_new_n45_), .B0(new_new_n676_), .Y(new_new_n680_));
  NA3        g0658(.A(new_new_n567_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n681_));
  NA2        g0659(.A(new_new_n139_), .B(i_9_), .Y(new_new_n682_));
  NA3        g0660(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n683_));
  NO2        g0661(.A(new_new_n47_), .B(i_1_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n682_), .B(new_new_n1092_), .Y(new_new_n685_));
  NA3        g0663(.A(new_new_n664_), .B(new_new_n327_), .C(i_6_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n686_), .B(new_new_n23_), .Y(new_new_n687_));
  AOI210     g0665(.A0(new_new_n500_), .A1(new_new_n440_), .B0(new_new_n246_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n688_), .B(new_new_n634_), .Y(new_new_n689_));
  NAi21      g0667(.An(new_new_n681_), .B(new_new_n93_), .Y(new_new_n690_));
  NA2        g0668(.A(new_new_n684_), .B(new_new_n275_), .Y(new_new_n691_));
  NO2        g0669(.A(i_11_), .B(new_new_n37_), .Y(new_new_n692_));
  NA2        g0670(.A(new_new_n692_), .B(new_new_n24_), .Y(new_new_n693_));
  OAI210     g0671(.A0(new_new_n693_), .A1(new_new_n691_), .B0(new_new_n690_), .Y(new_new_n694_));
  OR4        g0672(.A(new_new_n694_), .B(new_new_n689_), .C(new_new_n687_), .D(new_new_n685_), .Y(new_new_n695_));
  NO3        g0673(.A(new_new_n695_), .B(new_new_n680_), .C(new_new_n674_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n241_), .B(new_new_n103_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n697_), .B(new_new_n651_), .Y(new_new_n698_));
  NA2        g0676(.A(new_new_n698_), .B(i_1_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n699_), .B(new_new_n645_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n435_), .B(new_new_n87_), .Y(new_new_n701_));
  NA2        g0679(.A(new_new_n700_), .B(new_new_n47_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n237_), .B(new_new_n45_), .Y(new_new_n703_));
  NO3        g0681(.A(new_new_n703_), .B(new_new_n317_), .C(new_new_n242_), .Y(new_new_n704_));
  NO2        g0682(.A(new_new_n119_), .B(new_new_n37_), .Y(new_new_n705_));
  NO2        g0683(.A(new_new_n705_), .B(i_6_), .Y(new_new_n706_));
  NO2        g0684(.A(new_new_n87_), .B(i_9_), .Y(new_new_n707_));
  NO2        g0685(.A(new_new_n707_), .B(new_new_n64_), .Y(new_new_n708_));
  NO2        g0686(.A(new_new_n708_), .B(new_new_n667_), .Y(new_new_n709_));
  NO4        g0687(.A(new_new_n709_), .B(new_new_n706_), .C(new_new_n704_), .D(i_4_), .Y(new_new_n710_));
  NA2        g0688(.A(i_1_), .B(i_3_), .Y(new_new_n711_));
  INV        g0689(.A(new_new_n710_), .Y(new_new_n712_));
  NA4        g0690(.A(new_new_n712_), .B(new_new_n702_), .C(new_new_n696_), .D(new_new_n669_), .Y(new_new_n713_));
  AN2        g0691(.A(new_new_n250_), .B(new_new_n87_), .Y(new_new_n714_));
  NA2        g0692(.A(new_new_n387_), .B(new_new_n386_), .Y(new_new_n715_));
  NA3        g0693(.A(new_new_n509_), .B(new_new_n546_), .C(new_new_n47_), .Y(new_new_n716_));
  NO3        g0694(.A(new_new_n503_), .B(new_new_n637_), .C(new_new_n87_), .Y(new_new_n717_));
  NA2        g0695(.A(new_new_n717_), .B(new_new_n25_), .Y(new_new_n718_));
  NA3        g0696(.A(new_new_n162_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n719_));
  NA4        g0697(.A(new_new_n719_), .B(new_new_n718_), .C(new_new_n716_), .D(new_new_n715_), .Y(new_new_n720_));
  OAI210     g0698(.A0(new_new_n720_), .A1(new_new_n714_), .B0(i_1_), .Y(new_new_n721_));
  AOI210     g0699(.A0(new_new_n275_), .A1(new_new_n99_), .B0(i_1_), .Y(new_new_n722_));
  NO2        g0700(.A(new_new_n385_), .B(i_2_), .Y(new_new_n723_));
  NA2        g0701(.A(new_new_n723_), .B(new_new_n722_), .Y(new_new_n724_));
  OAI210     g0702(.A0(new_new_n686_), .A1(new_new_n470_), .B0(new_new_n724_), .Y(new_new_n725_));
  INV        g0703(.A(new_new_n725_), .Y(new_new_n726_));
  AOI210     g0704(.A0(new_new_n726_), .A1(new_new_n721_), .B0(i_13_), .Y(new_new_n727_));
  OR2        g0705(.A(i_11_), .B(i_7_), .Y(new_new_n728_));
  NA3        g0706(.A(new_new_n728_), .B(new_new_n108_), .C(new_new_n139_), .Y(new_new_n729_));
  AOI220     g0707(.A0(new_new_n495_), .A1(new_new_n162_), .B0(new_new_n472_), .B1(new_new_n139_), .Y(new_new_n730_));
  OAI210     g0708(.A0(new_new_n730_), .A1(new_new_n45_), .B0(new_new_n729_), .Y(new_new_n731_));
  AOI210     g0709(.A0(new_new_n683_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n732_));
  INV        g0710(.A(new_new_n732_), .Y(new_new_n733_));
  NO2        g0711(.A(new_new_n503_), .B(new_new_n24_), .Y(new_new_n734_));
  AOI220     g0712(.A0(new_new_n734_), .A1(new_new_n701_), .B0(new_new_n250_), .B1(new_new_n132_), .Y(new_new_n735_));
  OAI220     g0713(.A0(new_new_n735_), .A1(new_new_n41_), .B0(new_new_n733_), .B1(new_new_n94_), .Y(new_new_n736_));
  AOI210     g0714(.A0(new_new_n731_), .A1(new_new_n343_), .B0(new_new_n736_), .Y(new_new_n737_));
  INV        g0715(.A(new_new_n117_), .Y(new_new_n738_));
  AOI220     g0716(.A0(new_new_n738_), .A1(new_new_n73_), .B0(new_new_n403_), .B1(new_new_n684_), .Y(new_new_n739_));
  NO2        g0717(.A(new_new_n739_), .B(new_new_n247_), .Y(new_new_n740_));
  AOI210     g0718(.A0(new_new_n470_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n741_));
  NOi31      g0719(.An(new_new_n741_), .B(new_new_n626_), .C(new_new_n45_), .Y(new_new_n742_));
  NA2        g0720(.A(new_new_n128_), .B(i_13_), .Y(new_new_n743_));
  NO2        g0721(.A(new_new_n683_), .B(new_new_n117_), .Y(new_new_n744_));
  INV        g0722(.A(new_new_n744_), .Y(new_new_n745_));
  OAI220     g0723(.A0(new_new_n745_), .A1(new_new_n72_), .B0(new_new_n743_), .B1(new_new_n722_), .Y(new_new_n746_));
  NA2        g0724(.A(new_new_n26_), .B(new_new_n196_), .Y(new_new_n747_));
  NA2        g0725(.A(new_new_n747_), .B(i_7_), .Y(new_new_n748_));
  NO3        g0726(.A(new_new_n503_), .B(new_new_n241_), .C(new_new_n87_), .Y(new_new_n749_));
  NA2        g0727(.A(new_new_n749_), .B(new_new_n748_), .Y(new_new_n750_));
  AOI220     g0728(.A0(new_new_n403_), .A1(new_new_n684_), .B0(new_new_n93_), .B1(new_new_n104_), .Y(new_new_n751_));
  OAI220     g0729(.A0(new_new_n751_), .A1(new_new_n632_), .B0(new_new_n750_), .B1(new_new_n647_), .Y(new_new_n752_));
  NO4        g0730(.A(new_new_n752_), .B(new_new_n746_), .C(new_new_n742_), .D(new_new_n740_), .Y(new_new_n753_));
  OR2        g0731(.A(i_11_), .B(i_6_), .Y(new_new_n754_));
  NA3        g0732(.A(new_new_n631_), .B(new_new_n747_), .C(i_7_), .Y(new_new_n755_));
  AOI210     g0733(.A0(new_new_n755_), .A1(new_new_n745_), .B0(new_new_n754_), .Y(new_new_n756_));
  NA3        g0734(.A(new_new_n429_), .B(new_new_n636_), .C(new_new_n99_), .Y(new_new_n757_));
  NA2        g0735(.A(new_new_n673_), .B(i_13_), .Y(new_new_n758_));
  NA2        g0736(.A(new_new_n104_), .B(new_new_n747_), .Y(new_new_n759_));
  NAi21      g0737(.An(i_11_), .B(i_12_), .Y(new_new_n760_));
  NOi41      g0738(.An(new_new_n113_), .B(new_new_n760_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n761_));
  NO3        g0739(.A(new_new_n503_), .B(new_new_n609_), .C(new_new_n637_), .Y(new_new_n762_));
  AOI220     g0740(.A0(new_new_n762_), .A1(new_new_n321_), .B0(new_new_n761_), .B1(new_new_n759_), .Y(new_new_n763_));
  NA3        g0741(.A(new_new_n763_), .B(new_new_n758_), .C(new_new_n757_), .Y(new_new_n764_));
  OAI210     g0742(.A0(new_new_n764_), .A1(new_new_n756_), .B0(new_new_n64_), .Y(new_new_n765_));
  NO2        g0743(.A(i_2_), .B(i_12_), .Y(new_new_n766_));
  NA2        g0744(.A(new_new_n384_), .B(new_new_n766_), .Y(new_new_n767_));
  NA2        g0745(.A(i_8_), .B(new_new_n25_), .Y(new_new_n768_));
  NO3        g0746(.A(new_new_n768_), .B(new_new_n401_), .C(new_new_n631_), .Y(new_new_n769_));
  OAI210     g0747(.A0(new_new_n769_), .A1(new_new_n386_), .B0(new_new_n384_), .Y(new_new_n770_));
  NO2        g0748(.A(new_new_n129_), .B(i_2_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n771_), .B(new_new_n667_), .Y(new_new_n772_));
  NA3        g0750(.A(new_new_n772_), .B(new_new_n770_), .C(new_new_n767_), .Y(new_new_n773_));
  NA3        g0751(.A(new_new_n773_), .B(new_new_n46_), .C(new_new_n229_), .Y(new_new_n774_));
  NA4        g0752(.A(new_new_n774_), .B(new_new_n765_), .C(new_new_n753_), .D(new_new_n737_), .Y(new_new_n775_));
  OR4        g0753(.A(new_new_n775_), .B(new_new_n727_), .C(new_new_n713_), .D(new_new_n650_), .Y(men5));
  NA2        g0754(.A(new_new_n698_), .B(new_new_n278_), .Y(new_new_n777_));
  AN2        g0755(.A(new_new_n24_), .B(i_10_), .Y(new_new_n778_));
  NA3        g0756(.A(new_new_n778_), .B(new_new_n766_), .C(new_new_n110_), .Y(new_new_n779_));
  NO2        g0757(.A(new_new_n632_), .B(i_11_), .Y(new_new_n780_));
  NA2        g0758(.A(new_new_n88_), .B(new_new_n780_), .Y(new_new_n781_));
  NA3        g0759(.A(new_new_n781_), .B(new_new_n779_), .C(new_new_n777_), .Y(new_new_n782_));
  NO3        g0760(.A(i_11_), .B(new_new_n241_), .C(i_13_), .Y(new_new_n783_));
  NO2        g0761(.A(new_new_n125_), .B(new_new_n23_), .Y(new_new_n784_));
  NA2        g0762(.A(i_12_), .B(i_8_), .Y(new_new_n785_));
  OAI210     g0763(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n785_), .Y(new_new_n786_));
  INV        g0764(.A(new_new_n469_), .Y(new_new_n787_));
  AOI220     g0765(.A0(new_new_n327_), .A1(new_new_n603_), .B0(new_new_n786_), .B1(new_new_n784_), .Y(new_new_n788_));
  INV        g0766(.A(new_new_n788_), .Y(new_new_n789_));
  NO2        g0767(.A(new_new_n789_), .B(new_new_n782_), .Y(new_new_n790_));
  INV        g0768(.A(new_new_n173_), .Y(new_new_n791_));
  INV        g0769(.A(new_new_n250_), .Y(new_new_n792_));
  OAI210     g0770(.A0(new_new_n723_), .A1(new_new_n471_), .B0(new_new_n113_), .Y(new_new_n793_));
  AOI210     g0771(.A0(new_new_n793_), .A1(new_new_n792_), .B0(new_new_n791_), .Y(new_new_n794_));
  NO2        g0772(.A(new_new_n477_), .B(new_new_n26_), .Y(new_new_n795_));
  NO2        g0773(.A(new_new_n795_), .B(new_new_n440_), .Y(new_new_n796_));
  NA2        g0774(.A(new_new_n796_), .B(i_2_), .Y(new_new_n797_));
  INV        g0775(.A(new_new_n797_), .Y(new_new_n798_));
  AOI210     g0776(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n436_), .Y(new_new_n799_));
  AOI210     g0777(.A0(new_new_n799_), .A1(new_new_n798_), .B0(new_new_n794_), .Y(new_new_n800_));
  NO2        g0778(.A(new_new_n193_), .B(new_new_n126_), .Y(new_new_n801_));
  OAI210     g0779(.A0(new_new_n801_), .A1(new_new_n784_), .B0(i_2_), .Y(new_new_n802_));
  INV        g0780(.A(new_new_n174_), .Y(new_new_n803_));
  NO3        g0781(.A(new_new_n652_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n804_));
  AOI210     g0782(.A0(new_new_n803_), .A1(new_new_n88_), .B0(new_new_n804_), .Y(new_new_n805_));
  AOI210     g0783(.A0(new_new_n805_), .A1(new_new_n802_), .B0(new_new_n196_), .Y(new_new_n806_));
  OA210      g0784(.A0(new_new_n653_), .A1(new_new_n127_), .B0(i_13_), .Y(new_new_n807_));
  NA2        g0785(.A(new_new_n203_), .B(new_new_n206_), .Y(new_new_n808_));
  NA2        g0786(.A(new_new_n152_), .B(new_new_n627_), .Y(new_new_n809_));
  AOI210     g0787(.A0(new_new_n809_), .A1(new_new_n808_), .B0(new_new_n389_), .Y(new_new_n810_));
  AOI210     g0788(.A0(new_new_n211_), .A1(new_new_n149_), .B0(new_new_n546_), .Y(new_new_n811_));
  NA2        g0789(.A(new_new_n811_), .B(new_new_n440_), .Y(new_new_n812_));
  NO2        g0790(.A(new_new_n104_), .B(new_new_n45_), .Y(new_new_n813_));
  INV        g0791(.A(new_new_n310_), .Y(new_new_n814_));
  NA4        g0792(.A(new_new_n814_), .B(new_new_n314_), .C(new_new_n125_), .D(new_new_n43_), .Y(new_new_n815_));
  OAI210     g0793(.A0(new_new_n815_), .A1(new_new_n813_), .B0(new_new_n812_), .Y(new_new_n816_));
  NO4        g0794(.A(new_new_n816_), .B(new_new_n810_), .C(new_new_n807_), .D(new_new_n806_), .Y(new_new_n817_));
  NA2        g0795(.A(new_new_n603_), .B(new_new_n28_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n783_), .B(new_new_n282_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n819_), .B(new_new_n818_), .Y(new_new_n820_));
  NO2        g0798(.A(new_new_n63_), .B(i_12_), .Y(new_new_n821_));
  NO2        g0799(.A(new_new_n821_), .B(new_new_n127_), .Y(new_new_n822_));
  NO2        g0800(.A(new_new_n822_), .B(new_new_n627_), .Y(new_new_n823_));
  AOI220     g0801(.A0(new_new_n823_), .A1(new_new_n36_), .B0(new_new_n820_), .B1(new_new_n47_), .Y(new_new_n824_));
  NA4        g0802(.A(new_new_n824_), .B(new_new_n817_), .C(new_new_n800_), .D(new_new_n790_), .Y(men6));
  NO3        g0803(.A(new_new_n261_), .B(new_new_n316_), .C(i_1_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n188_), .B(new_new_n140_), .Y(new_new_n827_));
  OAI210     g0805(.A0(new_new_n827_), .A1(new_new_n826_), .B0(new_new_n771_), .Y(new_new_n828_));
  NA4        g0806(.A(new_new_n407_), .B(new_new_n508_), .C(new_new_n72_), .D(new_new_n103_), .Y(new_new_n829_));
  INV        g0807(.A(new_new_n829_), .Y(new_new_n830_));
  NO2        g0808(.A(new_new_n224_), .B(new_new_n513_), .Y(new_new_n831_));
  NO2        g0809(.A(i_11_), .B(i_9_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n830_), .B(new_new_n339_), .Y(new_new_n833_));
  AO210      g0811(.A0(new_new_n833_), .A1(new_new_n828_), .B0(i_12_), .Y(new_new_n834_));
  NA2        g0812(.A(new_new_n390_), .B(new_new_n346_), .Y(new_new_n835_));
  NA2        g0813(.A(new_new_n609_), .B(new_new_n64_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n836_), .B(new_new_n835_), .Y(new_new_n837_));
  INV        g0815(.A(new_new_n200_), .Y(new_new_n838_));
  AOI220     g0816(.A0(new_new_n838_), .A1(new_new_n832_), .B0(new_new_n837_), .B1(new_new_n74_), .Y(new_new_n839_));
  INV        g0817(.A(new_new_n338_), .Y(new_new_n840_));
  NA2        g0818(.A(new_new_n76_), .B(new_new_n132_), .Y(new_new_n841_));
  INV        g0819(.A(new_new_n125_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n842_), .B(new_new_n47_), .Y(new_new_n843_));
  AOI210     g0821(.A0(new_new_n843_), .A1(new_new_n841_), .B0(new_new_n840_), .Y(new_new_n844_));
  NO3        g0822(.A(new_new_n257_), .B(new_new_n133_), .C(i_9_), .Y(new_new_n845_));
  NA2        g0823(.A(new_new_n845_), .B(new_new_n821_), .Y(new_new_n846_));
  AOI210     g0824(.A0(new_new_n846_), .A1(new_new_n544_), .B0(new_new_n188_), .Y(new_new_n847_));
  NAi32      g0825(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n848_));
  NO2        g0826(.A(new_new_n754_), .B(new_new_n848_), .Y(new_new_n849_));
  OR3        g0827(.A(new_new_n849_), .B(new_new_n847_), .C(new_new_n844_), .Y(new_new_n850_));
  NO2        g0828(.A(new_new_n728_), .B(i_2_), .Y(new_new_n851_));
  NA2        g0829(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n852_));
  NO2        g0830(.A(new_new_n852_), .B(new_new_n428_), .Y(new_new_n853_));
  NA2        g0831(.A(new_new_n853_), .B(new_new_n851_), .Y(new_new_n854_));
  AO220      g0832(.A0(new_new_n374_), .A1(new_new_n364_), .B0(new_new_n415_), .B1(new_new_n627_), .Y(new_new_n855_));
  NA3        g0833(.A(new_new_n855_), .B(new_new_n262_), .C(i_7_), .Y(new_new_n856_));
  OR2        g0834(.A(new_new_n653_), .B(new_new_n471_), .Y(new_new_n857_));
  NA3        g0835(.A(new_new_n857_), .B(new_new_n148_), .C(new_new_n70_), .Y(new_new_n858_));
  AO210      g0836(.A0(new_new_n520_), .A1(new_new_n787_), .B0(new_new_n36_), .Y(new_new_n859_));
  NA4        g0837(.A(new_new_n859_), .B(new_new_n858_), .C(new_new_n856_), .D(new_new_n854_), .Y(new_new_n860_));
  NO2        g0838(.A(new_new_n672_), .B(i_11_), .Y(new_new_n861_));
  AOI220     g0839(.A0(new_new_n861_), .A1(new_new_n593_), .B0(new_new_n831_), .B1(new_new_n748_), .Y(new_new_n862_));
  NA3        g0840(.A(new_new_n389_), .B(new_new_n243_), .C(new_new_n148_), .Y(new_new_n863_));
  NA2        g0841(.A(new_new_n415_), .B(new_new_n71_), .Y(new_new_n864_));
  NA4        g0842(.A(new_new_n864_), .B(new_new_n863_), .C(new_new_n862_), .D(new_new_n635_), .Y(new_new_n865_));
  AOI210     g0843(.A0(new_new_n471_), .A1(new_new_n469_), .B0(new_new_n592_), .Y(new_new_n866_));
  NO2        g0844(.A(new_new_n643_), .B(new_new_n104_), .Y(new_new_n867_));
  OAI210     g0845(.A0(new_new_n867_), .A1(new_new_n114_), .B0(new_new_n426_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n249_), .B(new_new_n47_), .Y(new_new_n869_));
  INV        g0847(.A(new_new_n616_), .Y(new_new_n870_));
  NA3        g0848(.A(new_new_n870_), .B(new_new_n338_), .C(i_7_), .Y(new_new_n871_));
  NA3        g0849(.A(new_new_n871_), .B(new_new_n868_), .C(new_new_n866_), .Y(new_new_n872_));
  NO4        g0850(.A(new_new_n872_), .B(new_new_n865_), .C(new_new_n860_), .D(new_new_n850_), .Y(new_new_n873_));
  NA4        g0851(.A(new_new_n873_), .B(new_new_n839_), .C(new_new_n834_), .D(new_new_n397_), .Y(men3));
  NA2        g0852(.A(i_12_), .B(i_10_), .Y(new_new_n875_));
  NA2        g0853(.A(i_6_), .B(i_7_), .Y(new_new_n876_));
  NO2        g0854(.A(new_new_n876_), .B(i_0_), .Y(new_new_n877_));
  NO2        g0855(.A(i_11_), .B(new_new_n241_), .Y(new_new_n878_));
  OAI210     g0856(.A0(new_new_n877_), .A1(new_new_n298_), .B0(new_new_n878_), .Y(new_new_n879_));
  NO2        g0857(.A(new_new_n879_), .B(new_new_n196_), .Y(new_new_n880_));
  NO3        g0858(.A(new_new_n473_), .B(new_new_n91_), .C(new_new_n45_), .Y(new_new_n881_));
  OA210      g0859(.A0(new_new_n881_), .A1(new_new_n880_), .B0(new_new_n176_), .Y(new_new_n882_));
  NA2        g0860(.A(new_new_n863_), .B(new_new_n388_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n883_), .B(new_new_n40_), .Y(new_new_n884_));
  NOi21      g0862(.An(new_new_n98_), .B(new_new_n796_), .Y(new_new_n885_));
  NO3        g0863(.A(new_new_n662_), .B(new_new_n477_), .C(new_new_n132_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n429_), .B(new_new_n46_), .Y(new_new_n887_));
  AN2        g0865(.A(new_new_n475_), .B(new_new_n56_), .Y(new_new_n888_));
  NO3        g0866(.A(new_new_n888_), .B(new_new_n886_), .C(new_new_n885_), .Y(new_new_n889_));
  AOI210     g0867(.A0(new_new_n889_), .A1(new_new_n884_), .B0(new_new_n49_), .Y(new_new_n890_));
  NO4        g0868(.A(new_new_n393_), .B(new_new_n400_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n188_), .B(new_new_n601_), .Y(new_new_n892_));
  NOi21      g0870(.An(new_new_n892_), .B(new_new_n891_), .Y(new_new_n893_));
  NA2        g0871(.A(new_new_n741_), .B(new_new_n707_), .Y(new_new_n894_));
  NA2        g0872(.A(new_new_n344_), .B(new_new_n460_), .Y(new_new_n895_));
  OAI220     g0873(.A0(new_new_n895_), .A1(new_new_n894_), .B0(new_new_n893_), .B1(new_new_n64_), .Y(new_new_n896_));
  NOi21      g0874(.An(i_5_), .B(i_9_), .Y(new_new_n897_));
  NA2        g0875(.A(new_new_n897_), .B(new_new_n468_), .Y(new_new_n898_));
  BUFFER     g0876(.A(new_new_n275_), .Y(new_new_n899_));
  AOI210     g0877(.A0(new_new_n899_), .A1(new_new_n500_), .B0(new_new_n717_), .Y(new_new_n900_));
  NO2        g0878(.A(new_new_n177_), .B(new_new_n149_), .Y(new_new_n901_));
  NO2        g0879(.A(new_new_n900_), .B(new_new_n898_), .Y(new_new_n902_));
  NO4        g0880(.A(new_new_n902_), .B(new_new_n896_), .C(new_new_n890_), .D(new_new_n882_), .Y(new_new_n903_));
  NA2        g0881(.A(new_new_n188_), .B(new_new_n24_), .Y(new_new_n904_));
  NA2        g0882(.A(new_new_n321_), .B(new_new_n130_), .Y(new_new_n905_));
  NAi21      g0883(.An(new_new_n163_), .B(new_new_n460_), .Y(new_new_n906_));
  OAI220     g0884(.A0(new_new_n906_), .A1(new_new_n869_), .B0(new_new_n905_), .B1(new_new_n418_), .Y(new_new_n907_));
  INV        g0885(.A(new_new_n907_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n407_), .B(new_new_n302_), .Y(new_new_n909_));
  NA2        g0887(.A(new_new_n909_), .B(new_new_n744_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n602_), .B(i_0_), .Y(new_new_n911_));
  NO4        g0889(.A(new_new_n615_), .B(new_new_n218_), .C(new_new_n436_), .D(new_new_n428_), .Y(new_new_n912_));
  NA2        g0890(.A(new_new_n912_), .B(i_11_), .Y(new_new_n913_));
  INV        g0891(.A(new_new_n498_), .Y(new_new_n914_));
  AN2        g0892(.A(new_new_n98_), .B(new_new_n248_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n783_), .B(new_new_n339_), .Y(new_new_n916_));
  AOI210     g0894(.A0(new_new_n509_), .A1(new_new_n88_), .B0(new_new_n59_), .Y(new_new_n917_));
  OAI220     g0895(.A0(new_new_n917_), .A1(new_new_n916_), .B0(new_new_n693_), .B1(new_new_n569_), .Y(new_new_n918_));
  NO2        g0896(.A(new_new_n259_), .B(new_new_n154_), .Y(new_new_n919_));
  NA2        g0897(.A(i_0_), .B(i_10_), .Y(new_new_n920_));
  AN2        g0898(.A(new_new_n919_), .B(i_6_), .Y(new_new_n921_));
  AOI220     g0899(.A0(new_new_n344_), .A1(new_new_n100_), .B0(new_new_n188_), .B1(new_new_n85_), .Y(new_new_n922_));
  NA2        g0900(.A(new_new_n597_), .B(i_4_), .Y(new_new_n923_));
  NO2        g0901(.A(new_new_n923_), .B(new_new_n922_), .Y(new_new_n924_));
  NO4        g0902(.A(new_new_n924_), .B(new_new_n921_), .C(new_new_n918_), .D(new_new_n915_), .Y(new_new_n925_));
  NA4        g0903(.A(new_new_n925_), .B(new_new_n913_), .C(new_new_n910_), .D(new_new_n908_), .Y(new_new_n926_));
  NA2        g0904(.A(i_11_), .B(i_9_), .Y(new_new_n927_));
  NO2        g0905(.A(new_new_n49_), .B(i_7_), .Y(new_new_n928_));
  NA2        g0906(.A(new_new_n412_), .B(new_new_n181_), .Y(new_new_n929_));
  NA2        g0907(.A(new_new_n929_), .B(new_new_n161_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n927_), .B(new_new_n74_), .Y(new_new_n931_));
  NO2        g0909(.A(new_new_n177_), .B(i_0_), .Y(new_new_n932_));
  INV        g0910(.A(new_new_n932_), .Y(new_new_n933_));
  NA2        g0911(.A(new_new_n498_), .B(new_new_n235_), .Y(new_new_n934_));
  AOI210     g0912(.A0(new_new_n387_), .A1(new_new_n42_), .B0(new_new_n425_), .Y(new_new_n935_));
  OAI220     g0913(.A0(new_new_n935_), .A1(new_new_n898_), .B0(new_new_n934_), .B1(new_new_n933_), .Y(new_new_n936_));
  NO2        g0914(.A(new_new_n936_), .B(new_new_n930_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n692_), .B(new_new_n122_), .Y(new_new_n938_));
  NO2        g0916(.A(i_6_), .B(new_new_n938_), .Y(new_new_n939_));
  AOI210     g0917(.A0(new_new_n470_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n940_));
  NA2        g0918(.A(new_new_n173_), .B(new_new_n105_), .Y(new_new_n941_));
  NOi32      g0919(.An(new_new_n940_), .Bn(new_new_n191_), .C(new_new_n941_), .Y(new_new_n942_));
  NA2        g0920(.A(new_new_n636_), .B(new_new_n339_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n943_), .B(new_new_n887_), .Y(new_new_n944_));
  NO3        g0922(.A(new_new_n944_), .B(new_new_n942_), .C(new_new_n939_), .Y(new_new_n945_));
  NOi21      g0923(.An(i_7_), .B(i_5_), .Y(new_new_n946_));
  NOi31      g0924(.An(new_new_n946_), .B(i_0_), .C(new_new_n760_), .Y(new_new_n947_));
  NA3        g0925(.A(new_new_n947_), .B(new_new_n401_), .C(i_6_), .Y(new_new_n948_));
  OA210      g0926(.A0(new_new_n941_), .A1(new_new_n544_), .B0(new_new_n948_), .Y(new_new_n949_));
  NO3        g0927(.A(new_new_n421_), .B(new_new_n377_), .C(new_new_n373_), .Y(new_new_n950_));
  NO2        g0928(.A(new_new_n269_), .B(new_new_n328_), .Y(new_new_n951_));
  NO2        g0929(.A(new_new_n760_), .B(new_new_n264_), .Y(new_new_n952_));
  AOI210     g0930(.A0(new_new_n952_), .A1(new_new_n951_), .B0(new_new_n950_), .Y(new_new_n953_));
  NA4        g0931(.A(new_new_n953_), .B(new_new_n949_), .C(new_new_n945_), .D(new_new_n937_), .Y(new_new_n954_));
  NO2        g0932(.A(new_new_n904_), .B(new_new_n244_), .Y(new_new_n955_));
  AN2        g0933(.A(new_new_n343_), .B(new_new_n339_), .Y(new_new_n956_));
  AN2        g0934(.A(new_new_n956_), .B(new_new_n901_), .Y(new_new_n957_));
  OAI210     g0935(.A0(new_new_n957_), .A1(new_new_n955_), .B0(i_10_), .Y(new_new_n958_));
  NO2        g0936(.A(new_new_n875_), .B(new_new_n327_), .Y(new_new_n959_));
  NA2        g0937(.A(new_new_n959_), .B(new_new_n931_), .Y(new_new_n960_));
  NA3        g0938(.A(new_new_n497_), .B(new_new_n429_), .C(new_new_n46_), .Y(new_new_n961_));
  OAI210     g0939(.A0(new_new_n906_), .A1(new_new_n914_), .B0(new_new_n961_), .Y(new_new_n962_));
  NO2        g0940(.A(new_new_n262_), .B(new_new_n47_), .Y(new_new_n963_));
  NA2        g0941(.A(new_new_n931_), .B(new_new_n314_), .Y(new_new_n964_));
  OAI210     g0942(.A0(new_new_n963_), .A1(new_new_n190_), .B0(new_new_n964_), .Y(new_new_n965_));
  AOI220     g0943(.A0(new_new_n965_), .A1(new_new_n498_), .B0(new_new_n962_), .B1(new_new_n74_), .Y(new_new_n966_));
  NA3        g0944(.A(new_new_n852_), .B(new_new_n399_), .C(new_new_n672_), .Y(new_new_n967_));
  NO2        g0945(.A(new_new_n967_), .B(new_new_n48_), .Y(new_new_n968_));
  NO3        g0946(.A(new_new_n615_), .B(new_new_n372_), .C(new_new_n24_), .Y(new_new_n969_));
  AOI210     g0947(.A0(new_new_n734_), .A1(new_new_n576_), .B0(new_new_n969_), .Y(new_new_n970_));
  NAi21      g0948(.An(i_9_), .B(i_5_), .Y(new_new_n971_));
  NO2        g0949(.A(new_new_n971_), .B(new_new_n421_), .Y(new_new_n972_));
  NO2        g0950(.A(new_new_n630_), .B(new_new_n107_), .Y(new_new_n973_));
  AOI220     g0951(.A0(new_new_n973_), .A1(i_0_), .B0(new_new_n972_), .B1(new_new_n653_), .Y(new_new_n974_));
  OAI220     g0952(.A0(new_new_n974_), .A1(new_new_n87_), .B0(new_new_n970_), .B1(new_new_n174_), .Y(new_new_n975_));
  NO3        g0953(.A(new_new_n975_), .B(new_new_n968_), .C(new_new_n549_), .Y(new_new_n976_));
  NA4        g0954(.A(new_new_n976_), .B(new_new_n966_), .C(new_new_n960_), .D(new_new_n958_), .Y(new_new_n977_));
  NO3        g0955(.A(new_new_n977_), .B(new_new_n954_), .C(new_new_n926_), .Y(new_new_n978_));
  NO2        g0956(.A(i_0_), .B(new_new_n760_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n980_));
  NA2        g0958(.A(new_new_n920_), .B(new_new_n980_), .Y(new_new_n981_));
  NO3        g0959(.A(new_new_n107_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n982_));
  AO220      g0960(.A0(new_new_n982_), .A1(new_new_n981_), .B0(new_new_n979_), .B1(new_new_n176_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n836_), .A1(new_new_n715_), .B0(new_new_n941_), .Y(new_new_n984_));
  AOI210     g0962(.A0(new_new_n983_), .A1(new_new_n361_), .B0(new_new_n984_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n771_), .B(new_new_n147_), .Y(new_new_n986_));
  INV        g0964(.A(new_new_n986_), .Y(new_new_n987_));
  NA3        g0965(.A(new_new_n987_), .B(new_new_n707_), .C(new_new_n74_), .Y(new_new_n988_));
  NA3        g0966(.A(new_new_n877_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n989_));
  NA2        g0967(.A(new_new_n878_), .B(i_9_), .Y(new_new_n990_));
  AOI210     g0968(.A0(new_new_n989_), .A1(new_new_n525_), .B0(new_new_n990_), .Y(new_new_n991_));
  OAI210     g0969(.A0(new_new_n249_), .A1(i_9_), .B0(new_new_n234_), .Y(new_new_n992_));
  AOI210     g0970(.A0(new_new_n992_), .A1(new_new_n911_), .B0(new_new_n154_), .Y(new_new_n993_));
  NO2        g0971(.A(new_new_n993_), .B(new_new_n991_), .Y(new_new_n994_));
  NA3        g0972(.A(new_new_n994_), .B(new_new_n988_), .C(new_new_n985_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n956_), .B(new_new_n389_), .Y(new_new_n996_));
  AOI210     g0974(.A0(new_new_n309_), .A1(new_new_n163_), .B0(new_new_n996_), .Y(new_new_n997_));
  NA3        g0975(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n998_));
  NA2        g0976(.A(new_new_n928_), .B(new_new_n514_), .Y(new_new_n999_));
  AOI210     g0977(.A0(new_new_n998_), .A1(new_new_n163_), .B0(new_new_n999_), .Y(new_new_n1000_));
  NO2        g0978(.A(new_new_n1000_), .B(new_new_n997_), .Y(new_new_n1001_));
  NO3        g0979(.A(new_new_n920_), .B(new_new_n897_), .C(new_new_n193_), .Y(new_new_n1002_));
  AOI220     g0980(.A0(new_new_n1002_), .A1(i_11_), .B0(new_new_n598_), .B1(new_new_n76_), .Y(new_new_n1003_));
  NO3        g0981(.A(new_new_n212_), .B(new_new_n400_), .C(i_0_), .Y(new_new_n1004_));
  OAI210     g0982(.A0(new_new_n1004_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n1005_));
  INV        g0983(.A(new_new_n221_), .Y(new_new_n1006_));
  OAI220     g0984(.A0(new_new_n562_), .A1(new_new_n140_), .B0(new_new_n677_), .B1(new_new_n647_), .Y(new_new_n1007_));
  NA3        g0985(.A(new_new_n1007_), .B(new_new_n416_), .C(new_new_n1006_), .Y(new_new_n1008_));
  NA4        g0986(.A(new_new_n1008_), .B(new_new_n1005_), .C(new_new_n1003_), .D(new_new_n1001_), .Y(new_new_n1009_));
  INV        g0987(.A(new_new_n111_), .Y(new_new_n1010_));
  AOI220     g0988(.A0(new_new_n946_), .A1(new_new_n514_), .B0(new_new_n877_), .B1(new_new_n164_), .Y(new_new_n1011_));
  NA2        g0989(.A(new_new_n364_), .B(new_new_n178_), .Y(new_new_n1012_));
  OA220      g0990(.A0(new_new_n1012_), .A1(new_new_n1011_), .B0(new_new_n1010_), .B1(i_5_), .Y(new_new_n1013_));
  NA3        g0991(.A(new_new_n644_), .B(new_new_n188_), .C(new_new_n85_), .Y(new_new_n1014_));
  INV        g0992(.A(new_new_n1014_), .Y(new_new_n1015_));
  NO3        g0993(.A(new_new_n887_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n1016_));
  NA2        g0994(.A(new_new_n519_), .B(new_new_n512_), .Y(new_new_n1017_));
  NO3        g0995(.A(new_new_n1017_), .B(new_new_n1016_), .C(new_new_n1015_), .Y(new_new_n1018_));
  NA3        g0996(.A(new_new_n407_), .B(new_new_n173_), .C(new_new_n172_), .Y(new_new_n1019_));
  NA3        g0997(.A(new_new_n928_), .B(new_new_n298_), .C(new_new_n234_), .Y(new_new_n1020_));
  NA2        g0998(.A(new_new_n1020_), .B(new_new_n1019_), .Y(new_new_n1021_));
  NA3        g0999(.A(new_new_n407_), .B(new_new_n345_), .C(new_new_n225_), .Y(new_new_n1022_));
  INV        g1000(.A(new_new_n1022_), .Y(new_new_n1023_));
  NOi31      g1001(.An(new_new_n406_), .B(new_new_n980_), .C(new_new_n244_), .Y(new_new_n1024_));
  NO3        g1002(.A(new_new_n927_), .B(new_new_n221_), .C(new_new_n193_), .Y(new_new_n1025_));
  NO4        g1003(.A(new_new_n1025_), .B(new_new_n1024_), .C(new_new_n1023_), .D(new_new_n1021_), .Y(new_new_n1026_));
  NA3        g1004(.A(new_new_n1026_), .B(new_new_n1018_), .C(new_new_n1013_), .Y(new_new_n1027_));
  INV        g1005(.A(new_new_n646_), .Y(new_new_n1028_));
  NO3        g1006(.A(new_new_n1028_), .B(new_new_n588_), .C(new_new_n358_), .Y(new_new_n1029_));
  NO2        g1007(.A(new_new_n87_), .B(i_5_), .Y(new_new_n1030_));
  NA3        g1008(.A(new_new_n878_), .B(new_new_n112_), .C(new_new_n125_), .Y(new_new_n1031_));
  INV        g1009(.A(new_new_n1031_), .Y(new_new_n1032_));
  AOI210     g1010(.A0(new_new_n1032_), .A1(new_new_n1030_), .B0(new_new_n1029_), .Y(new_new_n1033_));
  NAi21      g1011(.An(new_new_n246_), .B(new_new_n247_), .Y(new_new_n1034_));
  NO4        g1012(.A(new_new_n244_), .B(new_new_n212_), .C(i_0_), .D(i_12_), .Y(new_new_n1035_));
  AOI220     g1013(.A0(new_new_n1035_), .A1(new_new_n1034_), .B0(new_new_n830_), .B1(new_new_n178_), .Y(new_new_n1036_));
  AN2        g1014(.A(new_new_n920_), .B(new_new_n154_), .Y(new_new_n1037_));
  NO4        g1015(.A(new_new_n1037_), .B(i_12_), .C(new_new_n681_), .D(new_new_n132_), .Y(new_new_n1038_));
  NA2        g1016(.A(new_new_n1038_), .B(new_new_n221_), .Y(new_new_n1039_));
  NA3        g1017(.A(new_new_n100_), .B(new_new_n601_), .C(i_11_), .Y(new_new_n1040_));
  NO2        g1018(.A(new_new_n1040_), .B(new_new_n156_), .Y(new_new_n1041_));
  NA2        g1019(.A(new_new_n946_), .B(new_new_n495_), .Y(new_new_n1042_));
  NO2        g1020(.A(new_new_n1042_), .B(new_new_n708_), .Y(new_new_n1043_));
  AOI210     g1021(.A0(new_new_n1043_), .A1(new_new_n932_), .B0(new_new_n1041_), .Y(new_new_n1044_));
  NA4        g1022(.A(new_new_n1044_), .B(new_new_n1039_), .C(new_new_n1036_), .D(new_new_n1033_), .Y(new_new_n1045_));
  NO4        g1023(.A(new_new_n1045_), .B(new_new_n1027_), .C(new_new_n1009_), .D(new_new_n995_), .Y(new_new_n1046_));
  NA2        g1024(.A(new_new_n851_), .B(new_new_n37_), .Y(new_new_n1047_));
  NA3        g1025(.A(new_new_n940_), .B(new_new_n384_), .C(i_5_), .Y(new_new_n1048_));
  NA3        g1026(.A(new_new_n1048_), .B(new_new_n1047_), .C(new_new_n642_), .Y(new_new_n1049_));
  NA2        g1027(.A(new_new_n1049_), .B(new_new_n209_), .Y(new_new_n1050_));
  AN2        g1028(.A(new_new_n728_), .B(new_new_n385_), .Y(new_new_n1051_));
  NA2        g1029(.A(new_new_n189_), .B(new_new_n191_), .Y(new_new_n1052_));
  AO210      g1030(.A0(new_new_n1051_), .A1(new_new_n33_), .B0(new_new_n1052_), .Y(new_new_n1053_));
  OAI210     g1031(.A0(new_new_n646_), .A1(new_new_n644_), .B0(new_new_n327_), .Y(new_new_n1054_));
  NAi31      g1032(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1055_));
  NO2        g1033(.A(new_new_n71_), .B(new_new_n1055_), .Y(new_new_n1056_));
  NO2        g1034(.A(new_new_n1056_), .B(new_new_n678_), .Y(new_new_n1057_));
  NA3        g1035(.A(new_new_n1057_), .B(new_new_n1054_), .C(new_new_n1053_), .Y(new_new_n1058_));
  NO4        g1036(.A(new_new_n237_), .B(new_new_n146_), .C(new_new_n711_), .D(new_new_n37_), .Y(new_new_n1059_));
  NO2        g1037(.A(new_new_n1059_), .B(new_new_n912_), .Y(new_new_n1060_));
  OAI210     g1038(.A0(new_new_n1040_), .A1(new_new_n149_), .B0(new_new_n1060_), .Y(new_new_n1061_));
  AOI210     g1039(.A0(new_new_n1058_), .A1(new_new_n49_), .B0(new_new_n1061_), .Y(new_new_n1062_));
  AOI210     g1040(.A0(new_new_n1062_), .A1(new_new_n1050_), .B0(new_new_n74_), .Y(new_new_n1063_));
  NO2        g1041(.A(new_new_n595_), .B(new_new_n396_), .Y(new_new_n1064_));
  NO2        g1042(.A(new_new_n1064_), .B(new_new_n791_), .Y(new_new_n1065_));
  OAI210     g1043(.A0(new_new_n81_), .A1(new_new_n55_), .B0(new_new_n110_), .Y(new_new_n1066_));
  NA2        g1044(.A(new_new_n1066_), .B(new_new_n77_), .Y(new_new_n1067_));
  INV        g1045(.A(new_new_n947_), .Y(new_new_n1068_));
  AOI210     g1046(.A0(new_new_n1068_), .A1(new_new_n1067_), .B0(new_new_n711_), .Y(new_new_n1069_));
  NA2        g1047(.A(new_new_n269_), .B(new_new_n58_), .Y(new_new_n1070_));
  AOI220     g1048(.A0(new_new_n1070_), .A1(new_new_n77_), .B0(new_new_n359_), .B1(new_new_n261_), .Y(new_new_n1071_));
  NO2        g1049(.A(new_new_n1071_), .B(new_new_n241_), .Y(new_new_n1072_));
  NA3        g1050(.A(new_new_n98_), .B(new_new_n316_), .C(new_new_n31_), .Y(new_new_n1073_));
  INV        g1051(.A(new_new_n1073_), .Y(new_new_n1074_));
  NO3        g1052(.A(new_new_n1074_), .B(new_new_n1072_), .C(new_new_n1069_), .Y(new_new_n1075_));
  OAI210     g1053(.A0(new_new_n277_), .A1(new_new_n159_), .B0(new_new_n88_), .Y(new_new_n1076_));
  NA3        g1054(.A(new_new_n795_), .B(new_new_n298_), .C(new_new_n81_), .Y(new_new_n1077_));
  AOI210     g1055(.A0(new_new_n1077_), .A1(new_new_n1076_), .B0(i_11_), .Y(new_new_n1078_));
  NA2        g1056(.A(new_new_n637_), .B(new_new_n218_), .Y(new_new_n1079_));
  OAI210     g1057(.A0(new_new_n1079_), .A1(new_new_n940_), .B0(new_new_n209_), .Y(new_new_n1080_));
  NA2        g1058(.A(new_new_n165_), .B(i_5_), .Y(new_new_n1081_));
  NO2        g1059(.A(new_new_n1080_), .B(new_new_n1081_), .Y(new_new_n1082_));
  NO4        g1060(.A(new_new_n971_), .B(new_new_n502_), .C(new_new_n258_), .D(new_new_n257_), .Y(new_new_n1083_));
  NO2        g1061(.A(new_new_n1083_), .B(new_new_n592_), .Y(new_new_n1084_));
  NO2        g1062(.A(new_new_n1084_), .B(new_new_n41_), .Y(new_new_n1085_));
  NO3        g1063(.A(new_new_n1085_), .B(new_new_n1082_), .C(new_new_n1078_), .Y(new_new_n1086_));
  OAI210     g1064(.A0(new_new_n1075_), .A1(i_4_), .B0(new_new_n1086_), .Y(new_new_n1087_));
  NO3        g1065(.A(new_new_n1087_), .B(new_new_n1065_), .C(new_new_n1063_), .Y(new_new_n1088_));
  NA4        g1066(.A(new_new_n1088_), .B(new_new_n1046_), .C(new_new_n978_), .D(new_new_n903_), .Y(men4));
  INV        g1067(.A(i_2_), .Y(new_new_n1092_));
  INV        g1068(.A(new_new_n119_), .Y(new_new_n1093_));
endmodule


