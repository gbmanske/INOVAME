//Benchmark atmr_misex3_1774_0.0156

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1374_, ori_ori_n1375_, ori_ori_n1376_, ori_ori_n1377_, ori_ori_n1378_, ori_ori_n1379_, ori_ori_n1380_, ori_ori_n1381_, ori_ori_n1382_, ori_ori_n1383_, ori_ori_n1384_, ori_ori_n1385_, ori_ori_n1386_, ori_ori_n1387_, ori_ori_n1388_, ori_ori_n1389_, ori_ori_n1390_, ori_ori_n1391_, ori_ori_n1392_, ori_ori_n1393_, ori_ori_n1394_, ori_ori_n1395_, ori_ori_n1396_, ori_ori_n1397_, ori_ori_n1398_, ori_ori_n1399_, ori_ori_n1400_, ori_ori_n1401_, ori_ori_n1402_, ori_ori_n1403_, ori_ori_n1404_, ori_ori_n1405_, ori_ori_n1406_, ori_ori_n1407_, ori_ori_n1408_, ori_ori_n1409_, ori_ori_n1410_, ori_ori_n1411_, ori_ori_n1412_, ori_ori_n1413_, ori_ori_n1414_, ori_ori_n1415_, ori_ori_n1416_, ori_ori_n1417_, ori_ori_n1418_, ori_ori_n1419_, ori_ori_n1420_, ori_ori_n1421_, ori_ori_n1422_, ori_ori_n1423_, ori_ori_n1424_, ori_ori_n1425_, ori_ori_n1426_, ori_ori_n1427_, ori_ori_n1428_, ori_ori_n1429_, ori_ori_n1430_, ori_ori_n1431_, ori_ori_n1432_, ori_ori_n1433_, ori_ori_n1434_, ori_ori_n1435_, ori_ori_n1436_, ori_ori_n1437_, ori_ori_n1438_, ori_ori_n1439_, ori_ori_n1440_, ori_ori_n1441_, ori_ori_n1442_, ori_ori_n1443_, ori_ori_n1444_, ori_ori_n1445_, ori_ori_n1446_, ori_ori_n1447_, ori_ori_n1448_, ori_ori_n1449_, ori_ori_n1450_, ori_ori_n1451_, ori_ori_n1452_, ori_ori_n1453_, ori_ori_n1454_, ori_ori_n1455_, ori_ori_n1456_, ori_ori_n1457_, ori_ori_n1458_, ori_ori_n1459_, ori_ori_n1460_, ori_ori_n1461_, ori_ori_n1462_, ori_ori_n1463_, ori_ori_n1464_, ori_ori_n1465_, ori_ori_n1466_, ori_ori_n1467_, ori_ori_n1469_, ori_ori_n1470_, ori_ori_n1471_, ori_ori_n1472_, ori_ori_n1476_, ori_ori_n1477_, ori_ori_n1478_, ori_ori_n1479_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1521_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1533_, mai_mai_n1534_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1540_, mai_mai_n1541_, mai_mai_n1542_, mai_mai_n1543_, mai_mai_n1547_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1562_, men_men_n1563_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  NO2        o0001(.A(d), .B(c), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(o), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(o), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  NO2        o0010(.A(ori_ori_n38_), .B(n), .Y(ori_ori_n39_));
  INV        o0011(.A(h), .Y(ori_ori_n40_));
  NAi21      o0012(.An(j), .B(l), .Y(ori_ori_n41_));
  NAi32      o0013(.An(n), .Bn(o), .C(m), .Y(ori_ori_n42_));
  NO3        o0014(.A(ori_ori_n42_), .B(ori_ori_n41_), .C(ori_ori_n40_), .Y(ori_ori_n43_));
  NAi31      o0015(.An(n), .B(m), .C(l), .Y(ori_ori_n44_));
  INV        o0016(.A(i), .Y(ori_ori_n45_));
  AN2        o0017(.A(h), .B(o), .Y(ori_ori_n46_));
  NA2        o0018(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o0019(.A(ori_ori_n47_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NAi21      o0020(.An(n), .B(m), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(l), .Y(ori_ori_n50_));
  NOi32      o0022(.An(k), .Bn(h), .C(o), .Y(ori_ori_n51_));
  INV        o0023(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NO2        o0024(.A(ori_ori_n52_), .B(ori_ori_n49_), .Y(ori_ori_n53_));
  NO4        o0025(.A(ori_ori_n53_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n54_));
  AOI210     o0026(.A0(ori_ori_n54_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n55_));
  INV        o0027(.A(c), .Y(ori_ori_n56_));
  NA2        o0028(.A(e), .B(b), .Y(ori_ori_n57_));
  NO2        o0029(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0030(.A(d), .Y(ori_ori_n59_));
  NA2        o0031(.A(o), .B(ori_ori_n59_), .Y(ori_ori_n60_));
  NAi21      o0032(.An(i), .B(h), .Y(ori_ori_n61_));
  NAi31      o0033(.An(i), .B(l), .C(j), .Y(ori_ori_n62_));
  OAI220     o0034(.A0(ori_ori_n62_), .A1(ori_ori_n49_), .B0(ori_ori_n61_), .B1(ori_ori_n44_), .Y(ori_ori_n63_));
  NAi31      o0035(.An(ori_ori_n60_), .B(ori_ori_n63_), .C(ori_ori_n58_), .Y(ori_ori_n64_));
  NAi41      o0036(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n65_));
  NA2        o0037(.A(o), .B(f), .Y(ori_ori_n66_));
  NO2        o0038(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n67_));
  NAi21      o0039(.An(i), .B(j), .Y(ori_ori_n68_));
  NAi32      o0040(.An(n), .Bn(k), .C(m), .Y(ori_ori_n69_));
  NAi31      o0041(.An(l), .B(m), .C(k), .Y(ori_ori_n70_));
  NAi21      o0042(.An(e), .B(h), .Y(ori_ori_n71_));
  NAi41      o0043(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n72_));
  INV        o0044(.A(m), .Y(ori_ori_n73_));
  NOi21      o0045(.An(k), .B(l), .Y(ori_ori_n74_));
  NA2        o0046(.A(ori_ori_n74_), .B(ori_ori_n73_), .Y(ori_ori_n75_));
  AN4        o0047(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n76_));
  NOi31      o0048(.An(h), .B(o), .C(f), .Y(ori_ori_n77_));
  NA2        o0049(.A(ori_ori_n77_), .B(ori_ori_n76_), .Y(ori_ori_n78_));
  NAi32      o0050(.An(m), .Bn(k), .C(j), .Y(ori_ori_n79_));
  NOi32      o0051(.An(h), .Bn(o), .C(f), .Y(ori_ori_n80_));
  NA2        o0052(.A(ori_ori_n80_), .B(ori_ori_n76_), .Y(ori_ori_n81_));
  OA220      o0053(.A0(ori_ori_n81_), .A1(ori_ori_n79_), .B0(ori_ori_n78_), .B1(ori_ori_n75_), .Y(ori_ori_n82_));
  NA2        o0054(.A(ori_ori_n82_), .B(ori_ori_n64_), .Y(ori_ori_n83_));
  INV        o0055(.A(n), .Y(ori_ori_n84_));
  NOi32      o0056(.An(e), .Bn(b), .C(d), .Y(ori_ori_n85_));
  NA2        o0057(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n86_));
  INV        o0058(.A(j), .Y(ori_ori_n87_));
  AN3        o0059(.A(m), .B(k), .C(i), .Y(ori_ori_n88_));
  NA3        o0060(.A(ori_ori_n88_), .B(ori_ori_n87_), .C(o), .Y(ori_ori_n89_));
  NO2        o0061(.A(ori_ori_n89_), .B(f), .Y(ori_ori_n90_));
  NAi32      o0062(.An(o), .Bn(f), .C(h), .Y(ori_ori_n91_));
  NAi31      o0063(.An(j), .B(m), .C(l), .Y(ori_ori_n92_));
  NO2        o0064(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  NA2        o0065(.A(m), .B(l), .Y(ori_ori_n94_));
  NAi31      o0066(.An(k), .B(j), .C(o), .Y(ori_ori_n95_));
  NO3        o0067(.A(ori_ori_n95_), .B(ori_ori_n94_), .C(f), .Y(ori_ori_n96_));
  AN2        o0068(.A(j), .B(o), .Y(ori_ori_n97_));
  NOi32      o0069(.An(m), .Bn(l), .C(i), .Y(ori_ori_n98_));
  NOi21      o0070(.An(o), .B(i), .Y(ori_ori_n99_));
  NOi32      o0071(.An(m), .Bn(j), .C(k), .Y(ori_ori_n100_));
  AOI220     o0072(.A0(ori_ori_n100_), .A1(ori_ori_n99_), .B0(ori_ori_n98_), .B1(ori_ori_n97_), .Y(ori_ori_n101_));
  NO3        o0073(.A(ori_ori_n96_), .B(ori_ori_n93_), .C(ori_ori_n90_), .Y(ori_ori_n102_));
  NAi41      o0074(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n103_));
  AN2        o0075(.A(e), .B(b), .Y(ori_ori_n104_));
  NOi31      o0076(.An(c), .B(h), .C(f), .Y(ori_ori_n105_));
  NA2        o0077(.A(ori_ori_n105_), .B(ori_ori_n104_), .Y(ori_ori_n106_));
  NO2        o0078(.A(ori_ori_n106_), .B(ori_ori_n103_), .Y(ori_ori_n107_));
  NOi21      o0079(.An(o), .B(f), .Y(ori_ori_n108_));
  NOi21      o0080(.An(i), .B(h), .Y(ori_ori_n109_));
  INV        o0081(.A(a), .Y(ori_ori_n110_));
  NA2        o0082(.A(ori_ori_n104_), .B(ori_ori_n110_), .Y(ori_ori_n111_));
  INV        o0083(.A(l), .Y(ori_ori_n112_));
  NOi21      o0084(.An(m), .B(n), .Y(ori_ori_n113_));
  AN2        o0085(.A(k), .B(h), .Y(ori_ori_n114_));
  INV        o0086(.A(b), .Y(ori_ori_n115_));
  NA2        o0087(.A(l), .B(j), .Y(ori_ori_n116_));
  AN2        o0088(.A(k), .B(i), .Y(ori_ori_n117_));
  NA2        o0089(.A(ori_ori_n117_), .B(ori_ori_n116_), .Y(ori_ori_n118_));
  NA2        o0090(.A(o), .B(e), .Y(ori_ori_n119_));
  NOi32      o0091(.An(c), .Bn(a), .C(d), .Y(ori_ori_n120_));
  NA2        o0092(.A(ori_ori_n120_), .B(ori_ori_n113_), .Y(ori_ori_n121_));
  INV        o0093(.A(ori_ori_n107_), .Y(ori_ori_n122_));
  OAI210     o0094(.A0(ori_ori_n102_), .A1(ori_ori_n86_), .B0(ori_ori_n122_), .Y(ori_ori_n123_));
  NOi31      o0095(.An(k), .B(m), .C(j), .Y(ori_ori_n124_));
  NA3        o0096(.A(ori_ori_n124_), .B(ori_ori_n77_), .C(ori_ori_n76_), .Y(ori_ori_n125_));
  NOi31      o0097(.An(k), .B(m), .C(i), .Y(ori_ori_n126_));
  NA3        o0098(.A(ori_ori_n126_), .B(ori_ori_n80_), .C(ori_ori_n76_), .Y(ori_ori_n127_));
  NA2        o0099(.A(ori_ori_n127_), .B(ori_ori_n125_), .Y(ori_ori_n128_));
  NOi32      o0100(.An(f), .Bn(b), .C(e), .Y(ori_ori_n129_));
  NAi21      o0101(.An(o), .B(h), .Y(ori_ori_n130_));
  NAi21      o0102(.An(m), .B(n), .Y(ori_ori_n131_));
  NAi21      o0103(.An(j), .B(k), .Y(ori_ori_n132_));
  NO3        o0104(.A(ori_ori_n132_), .B(ori_ori_n131_), .C(ori_ori_n130_), .Y(ori_ori_n133_));
  NAi41      o0105(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n134_));
  NAi31      o0106(.An(j), .B(k), .C(h), .Y(ori_ori_n135_));
  NO3        o0107(.A(ori_ori_n135_), .B(ori_ori_n134_), .C(ori_ori_n131_), .Y(ori_ori_n136_));
  AOI210     o0108(.A0(ori_ori_n133_), .A1(ori_ori_n129_), .B0(ori_ori_n136_), .Y(ori_ori_n137_));
  NO2        o0109(.A(k), .B(j), .Y(ori_ori_n138_));
  NO2        o0110(.A(ori_ori_n138_), .B(ori_ori_n131_), .Y(ori_ori_n139_));
  AN2        o0111(.A(k), .B(j), .Y(ori_ori_n140_));
  NAi21      o0112(.An(c), .B(b), .Y(ori_ori_n141_));
  NA2        o0113(.A(f), .B(d), .Y(ori_ori_n142_));
  NO4        o0114(.A(ori_ori_n142_), .B(ori_ori_n141_), .C(ori_ori_n140_), .D(ori_ori_n130_), .Y(ori_ori_n143_));
  NA2        o0115(.A(h), .B(c), .Y(ori_ori_n144_));
  NAi31      o0116(.An(f), .B(e), .C(b), .Y(ori_ori_n145_));
  NA2        o0117(.A(ori_ori_n143_), .B(ori_ori_n139_), .Y(ori_ori_n146_));
  NA2        o0118(.A(d), .B(b), .Y(ori_ori_n147_));
  NAi21      o0119(.An(e), .B(f), .Y(ori_ori_n148_));
  NO2        o0120(.A(ori_ori_n148_), .B(ori_ori_n147_), .Y(ori_ori_n149_));
  NA2        o0121(.A(b), .B(a), .Y(ori_ori_n150_));
  NAi21      o0122(.An(e), .B(o), .Y(ori_ori_n151_));
  NAi21      o0123(.An(c), .B(d), .Y(ori_ori_n152_));
  NAi31      o0124(.An(l), .B(k), .C(h), .Y(ori_ori_n153_));
  NO2        o0125(.A(ori_ori_n131_), .B(ori_ori_n153_), .Y(ori_ori_n154_));
  NA2        o0126(.A(ori_ori_n154_), .B(ori_ori_n149_), .Y(ori_ori_n155_));
  NAi41      o0127(.An(ori_ori_n128_), .B(ori_ori_n155_), .C(ori_ori_n146_), .D(ori_ori_n137_), .Y(ori_ori_n156_));
  NAi31      o0128(.An(e), .B(f), .C(b), .Y(ori_ori_n157_));
  NOi21      o0129(.An(o), .B(d), .Y(ori_ori_n158_));
  NO2        o0130(.A(ori_ori_n158_), .B(ori_ori_n157_), .Y(ori_ori_n159_));
  NOi21      o0131(.An(h), .B(i), .Y(ori_ori_n160_));
  NOi21      o0132(.An(k), .B(m), .Y(ori_ori_n161_));
  NA3        o0133(.A(ori_ori_n161_), .B(ori_ori_n160_), .C(n), .Y(ori_ori_n162_));
  NOi21      o0134(.An(ori_ori_n159_), .B(ori_ori_n162_), .Y(ori_ori_n163_));
  NOi21      o0135(.An(h), .B(o), .Y(ori_ori_n164_));
  NO2        o0136(.A(ori_ori_n142_), .B(ori_ori_n141_), .Y(ori_ori_n165_));
  NAi31      o0137(.An(l), .B(j), .C(h), .Y(ori_ori_n166_));
  NO2        o0138(.A(ori_ori_n166_), .B(ori_ori_n49_), .Y(ori_ori_n167_));
  NA2        o0139(.A(ori_ori_n167_), .B(ori_ori_n67_), .Y(ori_ori_n168_));
  NOi32      o0140(.An(n), .Bn(k), .C(m), .Y(ori_ori_n169_));
  NA2        o0141(.A(l), .B(i), .Y(ori_ori_n170_));
  INV        o0142(.A(ori_ori_n168_), .Y(ori_ori_n171_));
  NAi31      o0143(.An(d), .B(f), .C(c), .Y(ori_ori_n172_));
  NAi31      o0144(.An(e), .B(f), .C(c), .Y(ori_ori_n173_));
  NA2        o0145(.A(ori_ori_n173_), .B(ori_ori_n172_), .Y(ori_ori_n174_));
  NA2        o0146(.A(j), .B(h), .Y(ori_ori_n175_));
  OR3        o0147(.A(n), .B(m), .C(k), .Y(ori_ori_n176_));
  NO2        o0148(.A(ori_ori_n176_), .B(ori_ori_n175_), .Y(ori_ori_n177_));
  NAi32      o0149(.An(m), .Bn(k), .C(n), .Y(ori_ori_n178_));
  NO2        o0150(.A(ori_ori_n178_), .B(ori_ori_n175_), .Y(ori_ori_n179_));
  AOI220     o0151(.A0(ori_ori_n179_), .A1(ori_ori_n159_), .B0(ori_ori_n177_), .B1(ori_ori_n174_), .Y(ori_ori_n180_));
  NO2        o0152(.A(n), .B(m), .Y(ori_ori_n181_));
  NA2        o0153(.A(ori_ori_n181_), .B(ori_ori_n50_), .Y(ori_ori_n182_));
  NAi21      o0154(.An(f), .B(e), .Y(ori_ori_n183_));
  NA2        o0155(.A(d), .B(c), .Y(ori_ori_n184_));
  NO2        o0156(.A(ori_ori_n184_), .B(ori_ori_n183_), .Y(ori_ori_n185_));
  NOi21      o0157(.An(ori_ori_n185_), .B(ori_ori_n182_), .Y(ori_ori_n186_));
  NAi31      o0158(.An(m), .B(n), .C(b), .Y(ori_ori_n187_));
  NA2        o0159(.A(k), .B(i), .Y(ori_ori_n188_));
  NAi21      o0160(.An(h), .B(f), .Y(ori_ori_n189_));
  NO2        o0161(.A(ori_ori_n189_), .B(ori_ori_n188_), .Y(ori_ori_n190_));
  NO2        o0162(.A(ori_ori_n187_), .B(ori_ori_n152_), .Y(ori_ori_n191_));
  NA2        o0163(.A(ori_ori_n191_), .B(ori_ori_n190_), .Y(ori_ori_n192_));
  NOi32      o0164(.An(f), .Bn(c), .C(d), .Y(ori_ori_n193_));
  NOi32      o0165(.An(f), .Bn(c), .C(e), .Y(ori_ori_n194_));
  NO2        o0166(.A(ori_ori_n194_), .B(ori_ori_n193_), .Y(ori_ori_n195_));
  NO3        o0167(.A(n), .B(m), .C(j), .Y(ori_ori_n196_));
  NA2        o0168(.A(ori_ori_n196_), .B(ori_ori_n114_), .Y(ori_ori_n197_));
  AO210      o0169(.A0(ori_ori_n197_), .A1(ori_ori_n182_), .B0(ori_ori_n195_), .Y(ori_ori_n198_));
  NAi41      o0170(.An(ori_ori_n186_), .B(ori_ori_n198_), .C(ori_ori_n192_), .D(ori_ori_n180_), .Y(ori_ori_n199_));
  OR4        o0171(.A(ori_ori_n199_), .B(ori_ori_n171_), .C(ori_ori_n163_), .D(ori_ori_n156_), .Y(ori_ori_n200_));
  NO4        o0172(.A(ori_ori_n200_), .B(ori_ori_n123_), .C(ori_ori_n83_), .D(ori_ori_n55_), .Y(ori_ori_n201_));
  NA3        o0173(.A(m), .B(ori_ori_n112_), .C(j), .Y(ori_ori_n202_));
  NAi31      o0174(.An(n), .B(h), .C(o), .Y(ori_ori_n203_));
  NO2        o0175(.A(ori_ori_n203_), .B(ori_ori_n202_), .Y(ori_ori_n204_));
  NOi32      o0176(.An(m), .Bn(k), .C(l), .Y(ori_ori_n205_));
  NA3        o0177(.A(ori_ori_n205_), .B(ori_ori_n87_), .C(o), .Y(ori_ori_n206_));
  NO2        o0178(.A(ori_ori_n206_), .B(n), .Y(ori_ori_n207_));
  NOi21      o0179(.An(k), .B(j), .Y(ori_ori_n208_));
  NA4        o0180(.A(ori_ori_n208_), .B(ori_ori_n113_), .C(i), .D(o), .Y(ori_ori_n209_));
  AN2        o0181(.A(i), .B(o), .Y(ori_ori_n210_));
  NA3        o0182(.A(ori_ori_n74_), .B(ori_ori_n210_), .C(ori_ori_n113_), .Y(ori_ori_n211_));
  NA2        o0183(.A(ori_ori_n211_), .B(ori_ori_n209_), .Y(ori_ori_n212_));
  NO3        o0184(.A(ori_ori_n212_), .B(ori_ori_n207_), .C(ori_ori_n204_), .Y(ori_ori_n213_));
  NAi41      o0185(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n214_));
  INV        o0186(.A(ori_ori_n214_), .Y(ori_ori_n215_));
  INV        o0187(.A(f), .Y(ori_ori_n216_));
  INV        o0188(.A(o), .Y(ori_ori_n217_));
  NOi31      o0189(.An(i), .B(j), .C(h), .Y(ori_ori_n218_));
  NOi21      o0190(.An(l), .B(m), .Y(ori_ori_n219_));
  NA2        o0191(.A(ori_ori_n219_), .B(ori_ori_n218_), .Y(ori_ori_n220_));
  NO3        o0192(.A(ori_ori_n220_), .B(ori_ori_n217_), .C(ori_ori_n216_), .Y(ori_ori_n221_));
  NA2        o0193(.A(ori_ori_n221_), .B(ori_ori_n215_), .Y(ori_ori_n222_));
  OAI210     o0194(.A0(ori_ori_n213_), .A1(ori_ori_n32_), .B0(ori_ori_n222_), .Y(ori_ori_n223_));
  NOi21      o0195(.An(n), .B(m), .Y(ori_ori_n224_));
  NOi32      o0196(.An(l), .Bn(i), .C(j), .Y(ori_ori_n225_));
  NA2        o0197(.A(ori_ori_n225_), .B(ori_ori_n224_), .Y(ori_ori_n226_));
  OA220      o0198(.A0(ori_ori_n226_), .A1(ori_ori_n106_), .B0(ori_ori_n79_), .B1(ori_ori_n78_), .Y(ori_ori_n227_));
  NAi21      o0199(.An(j), .B(h), .Y(ori_ori_n228_));
  XN2        o0200(.A(i), .B(h), .Y(ori_ori_n229_));
  NA2        o0201(.A(ori_ori_n229_), .B(ori_ori_n228_), .Y(ori_ori_n230_));
  NOi31      o0202(.An(k), .B(n), .C(m), .Y(ori_ori_n231_));
  NOi31      o0203(.An(ori_ori_n231_), .B(ori_ori_n184_), .C(ori_ori_n183_), .Y(ori_ori_n232_));
  NA2        o0204(.A(ori_ori_n232_), .B(ori_ori_n230_), .Y(ori_ori_n233_));
  NAi31      o0205(.An(f), .B(e), .C(c), .Y(ori_ori_n234_));
  NO4        o0206(.A(ori_ori_n234_), .B(ori_ori_n176_), .C(ori_ori_n175_), .D(ori_ori_n59_), .Y(ori_ori_n235_));
  NA4        o0207(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n236_));
  NAi32      o0208(.An(m), .Bn(i), .C(k), .Y(ori_ori_n237_));
  NO3        o0209(.A(ori_ori_n237_), .B(ori_ori_n91_), .C(ori_ori_n236_), .Y(ori_ori_n238_));
  INV        o0210(.A(k), .Y(ori_ori_n239_));
  NO2        o0211(.A(ori_ori_n238_), .B(ori_ori_n235_), .Y(ori_ori_n240_));
  NAi21      o0212(.An(n), .B(a), .Y(ori_ori_n241_));
  NO2        o0213(.A(ori_ori_n241_), .B(ori_ori_n147_), .Y(ori_ori_n242_));
  NAi41      o0214(.An(o), .B(m), .C(k), .D(h), .Y(ori_ori_n243_));
  NO2        o0215(.A(ori_ori_n243_), .B(e), .Y(ori_ori_n244_));
  NA2        o0216(.A(ori_ori_n244_), .B(ori_ori_n242_), .Y(ori_ori_n245_));
  AN4        o0217(.A(ori_ori_n245_), .B(ori_ori_n240_), .C(ori_ori_n233_), .D(ori_ori_n227_), .Y(ori_ori_n246_));
  OR2        o0218(.A(h), .B(o), .Y(ori_ori_n247_));
  NO2        o0219(.A(ori_ori_n247_), .B(ori_ori_n103_), .Y(ori_ori_n248_));
  NA2        o0220(.A(ori_ori_n248_), .B(ori_ori_n129_), .Y(ori_ori_n249_));
  NAi41      o0221(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n250_));
  NO2        o0222(.A(ori_ori_n250_), .B(ori_ori_n216_), .Y(ori_ori_n251_));
  NA2        o0223(.A(ori_ori_n161_), .B(ori_ori_n109_), .Y(ori_ori_n252_));
  NAi21      o0224(.An(ori_ori_n252_), .B(ori_ori_n251_), .Y(ori_ori_n253_));
  NO2        o0225(.A(n), .B(a), .Y(ori_ori_n254_));
  NAi31      o0226(.An(ori_ori_n243_), .B(ori_ori_n254_), .C(ori_ori_n104_), .Y(ori_ori_n255_));
  AN2        o0227(.A(ori_ori_n255_), .B(ori_ori_n253_), .Y(ori_ori_n256_));
  NAi21      o0228(.An(h), .B(i), .Y(ori_ori_n257_));
  NA2        o0229(.A(ori_ori_n181_), .B(k), .Y(ori_ori_n258_));
  NO2        o0230(.A(ori_ori_n258_), .B(ori_ori_n257_), .Y(ori_ori_n259_));
  NA2        o0231(.A(ori_ori_n259_), .B(ori_ori_n193_), .Y(ori_ori_n260_));
  NA3        o0232(.A(ori_ori_n260_), .B(ori_ori_n256_), .C(ori_ori_n249_), .Y(ori_ori_n261_));
  NOi21      o0233(.An(o), .B(e), .Y(ori_ori_n262_));
  NO2        o0234(.A(ori_ori_n72_), .B(ori_ori_n73_), .Y(ori_ori_n263_));
  NA2        o0235(.A(ori_ori_n263_), .B(ori_ori_n262_), .Y(ori_ori_n264_));
  NOi32      o0236(.An(l), .Bn(j), .C(i), .Y(ori_ori_n265_));
  AOI210     o0237(.A0(ori_ori_n74_), .A1(ori_ori_n87_), .B0(ori_ori_n265_), .Y(ori_ori_n266_));
  NAi21      o0238(.An(f), .B(o), .Y(ori_ori_n267_));
  NO2        o0239(.A(ori_ori_n267_), .B(ori_ori_n65_), .Y(ori_ori_n268_));
  NO2        o0240(.A(ori_ori_n69_), .B(ori_ori_n116_), .Y(ori_ori_n269_));
  NO2        o0241(.A(ori_ori_n266_), .B(ori_ori_n264_), .Y(ori_ori_n270_));
  NO2        o0242(.A(ori_ori_n132_), .B(ori_ori_n49_), .Y(ori_ori_n271_));
  NOi41      o0243(.An(ori_ori_n246_), .B(ori_ori_n270_), .C(ori_ori_n261_), .D(ori_ori_n223_), .Y(ori_ori_n272_));
  NO4        o0244(.A(ori_ori_n204_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n273_));
  NO2        o0245(.A(ori_ori_n273_), .B(ori_ori_n111_), .Y(ori_ori_n274_));
  NA3        o0246(.A(ori_ori_n59_), .B(c), .C(b), .Y(ori_ori_n275_));
  NAi21      o0247(.An(h), .B(o), .Y(ori_ori_n276_));
  OR4        o0248(.A(ori_ori_n276_), .B(ori_ori_n275_), .C(ori_ori_n226_), .D(e), .Y(ori_ori_n277_));
  NO2        o0249(.A(ori_ori_n252_), .B(ori_ori_n267_), .Y(ori_ori_n278_));
  NAi31      o0250(.An(o), .B(k), .C(h), .Y(ori_ori_n279_));
  NAi31      o0251(.An(e), .B(d), .C(a), .Y(ori_ori_n280_));
  INV        o0252(.A(ori_ori_n277_), .Y(ori_ori_n281_));
  NA4        o0253(.A(ori_ori_n161_), .B(ori_ori_n80_), .C(ori_ori_n76_), .D(ori_ori_n116_), .Y(ori_ori_n282_));
  NA3        o0254(.A(ori_ori_n161_), .B(ori_ori_n160_), .C(ori_ori_n84_), .Y(ori_ori_n283_));
  NO2        o0255(.A(ori_ori_n283_), .B(ori_ori_n195_), .Y(ori_ori_n284_));
  NOi21      o0256(.An(ori_ori_n282_), .B(ori_ori_n284_), .Y(ori_ori_n285_));
  NA3        o0257(.A(e), .B(c), .C(b), .Y(ori_ori_n286_));
  NO2        o0258(.A(ori_ori_n60_), .B(ori_ori_n286_), .Y(ori_ori_n287_));
  NAi32      o0259(.An(k), .Bn(i), .C(j), .Y(ori_ori_n288_));
  NAi31      o0260(.An(h), .B(l), .C(i), .Y(ori_ori_n289_));
  NA3        o0261(.A(ori_ori_n289_), .B(ori_ori_n288_), .C(ori_ori_n166_), .Y(ori_ori_n290_));
  NOi21      o0262(.An(ori_ori_n290_), .B(ori_ori_n49_), .Y(ori_ori_n291_));
  OAI210     o0263(.A0(ori_ori_n268_), .A1(ori_ori_n287_), .B0(ori_ori_n291_), .Y(ori_ori_n292_));
  NAi21      o0264(.An(l), .B(k), .Y(ori_ori_n293_));
  NO2        o0265(.A(ori_ori_n293_), .B(ori_ori_n49_), .Y(ori_ori_n294_));
  NOi21      o0266(.An(l), .B(j), .Y(ori_ori_n295_));
  NA2        o0267(.A(ori_ori_n164_), .B(ori_ori_n295_), .Y(ori_ori_n296_));
  NA3        o0268(.A(ori_ori_n117_), .B(ori_ori_n116_), .C(o), .Y(ori_ori_n297_));
  OR3        o0269(.A(ori_ori_n72_), .B(ori_ori_n73_), .C(e), .Y(ori_ori_n298_));
  AOI210     o0270(.A0(ori_ori_n297_), .A1(ori_ori_n296_), .B0(ori_ori_n298_), .Y(ori_ori_n299_));
  INV        o0271(.A(ori_ori_n299_), .Y(ori_ori_n300_));
  NAi32      o0272(.An(j), .Bn(h), .C(i), .Y(ori_ori_n301_));
  NAi21      o0273(.An(m), .B(l), .Y(ori_ori_n302_));
  NO3        o0274(.A(ori_ori_n302_), .B(ori_ori_n301_), .C(ori_ori_n84_), .Y(ori_ori_n303_));
  NA2        o0275(.A(h), .B(o), .Y(ori_ori_n304_));
  NA2        o0276(.A(ori_ori_n169_), .B(ori_ori_n45_), .Y(ori_ori_n305_));
  NO2        o0277(.A(ori_ori_n305_), .B(ori_ori_n304_), .Y(ori_ori_n306_));
  NA2        o0278(.A(ori_ori_n306_), .B(ori_ori_n165_), .Y(ori_ori_n307_));
  NA4        o0279(.A(ori_ori_n307_), .B(ori_ori_n300_), .C(ori_ori_n292_), .D(ori_ori_n285_), .Y(ori_ori_n308_));
  NO2        o0280(.A(ori_ori_n145_), .B(d), .Y(ori_ori_n309_));
  NA2        o0281(.A(ori_ori_n309_), .B(ori_ori_n53_), .Y(ori_ori_n310_));
  NO2        o0282(.A(ori_ori_n106_), .B(ori_ori_n103_), .Y(ori_ori_n311_));
  NAi32      o0283(.An(n), .Bn(m), .C(l), .Y(ori_ori_n312_));
  NO2        o0284(.A(ori_ori_n312_), .B(ori_ori_n301_), .Y(ori_ori_n313_));
  NA2        o0285(.A(ori_ori_n313_), .B(ori_ori_n185_), .Y(ori_ori_n314_));
  NO2        o0286(.A(ori_ori_n121_), .B(ori_ori_n115_), .Y(ori_ori_n315_));
  NAi31      o0287(.An(k), .B(l), .C(j), .Y(ori_ori_n316_));
  OAI210     o0288(.A0(ori_ori_n293_), .A1(j), .B0(ori_ori_n316_), .Y(ori_ori_n317_));
  NOi21      o0289(.An(ori_ori_n317_), .B(ori_ori_n119_), .Y(ori_ori_n318_));
  NA2        o0290(.A(ori_ori_n318_), .B(ori_ori_n315_), .Y(ori_ori_n319_));
  NA3        o0291(.A(ori_ori_n319_), .B(ori_ori_n314_), .C(ori_ori_n310_), .Y(ori_ori_n320_));
  NO4        o0292(.A(ori_ori_n320_), .B(ori_ori_n308_), .C(ori_ori_n281_), .D(ori_ori_n274_), .Y(ori_ori_n321_));
  NA2        o0293(.A(ori_ori_n259_), .B(ori_ori_n194_), .Y(ori_ori_n322_));
  NAi21      o0294(.An(m), .B(k), .Y(ori_ori_n323_));
  NO2        o0295(.A(ori_ori_n229_), .B(ori_ori_n323_), .Y(ori_ori_n324_));
  NAi41      o0296(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n325_));
  NO2        o0297(.A(ori_ori_n325_), .B(ori_ori_n151_), .Y(ori_ori_n326_));
  NA2        o0298(.A(ori_ori_n326_), .B(ori_ori_n324_), .Y(ori_ori_n327_));
  NAi31      o0299(.An(i), .B(l), .C(h), .Y(ori_ori_n328_));
  NO4        o0300(.A(ori_ori_n328_), .B(ori_ori_n151_), .C(ori_ori_n72_), .D(ori_ori_n73_), .Y(ori_ori_n329_));
  NA2        o0301(.A(e), .B(c), .Y(ori_ori_n330_));
  NO3        o0302(.A(ori_ori_n330_), .B(n), .C(d), .Y(ori_ori_n331_));
  NOi21      o0303(.An(f), .B(h), .Y(ori_ori_n332_));
  NA2        o0304(.A(ori_ori_n332_), .B(ori_ori_n117_), .Y(ori_ori_n333_));
  NO2        o0305(.A(ori_ori_n333_), .B(ori_ori_n217_), .Y(ori_ori_n334_));
  NAi31      o0306(.An(d), .B(e), .C(b), .Y(ori_ori_n335_));
  NO2        o0307(.A(ori_ori_n131_), .B(ori_ori_n335_), .Y(ori_ori_n336_));
  NA2        o0308(.A(ori_ori_n336_), .B(ori_ori_n334_), .Y(ori_ori_n337_));
  NAi41      o0309(.An(ori_ori_n329_), .B(ori_ori_n337_), .C(ori_ori_n327_), .D(ori_ori_n322_), .Y(ori_ori_n338_));
  NO4        o0310(.A(ori_ori_n325_), .B(ori_ori_n79_), .C(ori_ori_n71_), .D(ori_ori_n217_), .Y(ori_ori_n339_));
  NA2        o0311(.A(ori_ori_n254_), .B(ori_ori_n104_), .Y(ori_ori_n340_));
  OR2        o0312(.A(ori_ori_n340_), .B(ori_ori_n206_), .Y(ori_ori_n341_));
  NOi31      o0313(.An(l), .B(n), .C(m), .Y(ori_ori_n342_));
  NA2        o0314(.A(ori_ori_n342_), .B(ori_ori_n218_), .Y(ori_ori_n343_));
  NO2        o0315(.A(ori_ori_n343_), .B(ori_ori_n195_), .Y(ori_ori_n344_));
  NAi32      o0316(.An(ori_ori_n344_), .Bn(ori_ori_n339_), .C(ori_ori_n341_), .Y(ori_ori_n345_));
  NAi32      o0317(.An(m), .Bn(j), .C(k), .Y(ori_ori_n346_));
  NAi41      o0318(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n347_));
  OAI210     o0319(.A0(ori_ori_n214_), .A1(ori_ori_n346_), .B0(ori_ori_n347_), .Y(ori_ori_n348_));
  NOi31      o0320(.An(j), .B(m), .C(k), .Y(ori_ori_n349_));
  NO2        o0321(.A(ori_ori_n124_), .B(ori_ori_n349_), .Y(ori_ori_n350_));
  AN3        o0322(.A(h), .B(o), .C(f), .Y(ori_ori_n351_));
  NAi31      o0323(.An(ori_ori_n350_), .B(ori_ori_n351_), .C(ori_ori_n348_), .Y(ori_ori_n352_));
  NOi32      o0324(.An(m), .Bn(j), .C(l), .Y(ori_ori_n353_));
  NO2        o0325(.A(ori_ori_n353_), .B(ori_ori_n98_), .Y(ori_ori_n354_));
  NAi32      o0326(.An(ori_ori_n354_), .Bn(ori_ori_n203_), .C(ori_ori_n309_), .Y(ori_ori_n355_));
  NO2        o0327(.A(ori_ori_n302_), .B(ori_ori_n301_), .Y(ori_ori_n356_));
  NO2        o0328(.A(ori_ori_n220_), .B(o), .Y(ori_ori_n357_));
  NO2        o0329(.A(ori_ori_n157_), .B(ori_ori_n84_), .Y(ori_ori_n358_));
  AOI220     o0330(.A0(ori_ori_n358_), .A1(ori_ori_n357_), .B0(ori_ori_n251_), .B1(ori_ori_n356_), .Y(ori_ori_n359_));
  NA2        o0331(.A(ori_ori_n237_), .B(ori_ori_n79_), .Y(ori_ori_n360_));
  NA3        o0332(.A(ori_ori_n360_), .B(ori_ori_n351_), .C(ori_ori_n215_), .Y(ori_ori_n361_));
  NA4        o0333(.A(ori_ori_n361_), .B(ori_ori_n359_), .C(ori_ori_n355_), .D(ori_ori_n352_), .Y(ori_ori_n362_));
  NA3        o0334(.A(h), .B(o), .C(f), .Y(ori_ori_n363_));
  NO2        o0335(.A(ori_ori_n363_), .B(ori_ori_n75_), .Y(ori_ori_n364_));
  INV        o0336(.A(ori_ori_n214_), .Y(ori_ori_n365_));
  NA2        o0337(.A(ori_ori_n164_), .B(e), .Y(ori_ori_n366_));
  NO2        o0338(.A(ori_ori_n366_), .B(ori_ori_n41_), .Y(ori_ori_n367_));
  AOI220     o0339(.A0(ori_ori_n367_), .A1(ori_ori_n315_), .B0(ori_ori_n365_), .B1(ori_ori_n364_), .Y(ori_ori_n368_));
  NOi32      o0340(.An(j), .Bn(o), .C(i), .Y(ori_ori_n369_));
  NA3        o0341(.A(ori_ori_n369_), .B(ori_ori_n293_), .C(ori_ori_n113_), .Y(ori_ori_n370_));
  AO210      o0342(.A0(ori_ori_n111_), .A1(ori_ori_n32_), .B0(ori_ori_n370_), .Y(ori_ori_n371_));
  NOi32      o0343(.An(e), .Bn(b), .C(a), .Y(ori_ori_n372_));
  AN2        o0344(.A(l), .B(j), .Y(ori_ori_n373_));
  NO2        o0345(.A(ori_ori_n323_), .B(ori_ori_n373_), .Y(ori_ori_n374_));
  NO3        o0346(.A(ori_ori_n325_), .B(ori_ori_n71_), .C(ori_ori_n217_), .Y(ori_ori_n375_));
  NA3        o0347(.A(ori_ori_n211_), .B(ori_ori_n209_), .C(ori_ori_n35_), .Y(ori_ori_n376_));
  AOI220     o0348(.A0(ori_ori_n376_), .A1(ori_ori_n372_), .B0(ori_ori_n375_), .B1(ori_ori_n374_), .Y(ori_ori_n377_));
  NO2        o0349(.A(ori_ori_n335_), .B(n), .Y(ori_ori_n378_));
  NA2        o0350(.A(ori_ori_n210_), .B(k), .Y(ori_ori_n379_));
  NA3        o0351(.A(m), .B(ori_ori_n112_), .C(ori_ori_n216_), .Y(ori_ori_n380_));
  NA4        o0352(.A(ori_ori_n205_), .B(ori_ori_n87_), .C(o), .D(ori_ori_n216_), .Y(ori_ori_n381_));
  OAI210     o0353(.A0(ori_ori_n380_), .A1(ori_ori_n379_), .B0(ori_ori_n381_), .Y(ori_ori_n382_));
  NAi41      o0354(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n383_));
  NA2        o0355(.A(ori_ori_n51_), .B(ori_ori_n113_), .Y(ori_ori_n384_));
  NO2        o0356(.A(ori_ori_n384_), .B(ori_ori_n383_), .Y(ori_ori_n385_));
  AOI220     o0357(.A0(ori_ori_n385_), .A1(b), .B0(ori_ori_n382_), .B1(ori_ori_n378_), .Y(ori_ori_n386_));
  NA4        o0358(.A(ori_ori_n386_), .B(ori_ori_n377_), .C(ori_ori_n371_), .D(ori_ori_n368_), .Y(ori_ori_n387_));
  NO4        o0359(.A(ori_ori_n387_), .B(ori_ori_n362_), .C(ori_ori_n345_), .D(ori_ori_n338_), .Y(ori_ori_n388_));
  NA4        o0360(.A(ori_ori_n388_), .B(ori_ori_n321_), .C(ori_ori_n272_), .D(ori_ori_n201_), .Y(ori10));
  NA3        o0361(.A(m), .B(k), .C(i), .Y(ori_ori_n390_));
  NO3        o0362(.A(ori_ori_n390_), .B(j), .C(ori_ori_n217_), .Y(ori_ori_n391_));
  NOi21      o0363(.An(e), .B(f), .Y(ori_ori_n392_));
  NO4        o0364(.A(ori_ori_n152_), .B(ori_ori_n392_), .C(n), .D(ori_ori_n110_), .Y(ori_ori_n393_));
  NAi31      o0365(.An(b), .B(f), .C(c), .Y(ori_ori_n394_));
  INV        o0366(.A(ori_ori_n394_), .Y(ori_ori_n395_));
  NOi32      o0367(.An(k), .Bn(h), .C(j), .Y(ori_ori_n396_));
  NA2        o0368(.A(ori_ori_n396_), .B(ori_ori_n224_), .Y(ori_ori_n397_));
  NA2        o0369(.A(ori_ori_n162_), .B(ori_ori_n397_), .Y(ori_ori_n398_));
  AOI220     o0370(.A0(ori_ori_n398_), .A1(ori_ori_n395_), .B0(ori_ori_n393_), .B1(ori_ori_n391_), .Y(ori_ori_n399_));
  AN2        o0371(.A(j), .B(h), .Y(ori_ori_n400_));
  NO3        o0372(.A(n), .B(m), .C(k), .Y(ori_ori_n401_));
  NA2        o0373(.A(ori_ori_n401_), .B(ori_ori_n400_), .Y(ori_ori_n402_));
  NO3        o0374(.A(ori_ori_n402_), .B(ori_ori_n152_), .C(ori_ori_n216_), .Y(ori_ori_n403_));
  OR2        o0375(.A(m), .B(k), .Y(ori_ori_n404_));
  NO2        o0376(.A(ori_ori_n175_), .B(ori_ori_n404_), .Y(ori_ori_n405_));
  NA4        o0377(.A(n), .B(f), .C(c), .D(ori_ori_n115_), .Y(ori_ori_n406_));
  NOi21      o0378(.An(ori_ori_n405_), .B(ori_ori_n406_), .Y(ori_ori_n407_));
  NOi32      o0379(.An(d), .Bn(a), .C(c), .Y(ori_ori_n408_));
  NA2        o0380(.A(ori_ori_n408_), .B(ori_ori_n183_), .Y(ori_ori_n409_));
  NAi21      o0381(.An(i), .B(o), .Y(ori_ori_n410_));
  NAi31      o0382(.An(k), .B(m), .C(j), .Y(ori_ori_n411_));
  NO3        o0383(.A(ori_ori_n411_), .B(ori_ori_n410_), .C(n), .Y(ori_ori_n412_));
  NOi21      o0384(.An(ori_ori_n412_), .B(ori_ori_n409_), .Y(ori_ori_n413_));
  NO3        o0385(.A(ori_ori_n413_), .B(ori_ori_n407_), .C(ori_ori_n403_), .Y(ori_ori_n414_));
  NO2        o0386(.A(ori_ori_n406_), .B(ori_ori_n302_), .Y(ori_ori_n415_));
  NOi32      o0387(.An(f), .Bn(d), .C(c), .Y(ori_ori_n416_));
  AOI220     o0388(.A0(ori_ori_n416_), .A1(ori_ori_n313_), .B0(ori_ori_n415_), .B1(ori_ori_n218_), .Y(ori_ori_n417_));
  NA3        o0389(.A(ori_ori_n417_), .B(ori_ori_n414_), .C(ori_ori_n399_), .Y(ori_ori_n418_));
  NO2        o0390(.A(ori_ori_n59_), .B(ori_ori_n115_), .Y(ori_ori_n419_));
  NA2        o0391(.A(ori_ori_n254_), .B(ori_ori_n419_), .Y(ori_ori_n420_));
  INV        o0392(.A(e), .Y(ori_ori_n421_));
  NA2        o0393(.A(ori_ori_n46_), .B(e), .Y(ori_ori_n422_));
  OAI220     o0394(.A0(ori_ori_n422_), .A1(ori_ori_n202_), .B0(ori_ori_n206_), .B1(ori_ori_n421_), .Y(ori_ori_n423_));
  AN2        o0395(.A(o), .B(e), .Y(ori_ori_n424_));
  NA3        o0396(.A(ori_ori_n424_), .B(ori_ori_n205_), .C(i), .Y(ori_ori_n425_));
  OAI210     o0397(.A0(ori_ori_n89_), .A1(ori_ori_n421_), .B0(ori_ori_n425_), .Y(ori_ori_n426_));
  NO2        o0398(.A(ori_ori_n101_), .B(ori_ori_n421_), .Y(ori_ori_n427_));
  NO3        o0399(.A(ori_ori_n427_), .B(ori_ori_n426_), .C(ori_ori_n423_), .Y(ori_ori_n428_));
  NOi32      o0400(.An(h), .Bn(e), .C(o), .Y(ori_ori_n429_));
  NA3        o0401(.A(ori_ori_n429_), .B(ori_ori_n295_), .C(m), .Y(ori_ori_n430_));
  NOi21      o0402(.An(o), .B(h), .Y(ori_ori_n431_));
  AN3        o0403(.A(m), .B(l), .C(i), .Y(ori_ori_n432_));
  NA3        o0404(.A(ori_ori_n432_), .B(ori_ori_n431_), .C(e), .Y(ori_ori_n433_));
  AN3        o0405(.A(h), .B(o), .C(e), .Y(ori_ori_n434_));
  NA2        o0406(.A(ori_ori_n434_), .B(ori_ori_n98_), .Y(ori_ori_n435_));
  AN3        o0407(.A(ori_ori_n435_), .B(ori_ori_n433_), .C(ori_ori_n430_), .Y(ori_ori_n436_));
  AOI210     o0408(.A0(ori_ori_n436_), .A1(ori_ori_n428_), .B0(ori_ori_n420_), .Y(ori_ori_n437_));
  NA3        o0409(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(e), .Y(ori_ori_n438_));
  NO2        o0410(.A(ori_ori_n438_), .B(ori_ori_n420_), .Y(ori_ori_n439_));
  NAi31      o0411(.An(b), .B(c), .C(a), .Y(ori_ori_n440_));
  NO2        o0412(.A(ori_ori_n440_), .B(n), .Y(ori_ori_n441_));
  NA2        o0413(.A(ori_ori_n51_), .B(m), .Y(ori_ori_n442_));
  NO2        o0414(.A(ori_ori_n442_), .B(ori_ori_n148_), .Y(ori_ori_n443_));
  NA2        o0415(.A(ori_ori_n443_), .B(ori_ori_n441_), .Y(ori_ori_n444_));
  INV        o0416(.A(ori_ori_n444_), .Y(ori_ori_n445_));
  NO4        o0417(.A(ori_ori_n445_), .B(ori_ori_n439_), .C(ori_ori_n437_), .D(ori_ori_n418_), .Y(ori_ori_n446_));
  NA2        o0418(.A(i), .B(o), .Y(ori_ori_n447_));
  NO3        o0419(.A(ori_ori_n280_), .B(ori_ori_n447_), .C(c), .Y(ori_ori_n448_));
  NOi21      o0420(.An(d), .B(c), .Y(ori_ori_n449_));
  NA3        o0421(.A(i), .B(o), .C(f), .Y(ori_ori_n450_));
  OR2        o0422(.A(ori_ori_n450_), .B(ori_ori_n70_), .Y(ori_ori_n451_));
  NA2        o0423(.A(ori_ori_n448_), .B(ori_ori_n294_), .Y(ori_ori_n452_));
  OR2        o0424(.A(n), .B(m), .Y(ori_ori_n453_));
  NO2        o0425(.A(ori_ori_n453_), .B(ori_ori_n153_), .Y(ori_ori_n454_));
  NO2        o0426(.A(ori_ori_n184_), .B(ori_ori_n148_), .Y(ori_ori_n455_));
  OAI210     o0427(.A0(ori_ori_n454_), .A1(ori_ori_n177_), .B0(ori_ori_n455_), .Y(ori_ori_n456_));
  INV        o0428(.A(ori_ori_n384_), .Y(ori_ori_n457_));
  NA3        o0429(.A(ori_ori_n457_), .B(ori_ori_n372_), .C(d), .Y(ori_ori_n458_));
  NO2        o0430(.A(ori_ori_n440_), .B(ori_ori_n49_), .Y(ori_ori_n459_));
  NAi21      o0431(.An(k), .B(j), .Y(ori_ori_n460_));
  NAi21      o0432(.An(e), .B(d), .Y(ori_ori_n461_));
  INV        o0433(.A(ori_ori_n461_), .Y(ori_ori_n462_));
  NO2        o0434(.A(ori_ori_n258_), .B(ori_ori_n216_), .Y(ori_ori_n463_));
  NA3        o0435(.A(ori_ori_n463_), .B(ori_ori_n462_), .C(ori_ori_n230_), .Y(ori_ori_n464_));
  NA3        o0436(.A(ori_ori_n464_), .B(ori_ori_n458_), .C(ori_ori_n456_), .Y(ori_ori_n465_));
  NO2        o0437(.A(ori_ori_n343_), .B(ori_ori_n216_), .Y(ori_ori_n466_));
  NA2        o0438(.A(ori_ori_n466_), .B(ori_ori_n462_), .Y(ori_ori_n467_));
  NOi31      o0439(.An(n), .B(m), .C(k), .Y(ori_ori_n468_));
  AOI220     o0440(.A0(ori_ori_n468_), .A1(ori_ori_n400_), .B0(ori_ori_n224_), .B1(ori_ori_n50_), .Y(ori_ori_n469_));
  NAi31      o0441(.An(o), .B(f), .C(c), .Y(ori_ori_n470_));
  OR3        o0442(.A(ori_ori_n470_), .B(ori_ori_n469_), .C(e), .Y(ori_ori_n471_));
  NA3        o0443(.A(ori_ori_n471_), .B(ori_ori_n467_), .C(ori_ori_n314_), .Y(ori_ori_n472_));
  NOi41      o0444(.An(ori_ori_n452_), .B(ori_ori_n472_), .C(ori_ori_n465_), .D(ori_ori_n270_), .Y(ori_ori_n473_));
  NOi32      o0445(.An(c), .Bn(a), .C(b), .Y(ori_ori_n474_));
  NA2        o0446(.A(ori_ori_n474_), .B(ori_ori_n113_), .Y(ori_ori_n475_));
  INV        o0447(.A(ori_ori_n279_), .Y(ori_ori_n476_));
  AN2        o0448(.A(e), .B(d), .Y(ori_ori_n477_));
  NA2        o0449(.A(ori_ori_n477_), .B(ori_ori_n476_), .Y(ori_ori_n478_));
  INV        o0450(.A(ori_ori_n148_), .Y(ori_ori_n479_));
  NO2        o0451(.A(ori_ori_n130_), .B(ori_ori_n41_), .Y(ori_ori_n480_));
  NO2        o0452(.A(ori_ori_n66_), .B(e), .Y(ori_ori_n481_));
  NOi31      o0453(.An(j), .B(k), .C(i), .Y(ori_ori_n482_));
  NOi21      o0454(.An(ori_ori_n166_), .B(ori_ori_n482_), .Y(ori_ori_n483_));
  NA4        o0455(.A(ori_ori_n328_), .B(ori_ori_n483_), .C(ori_ori_n266_), .D(ori_ori_n118_), .Y(ori_ori_n484_));
  AOI220     o0456(.A0(ori_ori_n484_), .A1(ori_ori_n481_), .B0(ori_ori_n480_), .B1(ori_ori_n479_), .Y(ori_ori_n485_));
  AOI210     o0457(.A0(ori_ori_n485_), .A1(ori_ori_n478_), .B0(ori_ori_n475_), .Y(ori_ori_n486_));
  NO2        o0458(.A(ori_ori_n212_), .B(ori_ori_n207_), .Y(ori_ori_n487_));
  NOi21      o0459(.An(a), .B(b), .Y(ori_ori_n488_));
  NA3        o0460(.A(e), .B(d), .C(c), .Y(ori_ori_n489_));
  NAi21      o0461(.An(ori_ori_n489_), .B(ori_ori_n488_), .Y(ori_ori_n490_));
  AOI210     o0462(.A0(ori_ori_n273_), .A1(ori_ori_n487_), .B0(ori_ori_n490_), .Y(ori_ori_n491_));
  NO4        o0463(.A(ori_ori_n189_), .B(ori_ori_n103_), .C(ori_ori_n56_), .D(b), .Y(ori_ori_n492_));
  NA2        o0464(.A(ori_ori_n395_), .B(ori_ori_n154_), .Y(ori_ori_n493_));
  OR2        o0465(.A(k), .B(j), .Y(ori_ori_n494_));
  NA2        o0466(.A(l), .B(k), .Y(ori_ori_n495_));
  NA3        o0467(.A(ori_ori_n495_), .B(ori_ori_n494_), .C(ori_ori_n224_), .Y(ori_ori_n496_));
  AOI210     o0468(.A0(ori_ori_n237_), .A1(ori_ori_n346_), .B0(ori_ori_n84_), .Y(ori_ori_n497_));
  NOi21      o0469(.An(ori_ori_n496_), .B(ori_ori_n497_), .Y(ori_ori_n498_));
  OR3        o0470(.A(ori_ori_n498_), .B(ori_ori_n144_), .C(ori_ori_n134_), .Y(ori_ori_n499_));
  NA3        o0471(.A(ori_ori_n282_), .B(ori_ori_n127_), .C(ori_ori_n125_), .Y(ori_ori_n500_));
  NA2        o0472(.A(ori_ori_n408_), .B(ori_ori_n113_), .Y(ori_ori_n501_));
  NO4        o0473(.A(ori_ori_n501_), .B(ori_ori_n95_), .C(ori_ori_n112_), .D(e), .Y(ori_ori_n502_));
  NO3        o0474(.A(ori_ori_n502_), .B(ori_ori_n500_), .C(ori_ori_n329_), .Y(ori_ori_n503_));
  NA3        o0475(.A(ori_ori_n503_), .B(ori_ori_n499_), .C(ori_ori_n493_), .Y(ori_ori_n504_));
  NO4        o0476(.A(ori_ori_n504_), .B(ori_ori_n492_), .C(ori_ori_n491_), .D(ori_ori_n486_), .Y(ori_ori_n505_));
  NOi21      o0477(.An(d), .B(e), .Y(ori_ori_n506_));
  NO2        o0478(.A(ori_ori_n189_), .B(ori_ori_n56_), .Y(ori_ori_n507_));
  NAi31      o0479(.An(j), .B(l), .C(i), .Y(ori_ori_n508_));
  OAI210     o0480(.A0(ori_ori_n508_), .A1(ori_ori_n131_), .B0(ori_ori_n103_), .Y(ori_ori_n509_));
  NA4        o0481(.A(ori_ori_n509_), .B(ori_ori_n507_), .C(ori_ori_n506_), .D(b), .Y(ori_ori_n510_));
  NO3        o0482(.A(ori_ori_n409_), .B(ori_ori_n354_), .C(ori_ori_n203_), .Y(ori_ori_n511_));
  NO2        o0483(.A(ori_ori_n409_), .B(ori_ori_n384_), .Y(ori_ori_n512_));
  NO4        o0484(.A(ori_ori_n512_), .B(ori_ori_n511_), .C(ori_ori_n186_), .D(ori_ori_n311_), .Y(ori_ori_n513_));
  NA3        o0485(.A(ori_ori_n513_), .B(ori_ori_n510_), .C(ori_ori_n246_), .Y(ori_ori_n514_));
  OAI210     o0486(.A0(ori_ori_n126_), .A1(ori_ori_n124_), .B0(n), .Y(ori_ori_n515_));
  NO2        o0487(.A(ori_ori_n515_), .B(ori_ori_n130_), .Y(ori_ori_n516_));
  OR2        o0488(.A(ori_ori_n303_), .B(ori_ori_n248_), .Y(ori_ori_n517_));
  OA210      o0489(.A0(ori_ori_n517_), .A1(ori_ori_n516_), .B0(ori_ori_n194_), .Y(ori_ori_n518_));
  XO2        o0490(.A(i), .B(h), .Y(ori_ori_n519_));
  NA3        o0491(.A(ori_ori_n519_), .B(ori_ori_n161_), .C(n), .Y(ori_ori_n520_));
  NAi41      o0492(.An(ori_ori_n303_), .B(ori_ori_n520_), .C(ori_ori_n469_), .D(ori_ori_n397_), .Y(ori_ori_n521_));
  NOi32      o0493(.An(ori_ori_n521_), .Bn(ori_ori_n481_), .C(ori_ori_n275_), .Y(ori_ori_n522_));
  NAi31      o0494(.An(c), .B(f), .C(d), .Y(ori_ori_n523_));
  AOI210     o0495(.A0(ori_ori_n283_), .A1(ori_ori_n197_), .B0(ori_ori_n523_), .Y(ori_ori_n524_));
  NOi21      o0496(.An(ori_ori_n82_), .B(ori_ori_n524_), .Y(ori_ori_n525_));
  NA2        o0497(.A(ori_ori_n231_), .B(ori_ori_n109_), .Y(ori_ori_n526_));
  AOI210     o0498(.A0(ori_ori_n526_), .A1(ori_ori_n182_), .B0(ori_ori_n523_), .Y(ori_ori_n527_));
  INV        o0499(.A(ori_ori_n527_), .Y(ori_ori_n528_));
  AO220      o0500(.A0(ori_ori_n291_), .A1(ori_ori_n268_), .B0(ori_ori_n167_), .B1(ori_ori_n67_), .Y(ori_ori_n529_));
  NA3        o0501(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(f), .Y(ori_ori_n530_));
  INV        o0502(.A(ori_ori_n299_), .Y(ori_ori_n531_));
  NAi41      o0503(.An(ori_ori_n529_), .B(ori_ori_n531_), .C(ori_ori_n528_), .D(ori_ori_n525_), .Y(ori_ori_n532_));
  NO4        o0504(.A(ori_ori_n532_), .B(ori_ori_n522_), .C(ori_ori_n518_), .D(ori_ori_n514_), .Y(ori_ori_n533_));
  NA4        o0505(.A(ori_ori_n533_), .B(ori_ori_n505_), .C(ori_ori_n473_), .D(ori_ori_n446_), .Y(ori11));
  NO2        o0506(.A(ori_ori_n72_), .B(f), .Y(ori_ori_n535_));
  NA2        o0507(.A(j), .B(o), .Y(ori_ori_n536_));
  NAi31      o0508(.An(i), .B(m), .C(l), .Y(ori_ori_n537_));
  NA3        o0509(.A(m), .B(k), .C(j), .Y(ori_ori_n538_));
  OAI220     o0510(.A0(ori_ori_n538_), .A1(ori_ori_n130_), .B0(ori_ori_n537_), .B1(ori_ori_n536_), .Y(ori_ori_n539_));
  NA2        o0511(.A(ori_ori_n539_), .B(ori_ori_n535_), .Y(ori_ori_n540_));
  NOi32      o0512(.An(e), .Bn(b), .C(f), .Y(ori_ori_n541_));
  NA2        o0513(.A(ori_ori_n46_), .B(j), .Y(ori_ori_n542_));
  NO2        o0514(.A(ori_ori_n542_), .B(ori_ori_n305_), .Y(ori_ori_n543_));
  NAi31      o0515(.An(d), .B(e), .C(a), .Y(ori_ori_n544_));
  NO2        o0516(.A(ori_ori_n544_), .B(n), .Y(ori_ori_n545_));
  NA2        o0517(.A(ori_ori_n543_), .B(ori_ori_n541_), .Y(ori_ori_n546_));
  NAi41      o0518(.An(f), .B(e), .C(c), .D(a), .Y(ori_ori_n547_));
  AN2        o0519(.A(ori_ori_n547_), .B(ori_ori_n383_), .Y(ori_ori_n548_));
  NA2        o0520(.A(j), .B(i), .Y(ori_ori_n549_));
  NAi31      o0521(.An(n), .B(m), .C(k), .Y(ori_ori_n550_));
  NO3        o0522(.A(ori_ori_n550_), .B(ori_ori_n549_), .C(ori_ori_n112_), .Y(ori_ori_n551_));
  NO4        o0523(.A(n), .B(d), .C(ori_ori_n115_), .D(a), .Y(ori_ori_n552_));
  OR2        o0524(.A(n), .B(c), .Y(ori_ori_n553_));
  NO2        o0525(.A(ori_ori_n553_), .B(ori_ori_n150_), .Y(ori_ori_n554_));
  NO2        o0526(.A(ori_ori_n554_), .B(ori_ori_n552_), .Y(ori_ori_n555_));
  NOi32      o0527(.An(o), .Bn(f), .C(i), .Y(ori_ori_n556_));
  AOI220     o0528(.A0(ori_ori_n556_), .A1(ori_ori_n100_), .B0(ori_ori_n539_), .B1(f), .Y(ori_ori_n557_));
  NO2        o0529(.A(ori_ori_n279_), .B(ori_ori_n49_), .Y(ori_ori_n558_));
  NO2        o0530(.A(ori_ori_n557_), .B(ori_ori_n555_), .Y(ori_ori_n559_));
  INV        o0531(.A(ori_ori_n559_), .Y(ori_ori_n560_));
  NA2        o0532(.A(ori_ori_n140_), .B(ori_ori_n34_), .Y(ori_ori_n561_));
  OAI220     o0533(.A0(ori_ori_n561_), .A1(m), .B0(ori_ori_n542_), .B1(ori_ori_n237_), .Y(ori_ori_n562_));
  NOi41      o0534(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n563_));
  NAi32      o0535(.An(e), .Bn(b), .C(c), .Y(ori_ori_n564_));
  OR2        o0536(.A(ori_ori_n564_), .B(ori_ori_n84_), .Y(ori_ori_n565_));
  AN2        o0537(.A(ori_ori_n347_), .B(ori_ori_n325_), .Y(ori_ori_n566_));
  NA2        o0538(.A(ori_ori_n566_), .B(ori_ori_n565_), .Y(ori_ori_n567_));
  OA210      o0539(.A0(ori_ori_n567_), .A1(ori_ori_n563_), .B0(ori_ori_n562_), .Y(ori_ori_n568_));
  OAI220     o0540(.A0(ori_ori_n411_), .A1(ori_ori_n410_), .B0(ori_ori_n537_), .B1(ori_ori_n536_), .Y(ori_ori_n569_));
  NAi31      o0541(.An(d), .B(c), .C(a), .Y(ori_ori_n570_));
  NO2        o0542(.A(ori_ori_n570_), .B(n), .Y(ori_ori_n571_));
  NA3        o0543(.A(ori_ori_n571_), .B(ori_ori_n569_), .C(e), .Y(ori_ori_n572_));
  INV        o0544(.A(ori_ori_n572_), .Y(ori_ori_n573_));
  NO2        o0545(.A(ori_ori_n280_), .B(n), .Y(ori_ori_n574_));
  NO2        o0546(.A(ori_ori_n441_), .B(ori_ori_n574_), .Y(ori_ori_n575_));
  NA2        o0547(.A(ori_ori_n569_), .B(f), .Y(ori_ori_n576_));
  NAi32      o0548(.An(d), .Bn(a), .C(b), .Y(ori_ori_n577_));
  NA2        o0549(.A(h), .B(f), .Y(ori_ori_n578_));
  NO2        o0550(.A(ori_ori_n578_), .B(ori_ori_n95_), .Y(ori_ori_n579_));
  NO3        o0551(.A(ori_ori_n178_), .B(ori_ori_n175_), .C(o), .Y(ori_ori_n580_));
  NA2        o0552(.A(ori_ori_n580_), .B(ori_ori_n58_), .Y(ori_ori_n581_));
  OAI210     o0553(.A0(ori_ori_n576_), .A1(ori_ori_n575_), .B0(ori_ori_n581_), .Y(ori_ori_n582_));
  AN3        o0554(.A(j), .B(h), .C(o), .Y(ori_ori_n583_));
  NO2        o0555(.A(ori_ori_n147_), .B(c), .Y(ori_ori_n584_));
  NA3        o0556(.A(ori_ori_n584_), .B(ori_ori_n583_), .C(ori_ori_n468_), .Y(ori_ori_n585_));
  NA3        o0557(.A(f), .B(d), .C(b), .Y(ori_ori_n586_));
  NO4        o0558(.A(ori_ori_n586_), .B(ori_ori_n178_), .C(ori_ori_n175_), .D(o), .Y(ori_ori_n587_));
  NAi21      o0559(.An(ori_ori_n587_), .B(ori_ori_n585_), .Y(ori_ori_n588_));
  NO4        o0560(.A(ori_ori_n588_), .B(ori_ori_n582_), .C(ori_ori_n573_), .D(ori_ori_n568_), .Y(ori_ori_n589_));
  AN4        o0561(.A(ori_ori_n589_), .B(ori_ori_n560_), .C(ori_ori_n546_), .D(ori_ori_n540_), .Y(ori_ori_n590_));
  INV        o0562(.A(k), .Y(ori_ori_n591_));
  NA3        o0563(.A(l), .B(ori_ori_n591_), .C(i), .Y(ori_ori_n592_));
  INV        o0564(.A(ori_ori_n592_), .Y(ori_ori_n593_));
  NAi32      o0565(.An(h), .Bn(f), .C(o), .Y(ori_ori_n594_));
  NAi41      o0566(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n595_));
  OAI210     o0567(.A0(ori_ori_n544_), .A1(n), .B0(ori_ori_n595_), .Y(ori_ori_n596_));
  NA2        o0568(.A(ori_ori_n596_), .B(m), .Y(ori_ori_n597_));
  NAi31      o0569(.An(h), .B(o), .C(f), .Y(ori_ori_n598_));
  OR3        o0570(.A(ori_ori_n598_), .B(ori_ori_n280_), .C(ori_ori_n49_), .Y(ori_ori_n599_));
  NA4        o0571(.A(ori_ori_n431_), .B(ori_ori_n120_), .C(ori_ori_n113_), .D(e), .Y(ori_ori_n600_));
  AN2        o0572(.A(ori_ori_n600_), .B(ori_ori_n599_), .Y(ori_ori_n601_));
  NO3        o0573(.A(ori_ori_n594_), .B(ori_ori_n72_), .C(ori_ori_n73_), .Y(ori_ori_n602_));
  NO4        o0574(.A(ori_ori_n598_), .B(ori_ori_n553_), .C(ori_ori_n150_), .D(ori_ori_n73_), .Y(ori_ori_n603_));
  OR2        o0575(.A(ori_ori_n603_), .B(ori_ori_n602_), .Y(ori_ori_n604_));
  NAi21      o0576(.An(ori_ori_n604_), .B(ori_ori_n601_), .Y(ori_ori_n605_));
  NAi31      o0577(.An(f), .B(h), .C(o), .Y(ori_ori_n606_));
  NOi32      o0578(.An(b), .Bn(a), .C(c), .Y(ori_ori_n607_));
  NOi41      o0579(.An(ori_ori_n607_), .B(ori_ori_n363_), .C(ori_ori_n69_), .D(ori_ori_n116_), .Y(ori_ori_n608_));
  NOi32      o0580(.An(d), .Bn(a), .C(e), .Y(ori_ori_n609_));
  NA2        o0581(.A(ori_ori_n609_), .B(ori_ori_n113_), .Y(ori_ori_n610_));
  NO2        o0582(.A(n), .B(c), .Y(ori_ori_n611_));
  NA3        o0583(.A(ori_ori_n611_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n612_));
  NAi32      o0584(.An(n), .Bn(f), .C(m), .Y(ori_ori_n613_));
  NA3        o0585(.A(ori_ori_n613_), .B(ori_ori_n612_), .C(ori_ori_n610_), .Y(ori_ori_n614_));
  NOi32      o0586(.An(e), .Bn(a), .C(d), .Y(ori_ori_n615_));
  AOI210     o0587(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n615_), .Y(ori_ori_n616_));
  AOI210     o0588(.A0(ori_ori_n616_), .A1(ori_ori_n216_), .B0(ori_ori_n561_), .Y(ori_ori_n617_));
  AOI210     o0589(.A0(ori_ori_n617_), .A1(ori_ori_n614_), .B0(ori_ori_n608_), .Y(ori_ori_n618_));
  OAI210     o0590(.A0(ori_ori_n253_), .A1(ori_ori_n87_), .B0(ori_ori_n618_), .Y(ori_ori_n619_));
  AOI210     o0591(.A0(ori_ori_n605_), .A1(ori_ori_n593_), .B0(ori_ori_n619_), .Y(ori_ori_n620_));
  NO3        o0592(.A(ori_ori_n323_), .B(ori_ori_n61_), .C(n), .Y(ori_ori_n621_));
  NA3        o0593(.A(ori_ori_n523_), .B(ori_ori_n173_), .C(ori_ori_n172_), .Y(ori_ori_n622_));
  NA2        o0594(.A(ori_ori_n470_), .B(ori_ori_n234_), .Y(ori_ori_n623_));
  OR2        o0595(.A(ori_ori_n623_), .B(ori_ori_n622_), .Y(ori_ori_n624_));
  NA2        o0596(.A(ori_ori_n74_), .B(ori_ori_n113_), .Y(ori_ori_n625_));
  NA2        o0597(.A(ori_ori_n624_), .B(ori_ori_n621_), .Y(ori_ori_n626_));
  NO2        o0598(.A(ori_ori_n626_), .B(ori_ori_n87_), .Y(ori_ori_n627_));
  NA3        o0599(.A(ori_ori_n563_), .B(ori_ori_n349_), .C(ori_ori_n46_), .Y(ori_ori_n628_));
  NOi32      o0600(.An(e), .Bn(c), .C(f), .Y(ori_ori_n629_));
  NOi21      o0601(.An(f), .B(o), .Y(ori_ori_n630_));
  NO2        o0602(.A(ori_ori_n630_), .B(ori_ori_n214_), .Y(ori_ori_n631_));
  AOI220     o0603(.A0(ori_ori_n631_), .A1(ori_ori_n405_), .B0(ori_ori_n629_), .B1(ori_ori_n177_), .Y(ori_ori_n632_));
  NA3        o0604(.A(ori_ori_n632_), .B(ori_ori_n628_), .C(ori_ori_n180_), .Y(ori_ori_n633_));
  AOI210     o0605(.A0(ori_ori_n548_), .A1(ori_ori_n409_), .B0(ori_ori_n304_), .Y(ori_ori_n634_));
  NA2        o0606(.A(ori_ori_n634_), .B(ori_ori_n269_), .Y(ori_ori_n635_));
  NOi21      o0607(.An(j), .B(l), .Y(ori_ori_n636_));
  NAi21      o0608(.An(k), .B(h), .Y(ori_ori_n637_));
  NO2        o0609(.A(ori_ori_n637_), .B(ori_ori_n267_), .Y(ori_ori_n638_));
  NA2        o0610(.A(ori_ori_n638_), .B(ori_ori_n636_), .Y(ori_ori_n639_));
  OR2        o0611(.A(ori_ori_n639_), .B(ori_ori_n597_), .Y(ori_ori_n640_));
  NOi31      o0612(.An(m), .B(n), .C(k), .Y(ori_ori_n641_));
  NA2        o0613(.A(ori_ori_n636_), .B(ori_ori_n641_), .Y(ori_ori_n642_));
  AOI210     o0614(.A0(ori_ori_n409_), .A1(ori_ori_n383_), .B0(ori_ori_n304_), .Y(ori_ori_n643_));
  NAi21      o0615(.An(ori_ori_n642_), .B(ori_ori_n643_), .Y(ori_ori_n644_));
  NO2        o0616(.A(ori_ori_n280_), .B(ori_ori_n49_), .Y(ori_ori_n645_));
  NO2        o0617(.A(ori_ori_n316_), .B(ori_ori_n606_), .Y(ori_ori_n646_));
  NO2        o0618(.A(ori_ori_n544_), .B(ori_ori_n49_), .Y(ori_ori_n647_));
  NA2        o0619(.A(ori_ori_n647_), .B(ori_ori_n646_), .Y(ori_ori_n648_));
  NA4        o0620(.A(ori_ori_n648_), .B(ori_ori_n644_), .C(ori_ori_n640_), .D(ori_ori_n635_), .Y(ori_ori_n649_));
  NA2        o0621(.A(ori_ori_n109_), .B(ori_ori_n36_), .Y(ori_ori_n650_));
  NO2        o0622(.A(k), .B(ori_ori_n217_), .Y(ori_ori_n651_));
  INV        o0623(.A(ori_ori_n372_), .Y(ori_ori_n652_));
  NO2        o0624(.A(ori_ori_n652_), .B(n), .Y(ori_ori_n653_));
  NAi31      o0625(.An(ori_ori_n650_), .B(ori_ori_n653_), .C(ori_ori_n651_), .Y(ori_ori_n654_));
  NO2        o0626(.A(ori_ori_n542_), .B(ori_ori_n178_), .Y(ori_ori_n655_));
  NA3        o0627(.A(ori_ori_n564_), .B(ori_ori_n275_), .C(ori_ori_n145_), .Y(ori_ori_n656_));
  NA2        o0628(.A(ori_ori_n519_), .B(ori_ori_n161_), .Y(ori_ori_n657_));
  NO3        o0629(.A(ori_ori_n406_), .B(ori_ori_n657_), .C(ori_ori_n87_), .Y(ori_ori_n658_));
  AOI210     o0630(.A0(ori_ori_n656_), .A1(ori_ori_n655_), .B0(ori_ori_n658_), .Y(ori_ori_n659_));
  AN3        o0631(.A(f), .B(d), .C(b), .Y(ori_ori_n660_));
  OAI210     o0632(.A0(ori_ori_n660_), .A1(ori_ori_n129_), .B0(n), .Y(ori_ori_n661_));
  NA3        o0633(.A(ori_ori_n519_), .B(ori_ori_n161_), .C(ori_ori_n217_), .Y(ori_ori_n662_));
  AOI210     o0634(.A0(ori_ori_n661_), .A1(ori_ori_n236_), .B0(ori_ori_n662_), .Y(ori_ori_n663_));
  NAi31      o0635(.An(m), .B(n), .C(k), .Y(ori_ori_n664_));
  OR2        o0636(.A(ori_ori_n134_), .B(ori_ori_n61_), .Y(ori_ori_n665_));
  OAI210     o0637(.A0(ori_ori_n665_), .A1(ori_ori_n664_), .B0(ori_ori_n255_), .Y(ori_ori_n666_));
  OAI210     o0638(.A0(ori_ori_n666_), .A1(ori_ori_n663_), .B0(j), .Y(ori_ori_n667_));
  NA3        o0639(.A(ori_ori_n667_), .B(ori_ori_n659_), .C(ori_ori_n654_), .Y(ori_ori_n668_));
  NO4        o0640(.A(ori_ori_n668_), .B(ori_ori_n649_), .C(ori_ori_n633_), .D(ori_ori_n627_), .Y(ori_ori_n669_));
  NA2        o0641(.A(ori_ori_n393_), .B(ori_ori_n164_), .Y(ori_ori_n670_));
  NAi31      o0642(.An(o), .B(h), .C(f), .Y(ori_ori_n671_));
  OR3        o0643(.A(ori_ori_n671_), .B(ori_ori_n280_), .C(n), .Y(ori_ori_n672_));
  OA210      o0644(.A0(ori_ori_n544_), .A1(n), .B0(ori_ori_n595_), .Y(ori_ori_n673_));
  NA3        o0645(.A(ori_ori_n429_), .B(ori_ori_n120_), .C(ori_ori_n84_), .Y(ori_ori_n674_));
  OAI210     o0646(.A0(ori_ori_n673_), .A1(ori_ori_n91_), .B0(ori_ori_n674_), .Y(ori_ori_n675_));
  NOi21      o0647(.An(ori_ori_n672_), .B(ori_ori_n675_), .Y(ori_ori_n676_));
  AOI210     o0648(.A0(ori_ori_n676_), .A1(ori_ori_n670_), .B0(ori_ori_n538_), .Y(ori_ori_n677_));
  NO3        o0649(.A(o), .B(ori_ori_n216_), .C(ori_ori_n56_), .Y(ori_ori_n678_));
  NAi21      o0650(.An(h), .B(j), .Y(ori_ori_n679_));
  NO2        o0651(.A(ori_ori_n526_), .B(ori_ori_n87_), .Y(ori_ori_n680_));
  OAI210     o0652(.A0(ori_ori_n680_), .A1(ori_ori_n405_), .B0(ori_ori_n678_), .Y(ori_ori_n681_));
  OR2        o0653(.A(ori_ori_n72_), .B(ori_ori_n73_), .Y(ori_ori_n682_));
  NA2        o0654(.A(ori_ori_n607_), .B(ori_ori_n351_), .Y(ori_ori_n683_));
  OA220      o0655(.A0(ori_ori_n642_), .A1(ori_ori_n683_), .B0(ori_ori_n639_), .B1(ori_ori_n682_), .Y(ori_ori_n684_));
  NA3        o0656(.A(ori_ori_n535_), .B(ori_ori_n100_), .C(ori_ori_n99_), .Y(ori_ori_n685_));
  AN2        o0657(.A(h), .B(f), .Y(ori_ori_n686_));
  NA2        o0658(.A(ori_ori_n686_), .B(ori_ori_n37_), .Y(ori_ori_n687_));
  NA2        o0659(.A(ori_ori_n100_), .B(ori_ori_n46_), .Y(ori_ori_n688_));
  OAI220     o0660(.A0(ori_ori_n688_), .A1(ori_ori_n340_), .B0(ori_ori_n687_), .B1(ori_ori_n475_), .Y(ori_ori_n689_));
  AOI210     o0661(.A0(ori_ori_n577_), .A1(ori_ori_n440_), .B0(ori_ori_n49_), .Y(ori_ori_n690_));
  OAI220     o0662(.A0(ori_ori_n598_), .A1(ori_ori_n592_), .B0(ori_ori_n333_), .B1(ori_ori_n536_), .Y(ori_ori_n691_));
  AOI210     o0663(.A0(ori_ori_n691_), .A1(ori_ori_n690_), .B0(ori_ori_n689_), .Y(ori_ori_n692_));
  NA4        o0664(.A(ori_ori_n692_), .B(ori_ori_n685_), .C(ori_ori_n684_), .D(ori_ori_n681_), .Y(ori_ori_n693_));
  NO2        o0665(.A(ori_ori_n630_), .B(ori_ori_n61_), .Y(ori_ori_n694_));
  NO2        o0666(.A(ori_ori_n694_), .B(ori_ori_n34_), .Y(ori_ori_n695_));
  NA2        o0667(.A(ori_ori_n336_), .B(ori_ori_n140_), .Y(ori_ori_n696_));
  NA2        o0668(.A(ori_ori_n131_), .B(ori_ori_n49_), .Y(ori_ori_n697_));
  AOI220     o0669(.A0(ori_ori_n697_), .A1(ori_ori_n541_), .B0(ori_ori_n372_), .B1(ori_ori_n113_), .Y(ori_ori_n698_));
  OA220      o0670(.A0(ori_ori_n698_), .A1(ori_ori_n561_), .B0(ori_ori_n370_), .B1(ori_ori_n111_), .Y(ori_ori_n699_));
  OAI210     o0671(.A0(ori_ori_n696_), .A1(ori_ori_n695_), .B0(ori_ori_n699_), .Y(ori_ori_n700_));
  NO3        o0672(.A(ori_ori_n416_), .B(ori_ori_n194_), .C(ori_ori_n193_), .Y(ori_ori_n701_));
  NA2        o0673(.A(ori_ori_n701_), .B(ori_ori_n234_), .Y(ori_ori_n702_));
  NA3        o0674(.A(ori_ori_n702_), .B(ori_ori_n259_), .C(j), .Y(ori_ori_n703_));
  NO3        o0675(.A(ori_ori_n470_), .B(ori_ori_n175_), .C(i), .Y(ori_ori_n704_));
  NA2        o0676(.A(ori_ori_n474_), .B(ori_ori_n84_), .Y(ori_ori_n705_));
  NA2        o0677(.A(ori_ori_n703_), .B(ori_ori_n414_), .Y(ori_ori_n706_));
  NO4        o0678(.A(ori_ori_n706_), .B(ori_ori_n700_), .C(ori_ori_n693_), .D(ori_ori_n677_), .Y(ori_ori_n707_));
  NA4        o0679(.A(ori_ori_n707_), .B(ori_ori_n669_), .C(ori_ori_n620_), .D(ori_ori_n590_), .Y(ori08));
  NO2        o0680(.A(k), .B(h), .Y(ori_ori_n709_));
  AO210      o0681(.A0(ori_ori_n257_), .A1(ori_ori_n460_), .B0(ori_ori_n709_), .Y(ori_ori_n710_));
  NO2        o0682(.A(ori_ori_n710_), .B(ori_ori_n302_), .Y(ori_ori_n711_));
  NA2        o0683(.A(ori_ori_n629_), .B(ori_ori_n84_), .Y(ori_ori_n712_));
  NA2        o0684(.A(ori_ori_n712_), .B(ori_ori_n470_), .Y(ori_ori_n713_));
  NA2        o0685(.A(ori_ori_n713_), .B(ori_ori_n711_), .Y(ori_ori_n714_));
  NA2        o0686(.A(ori_ori_n84_), .B(ori_ori_n110_), .Y(ori_ori_n715_));
  NO2        o0687(.A(ori_ori_n715_), .B(ori_ori_n57_), .Y(ori_ori_n716_));
  NO4        o0688(.A(ori_ori_n390_), .B(ori_ori_n112_), .C(j), .D(ori_ori_n217_), .Y(ori_ori_n717_));
  NA2        o0689(.A(ori_ori_n586_), .B(ori_ori_n236_), .Y(ori_ori_n718_));
  AOI220     o0690(.A0(ori_ori_n718_), .A1(ori_ori_n357_), .B0(ori_ori_n717_), .B1(ori_ori_n716_), .Y(ori_ori_n719_));
  AOI210     o0691(.A0(ori_ori_n586_), .A1(ori_ori_n157_), .B0(ori_ori_n84_), .Y(ori_ori_n720_));
  NA4        o0692(.A(ori_ori_n219_), .B(ori_ori_n140_), .C(ori_ori_n45_), .D(h), .Y(ori_ori_n721_));
  AN2        o0693(.A(l), .B(k), .Y(ori_ori_n722_));
  NA4        o0694(.A(ori_ori_n722_), .B(ori_ori_n109_), .C(ori_ori_n73_), .D(ori_ori_n217_), .Y(ori_ori_n723_));
  NA3        o0695(.A(ori_ori_n719_), .B(ori_ori_n714_), .C(ori_ori_n359_), .Y(ori_ori_n724_));
  AN2        o0696(.A(ori_ori_n545_), .B(ori_ori_n96_), .Y(ori_ori_n725_));
  NO4        o0697(.A(ori_ori_n175_), .B(ori_ori_n404_), .C(ori_ori_n112_), .D(o), .Y(ori_ori_n726_));
  NA2        o0698(.A(ori_ori_n726_), .B(ori_ori_n718_), .Y(ori_ori_n727_));
  NA2        o0699(.A(ori_ori_n631_), .B(ori_ori_n356_), .Y(ori_ori_n728_));
  NAi31      o0700(.An(ori_ori_n725_), .B(ori_ori_n728_), .C(ori_ori_n727_), .Y(ori_ori_n729_));
  NO2        o0701(.A(ori_ori_n548_), .B(ori_ori_n35_), .Y(ori_ori_n730_));
  OAI210     o0702(.A0(ori_ori_n564_), .A1(ori_ori_n47_), .B0(ori_ori_n665_), .Y(ori_ori_n731_));
  NO2        o0703(.A(ori_ori_n495_), .B(ori_ori_n131_), .Y(ori_ori_n732_));
  AOI210     o0704(.A0(ori_ori_n732_), .A1(ori_ori_n731_), .B0(ori_ori_n730_), .Y(ori_ori_n733_));
  NO3        o0705(.A(ori_ori_n323_), .B(ori_ori_n130_), .C(ori_ori_n41_), .Y(ori_ori_n734_));
  NAi21      o0706(.An(ori_ori_n734_), .B(ori_ori_n723_), .Y(ori_ori_n735_));
  NA2        o0707(.A(ori_ori_n710_), .B(ori_ori_n135_), .Y(ori_ori_n736_));
  AOI220     o0708(.A0(ori_ori_n736_), .A1(ori_ori_n415_), .B0(ori_ori_n735_), .B1(ori_ori_n76_), .Y(ori_ori_n737_));
  OAI210     o0709(.A0(ori_ori_n733_), .A1(ori_ori_n87_), .B0(ori_ori_n737_), .Y(ori_ori_n738_));
  NA2        o0710(.A(ori_ori_n372_), .B(ori_ori_n43_), .Y(ori_ori_n739_));
  NA3        o0711(.A(ori_ori_n702_), .B(ori_ori_n342_), .C(ori_ori_n396_), .Y(ori_ori_n740_));
  INV        o0712(.A(ori_ori_n502_), .Y(ori_ori_n741_));
  NA3        o0713(.A(m), .B(l), .C(k), .Y(ori_ori_n742_));
  AOI210     o0714(.A0(ori_ori_n674_), .A1(ori_ori_n672_), .B0(ori_ori_n742_), .Y(ori_ori_n743_));
  NA4        o0715(.A(ori_ori_n113_), .B(l), .C(k), .D(ori_ori_n87_), .Y(ori_ori_n744_));
  INV        o0716(.A(ori_ori_n743_), .Y(ori_ori_n745_));
  NA4        o0717(.A(ori_ori_n745_), .B(ori_ori_n741_), .C(ori_ori_n740_), .D(ori_ori_n739_), .Y(ori_ori_n746_));
  NO4        o0718(.A(ori_ori_n746_), .B(ori_ori_n738_), .C(ori_ori_n729_), .D(ori_ori_n724_), .Y(ori_ori_n747_));
  NA2        o0719(.A(ori_ori_n631_), .B(ori_ori_n405_), .Y(ori_ori_n748_));
  INV        o0720(.A(ori_ori_n512_), .Y(ori_ori_n749_));
  NA3        o0721(.A(ori_ori_n749_), .B(ori_ori_n748_), .C(ori_ori_n256_), .Y(ori_ori_n750_));
  NA2        o0722(.A(ori_ori_n722_), .B(ori_ori_n73_), .Y(ori_ori_n751_));
  NO4        o0723(.A(ori_ori_n701_), .B(ori_ori_n175_), .C(n), .D(i), .Y(ori_ori_n752_));
  NOi21      o0724(.An(h), .B(j), .Y(ori_ori_n753_));
  NA2        o0725(.A(ori_ori_n753_), .B(f), .Y(ori_ori_n754_));
  NO2        o0726(.A(ori_ori_n754_), .B(ori_ori_n250_), .Y(ori_ori_n755_));
  NO3        o0727(.A(ori_ori_n755_), .B(ori_ori_n752_), .C(ori_ori_n704_), .Y(ori_ori_n756_));
  OAI220     o0728(.A0(ori_ori_n756_), .A1(ori_ori_n751_), .B0(ori_ori_n601_), .B1(ori_ori_n62_), .Y(ori_ori_n757_));
  AOI210     o0729(.A0(ori_ori_n750_), .A1(l), .B0(ori_ori_n757_), .Y(ori_ori_n758_));
  NO2        o0730(.A(j), .B(i), .Y(ori_ori_n759_));
  NA3        o0731(.A(ori_ori_n759_), .B(ori_ori_n80_), .C(l), .Y(ori_ori_n760_));
  NA2        o0732(.A(ori_ori_n759_), .B(ori_ori_n33_), .Y(ori_ori_n761_));
  NA2        o0733(.A(ori_ori_n434_), .B(ori_ori_n120_), .Y(ori_ori_n762_));
  OA220      o0734(.A0(ori_ori_n762_), .A1(ori_ori_n761_), .B0(ori_ori_n760_), .B1(ori_ori_n597_), .Y(ori_ori_n763_));
  NO3        o0735(.A(ori_ori_n152_), .B(ori_ori_n49_), .C(ori_ori_n110_), .Y(ori_ori_n764_));
  NO3        o0736(.A(ori_ori_n553_), .B(ori_ori_n150_), .C(ori_ori_n73_), .Y(ori_ori_n765_));
  NO3        o0737(.A(ori_ori_n495_), .B(ori_ori_n450_), .C(j), .Y(ori_ori_n766_));
  OAI210     o0738(.A0(ori_ori_n765_), .A1(ori_ori_n764_), .B0(ori_ori_n766_), .Y(ori_ori_n767_));
  INV        o0739(.A(ori_ori_n767_), .Y(ori_ori_n768_));
  NA2        o0740(.A(k), .B(j), .Y(ori_ori_n769_));
  NO3        o0741(.A(ori_ori_n302_), .B(ori_ori_n769_), .C(ori_ori_n40_), .Y(ori_ori_n770_));
  AOI210     o0742(.A0(ori_ori_n541_), .A1(n), .B0(ori_ori_n563_), .Y(ori_ori_n771_));
  NA2        o0743(.A(ori_ori_n771_), .B(ori_ori_n566_), .Y(ori_ori_n772_));
  AN3        o0744(.A(ori_ori_n772_), .B(ori_ori_n770_), .C(ori_ori_n99_), .Y(ori_ori_n773_));
  NO3        o0745(.A(ori_ori_n175_), .B(ori_ori_n404_), .C(ori_ori_n112_), .Y(ori_ori_n774_));
  AOI220     o0746(.A0(ori_ori_n774_), .A1(ori_ori_n251_), .B0(ori_ori_n623_), .B1(ori_ori_n313_), .Y(ori_ori_n775_));
  NAi31      o0747(.An(ori_ori_n616_), .B(ori_ori_n93_), .C(ori_ori_n84_), .Y(ori_ori_n776_));
  NA2        o0748(.A(ori_ori_n776_), .B(ori_ori_n775_), .Y(ori_ori_n777_));
  NO2        o0749(.A(ori_ori_n302_), .B(ori_ori_n135_), .Y(ori_ori_n778_));
  AOI220     o0750(.A0(ori_ori_n778_), .A1(ori_ori_n631_), .B0(ori_ori_n734_), .B1(ori_ori_n720_), .Y(ori_ori_n779_));
  NO2        o0751(.A(ori_ori_n742_), .B(ori_ori_n91_), .Y(ori_ori_n780_));
  NA2        o0752(.A(ori_ori_n780_), .B(ori_ori_n596_), .Y(ori_ori_n781_));
  NO2        o0753(.A(ori_ori_n598_), .B(ori_ori_n116_), .Y(ori_ori_n782_));
  OAI210     o0754(.A0(ori_ori_n782_), .A1(ori_ori_n766_), .B0(ori_ori_n690_), .Y(ori_ori_n783_));
  NA3        o0755(.A(ori_ori_n783_), .B(ori_ori_n781_), .C(ori_ori_n779_), .Y(ori_ori_n784_));
  OR4        o0756(.A(ori_ori_n784_), .B(ori_ori_n777_), .C(ori_ori_n773_), .D(ori_ori_n768_), .Y(ori_ori_n785_));
  NA3        o0757(.A(ori_ori_n771_), .B(ori_ori_n566_), .C(ori_ori_n565_), .Y(ori_ori_n786_));
  NA4        o0758(.A(ori_ori_n786_), .B(ori_ori_n219_), .C(ori_ori_n460_), .D(ori_ori_n34_), .Y(ori_ori_n787_));
  NO4        o0759(.A(ori_ori_n495_), .B(ori_ori_n447_), .C(j), .D(f), .Y(ori_ori_n788_));
  OAI220     o0760(.A0(ori_ori_n721_), .A1(ori_ori_n712_), .B0(ori_ori_n340_), .B1(ori_ori_n38_), .Y(ori_ori_n789_));
  INV        o0761(.A(ori_ori_n789_), .Y(ori_ori_n790_));
  NA3        o0762(.A(ori_ori_n556_), .B(ori_ori_n295_), .C(h), .Y(ori_ori_n791_));
  NO2        o0763(.A(ori_ori_n92_), .B(ori_ori_n47_), .Y(ori_ori_n792_));
  NO2        o0764(.A(ori_ori_n791_), .B(ori_ori_n612_), .Y(ori_ori_n793_));
  AOI210     o0765(.A0(ori_ori_n792_), .A1(ori_ori_n653_), .B0(ori_ori_n793_), .Y(ori_ori_n794_));
  NA3        o0766(.A(ori_ori_n794_), .B(ori_ori_n790_), .C(ori_ori_n787_), .Y(ori_ori_n795_));
  NA2        o0767(.A(ori_ori_n780_), .B(ori_ori_n242_), .Y(ori_ori_n796_));
  NO2        o0768(.A(ori_ori_n673_), .B(ori_ori_n73_), .Y(ori_ori_n797_));
  AOI210     o0769(.A0(ori_ori_n788_), .A1(ori_ori_n797_), .B0(ori_ori_n344_), .Y(ori_ori_n798_));
  OAI210     o0770(.A0(ori_ori_n742_), .A1(ori_ori_n671_), .B0(ori_ori_n530_), .Y(ori_ori_n799_));
  NA3        o0771(.A(ori_ori_n254_), .B(ori_ori_n59_), .C(b), .Y(ori_ori_n800_));
  AOI220     o0772(.A0(ori_ori_n611_), .A1(ori_ori_n29_), .B0(ori_ori_n474_), .B1(ori_ori_n84_), .Y(ori_ori_n801_));
  NA2        o0773(.A(ori_ori_n801_), .B(ori_ori_n800_), .Y(ori_ori_n802_));
  NO2        o0774(.A(ori_ori_n791_), .B(ori_ori_n501_), .Y(ori_ori_n803_));
  AOI210     o0775(.A0(ori_ori_n802_), .A1(ori_ori_n799_), .B0(ori_ori_n803_), .Y(ori_ori_n804_));
  NA3        o0776(.A(ori_ori_n804_), .B(ori_ori_n798_), .C(ori_ori_n796_), .Y(ori_ori_n805_));
  NOi41      o0777(.An(ori_ori_n763_), .B(ori_ori_n805_), .C(ori_ori_n795_), .D(ori_ori_n785_), .Y(ori_ori_n806_));
  OR2        o0778(.A(ori_ori_n721_), .B(ori_ori_n236_), .Y(ori_ori_n807_));
  NO3        o0779(.A(ori_ori_n350_), .B(ori_ori_n304_), .C(ori_ori_n112_), .Y(ori_ori_n808_));
  NA2        o0780(.A(ori_ori_n808_), .B(ori_ori_n772_), .Y(ori_ori_n809_));
  NA2        o0781(.A(ori_ori_n46_), .B(ori_ori_n56_), .Y(ori_ori_n810_));
  NO3        o0782(.A(ori_ori_n810_), .B(ori_ori_n761_), .C(ori_ori_n280_), .Y(ori_ori_n811_));
  NO3        o0783(.A(ori_ori_n536_), .B(ori_ori_n94_), .C(h), .Y(ori_ori_n812_));
  AOI210     o0784(.A0(ori_ori_n812_), .A1(ori_ori_n716_), .B0(ori_ori_n811_), .Y(ori_ori_n813_));
  NA4        o0785(.A(ori_ori_n813_), .B(ori_ori_n809_), .C(ori_ori_n807_), .D(ori_ori_n417_), .Y(ori_ori_n814_));
  OR2        o0786(.A(ori_ori_n671_), .B(ori_ori_n92_), .Y(ori_ori_n815_));
  NOi31      o0787(.An(b), .B(d), .C(a), .Y(ori_ori_n816_));
  NO2        o0788(.A(ori_ori_n816_), .B(ori_ori_n609_), .Y(ori_ori_n817_));
  NO2        o0789(.A(ori_ori_n817_), .B(n), .Y(ori_ori_n818_));
  NOi21      o0790(.An(ori_ori_n801_), .B(ori_ori_n818_), .Y(ori_ori_n819_));
  OAI220     o0791(.A0(ori_ori_n819_), .A1(ori_ori_n815_), .B0(ori_ori_n791_), .B1(ori_ori_n610_), .Y(ori_ori_n820_));
  NO2        o0792(.A(ori_ori_n564_), .B(ori_ori_n84_), .Y(ori_ori_n821_));
  NO3        o0793(.A(ori_ori_n630_), .B(ori_ori_n335_), .C(ori_ori_n116_), .Y(ori_ori_n822_));
  NOi21      o0794(.An(ori_ori_n822_), .B(ori_ori_n162_), .Y(ori_ori_n823_));
  AOI210     o0795(.A0(ori_ori_n808_), .A1(ori_ori_n821_), .B0(ori_ori_n823_), .Y(ori_ori_n824_));
  OAI210     o0796(.A0(ori_ori_n721_), .A1(ori_ori_n406_), .B0(ori_ori_n824_), .Y(ori_ori_n825_));
  NO2        o0797(.A(ori_ori_n701_), .B(n), .Y(ori_ori_n826_));
  AOI220     o0798(.A0(ori_ori_n778_), .A1(ori_ori_n678_), .B0(ori_ori_n826_), .B1(ori_ori_n711_), .Y(ori_ori_n827_));
  NO2        o0799(.A(ori_ori_n330_), .B(ori_ori_n241_), .Y(ori_ori_n828_));
  OAI210     o0800(.A0(ori_ori_n96_), .A1(ori_ori_n93_), .B0(ori_ori_n828_), .Y(ori_ori_n829_));
  NA2        o0801(.A(ori_ori_n120_), .B(ori_ori_n84_), .Y(ori_ori_n830_));
  AOI210     o0802(.A0(ori_ori_n438_), .A1(ori_ori_n430_), .B0(ori_ori_n830_), .Y(ori_ori_n831_));
  NAi21      o0803(.An(ori_ori_n831_), .B(ori_ori_n829_), .Y(ori_ori_n832_));
  NAi21      o0804(.An(ori_ori_n744_), .B(ori_ori_n448_), .Y(ori_ori_n833_));
  NO2        o0805(.A(ori_ori_n276_), .B(i), .Y(ori_ori_n834_));
  NA2        o0806(.A(ori_ori_n726_), .B(ori_ori_n358_), .Y(ori_ori_n835_));
  OAI210     o0807(.A0(ori_ori_n603_), .A1(ori_ori_n602_), .B0(ori_ori_n373_), .Y(ori_ori_n836_));
  AN3        o0808(.A(ori_ori_n836_), .B(ori_ori_n835_), .C(ori_ori_n833_), .Y(ori_ori_n837_));
  NAi31      o0809(.An(ori_ori_n832_), .B(ori_ori_n837_), .C(ori_ori_n827_), .Y(ori_ori_n838_));
  NO4        o0810(.A(ori_ori_n838_), .B(ori_ori_n825_), .C(ori_ori_n820_), .D(ori_ori_n814_), .Y(ori_ori_n839_));
  NA4        o0811(.A(ori_ori_n839_), .B(ori_ori_n806_), .C(ori_ori_n758_), .D(ori_ori_n747_), .Y(ori09));
  INV        o0812(.A(ori_ori_n121_), .Y(ori_ori_n841_));
  NA2        o0813(.A(f), .B(e), .Y(ori_ori_n842_));
  NO2        o0814(.A(ori_ori_n229_), .B(ori_ori_n112_), .Y(ori_ori_n843_));
  NA2        o0815(.A(ori_ori_n843_), .B(o), .Y(ori_ori_n844_));
  NA4        o0816(.A(ori_ori_n316_), .B(ori_ori_n483_), .C(ori_ori_n266_), .D(ori_ori_n118_), .Y(ori_ori_n845_));
  AOI210     o0817(.A0(ori_ori_n845_), .A1(o), .B0(ori_ori_n480_), .Y(ori_ori_n846_));
  AOI210     o0818(.A0(ori_ori_n846_), .A1(ori_ori_n844_), .B0(ori_ori_n842_), .Y(ori_ori_n847_));
  NA2        o0819(.A(ori_ori_n454_), .B(e), .Y(ori_ori_n848_));
  NO2        o0820(.A(ori_ori_n848_), .B(ori_ori_n523_), .Y(ori_ori_n849_));
  AOI210     o0821(.A0(ori_ori_n847_), .A1(ori_ori_n841_), .B0(ori_ori_n849_), .Y(ori_ori_n850_));
  NA3        o0822(.A(m), .B(l), .C(i), .Y(ori_ori_n851_));
  OAI220     o0823(.A0(ori_ori_n598_), .A1(ori_ori_n851_), .B0(ori_ori_n363_), .B1(ori_ori_n537_), .Y(ori_ori_n852_));
  NA4        o0824(.A(ori_ori_n88_), .B(ori_ori_n87_), .C(o), .D(f), .Y(ori_ori_n853_));
  NAi31      o0825(.An(ori_ori_n852_), .B(ori_ori_n853_), .C(ori_ori_n451_), .Y(ori_ori_n854_));
  NA3        o0826(.A(ori_ori_n815_), .B(ori_ori_n576_), .C(ori_ori_n530_), .Y(ori_ori_n855_));
  OA210      o0827(.A0(ori_ori_n855_), .A1(ori_ori_n854_), .B0(ori_ori_n818_), .Y(ori_ori_n856_));
  INV        o0828(.A(ori_ori_n347_), .Y(ori_ori_n857_));
  NO2        o0829(.A(ori_ori_n126_), .B(ori_ori_n124_), .Y(ori_ori_n858_));
  NOi31      o0830(.An(k), .B(m), .C(l), .Y(ori_ori_n859_));
  NO2        o0831(.A(ori_ori_n349_), .B(ori_ori_n859_), .Y(ori_ori_n860_));
  AOI210     o0832(.A0(ori_ori_n860_), .A1(ori_ori_n858_), .B0(ori_ori_n606_), .Y(ori_ori_n861_));
  NA2        o0833(.A(ori_ori_n800_), .B(ori_ori_n340_), .Y(ori_ori_n862_));
  NA2        o0834(.A(ori_ori_n351_), .B(ori_ori_n353_), .Y(ori_ori_n863_));
  OAI210     o0835(.A0(ori_ori_n206_), .A1(ori_ori_n216_), .B0(ori_ori_n863_), .Y(ori_ori_n864_));
  AOI220     o0836(.A0(ori_ori_n864_), .A1(ori_ori_n862_), .B0(ori_ori_n861_), .B1(ori_ori_n857_), .Y(ori_ori_n865_));
  NA2        o0837(.A(ori_ori_n170_), .B(ori_ori_n114_), .Y(ori_ori_n866_));
  NA3        o0838(.A(ori_ori_n866_), .B(ori_ori_n710_), .C(ori_ori_n135_), .Y(ori_ori_n867_));
  NA3        o0839(.A(ori_ori_n867_), .B(ori_ori_n191_), .C(ori_ori_n31_), .Y(ori_ori_n868_));
  NA4        o0840(.A(ori_ori_n868_), .B(ori_ori_n865_), .C(ori_ori_n632_), .D(ori_ori_n82_), .Y(ori_ori_n869_));
  NO2        o0841(.A(ori_ori_n594_), .B(ori_ori_n508_), .Y(ori_ori_n870_));
  NOi21      o0842(.An(f), .B(d), .Y(ori_ori_n871_));
  NA2        o0843(.A(ori_ori_n871_), .B(m), .Y(ori_ori_n872_));
  NO2        o0844(.A(ori_ori_n872_), .B(ori_ori_n52_), .Y(ori_ori_n873_));
  NOi32      o0845(.An(o), .Bn(f), .C(d), .Y(ori_ori_n874_));
  NA4        o0846(.A(ori_ori_n874_), .B(ori_ori_n611_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n875_));
  NOi21      o0847(.An(ori_ori_n317_), .B(ori_ori_n875_), .Y(ori_ori_n876_));
  AOI210     o0848(.A0(ori_ori_n873_), .A1(ori_ori_n554_), .B0(ori_ori_n876_), .Y(ori_ori_n877_));
  NA2        o0849(.A(ori_ori_n266_), .B(ori_ori_n118_), .Y(ori_ori_n878_));
  AN2        o0850(.A(f), .B(d), .Y(ori_ori_n879_));
  NA3        o0851(.A(ori_ori_n488_), .B(ori_ori_n879_), .C(ori_ori_n84_), .Y(ori_ori_n880_));
  NO3        o0852(.A(ori_ori_n880_), .B(ori_ori_n73_), .C(ori_ori_n217_), .Y(ori_ori_n881_));
  NO2        o0853(.A(ori_ori_n288_), .B(ori_ori_n56_), .Y(ori_ori_n882_));
  NA2        o0854(.A(ori_ori_n878_), .B(ori_ori_n881_), .Y(ori_ori_n883_));
  NAi31      o0855(.An(ori_ori_n500_), .B(ori_ori_n883_), .C(ori_ori_n877_), .Y(ori_ori_n884_));
  NO4        o0856(.A(ori_ori_n630_), .B(ori_ori_n131_), .C(ori_ori_n335_), .D(ori_ori_n153_), .Y(ori_ori_n885_));
  NO2        o0857(.A(ori_ori_n664_), .B(ori_ori_n335_), .Y(ori_ori_n886_));
  NO2        o0858(.A(ori_ori_n885_), .B(ori_ori_n238_), .Y(ori_ori_n887_));
  NA2        o0859(.A(ori_ori_n609_), .B(ori_ori_n84_), .Y(ori_ori_n888_));
  NO2        o0860(.A(ori_ori_n863_), .B(ori_ori_n888_), .Y(ori_ori_n889_));
  NA3        o0861(.A(ori_ori_n161_), .B(ori_ori_n109_), .C(ori_ori_n108_), .Y(ori_ori_n890_));
  OAI220     o0862(.A0(ori_ori_n880_), .A1(ori_ori_n442_), .B0(ori_ori_n347_), .B1(ori_ori_n890_), .Y(ori_ori_n891_));
  NOi41      o0863(.An(ori_ori_n227_), .B(ori_ori_n891_), .C(ori_ori_n889_), .D(ori_ori_n311_), .Y(ori_ori_n892_));
  NA2        o0864(.A(c), .B(ori_ori_n115_), .Y(ori_ori_n893_));
  NO2        o0865(.A(ori_ori_n893_), .B(ori_ori_n421_), .Y(ori_ori_n894_));
  NA3        o0866(.A(ori_ori_n894_), .B(ori_ori_n521_), .C(f), .Y(ori_ori_n895_));
  OR2        o0867(.A(ori_ori_n671_), .B(ori_ori_n550_), .Y(ori_ori_n896_));
  INV        o0868(.A(ori_ori_n896_), .Y(ori_ori_n897_));
  NA2        o0869(.A(ori_ori_n817_), .B(ori_ori_n111_), .Y(ori_ori_n898_));
  NA2        o0870(.A(ori_ori_n898_), .B(ori_ori_n897_), .Y(ori_ori_n899_));
  NA4        o0871(.A(ori_ori_n899_), .B(ori_ori_n895_), .C(ori_ori_n892_), .D(ori_ori_n887_), .Y(ori_ori_n900_));
  NO4        o0872(.A(ori_ori_n900_), .B(ori_ori_n884_), .C(ori_ori_n869_), .D(ori_ori_n856_), .Y(ori_ori_n901_));
  NA2        o0873(.A(ori_ori_n112_), .B(j), .Y(ori_ori_n902_));
  NO2        o0874(.A(ori_ori_n340_), .B(ori_ori_n853_), .Y(ori_ori_n903_));
  NO2        o0875(.A(ori_ori_n234_), .B(ori_ori_n228_), .Y(ori_ori_n904_));
  NA2        o0876(.A(ori_ori_n904_), .B(ori_ori_n231_), .Y(ori_ori_n905_));
  NO2        o0877(.A(ori_ori_n442_), .B(ori_ori_n842_), .Y(ori_ori_n906_));
  NA2        o0878(.A(ori_ori_n906_), .B(ori_ori_n571_), .Y(ori_ori_n907_));
  NA2        o0879(.A(ori_ori_n907_), .B(ori_ori_n905_), .Y(ori_ori_n908_));
  NA2        o0880(.A(e), .B(d), .Y(ori_ori_n909_));
  OAI220     o0881(.A0(ori_ori_n909_), .A1(c), .B0(ori_ori_n330_), .B1(d), .Y(ori_ori_n910_));
  NA3        o0882(.A(ori_ori_n910_), .B(ori_ori_n463_), .C(ori_ori_n519_), .Y(ori_ori_n911_));
  AOI210     o0883(.A0(ori_ori_n526_), .A1(ori_ori_n182_), .B0(ori_ori_n234_), .Y(ori_ori_n912_));
  AOI210     o0884(.A0(ori_ori_n631_), .A1(ori_ori_n356_), .B0(ori_ori_n912_), .Y(ori_ori_n913_));
  NA2        o0885(.A(ori_ori_n288_), .B(ori_ori_n166_), .Y(ori_ori_n914_));
  NA2        o0886(.A(ori_ori_n881_), .B(ori_ori_n914_), .Y(ori_ori_n915_));
  NA3        o0887(.A(ori_ori_n169_), .B(ori_ori_n85_), .C(ori_ori_n34_), .Y(ori_ori_n916_));
  NA4        o0888(.A(ori_ori_n916_), .B(ori_ori_n915_), .C(ori_ori_n913_), .D(ori_ori_n911_), .Y(ori_ori_n917_));
  NO3        o0889(.A(ori_ori_n917_), .B(ori_ori_n908_), .C(ori_ori_n903_), .Y(ori_ori_n918_));
  OR2        o0890(.A(ori_ori_n712_), .B(ori_ori_n220_), .Y(ori_ori_n919_));
  OAI220     o0891(.A0(ori_ori_n630_), .A1(ori_ori_n61_), .B0(ori_ori_n304_), .B1(j), .Y(ori_ori_n920_));
  AOI220     o0892(.A0(ori_ori_n920_), .A1(ori_ori_n886_), .B0(ori_ori_n621_), .B1(ori_ori_n629_), .Y(ori_ori_n921_));
  OAI210     o0893(.A0(ori_ori_n848_), .A1(ori_ori_n172_), .B0(ori_ori_n921_), .Y(ori_ori_n922_));
  OAI210     o0894(.A0(ori_ori_n843_), .A1(ori_ori_n914_), .B0(ori_ori_n874_), .Y(ori_ori_n923_));
  NO2        o0895(.A(ori_ori_n923_), .B(ori_ori_n612_), .Y(ori_ori_n924_));
  AOI210     o0896(.A0(ori_ori_n117_), .A1(ori_ori_n116_), .B0(ori_ori_n265_), .Y(ori_ori_n925_));
  NO2        o0897(.A(ori_ori_n925_), .B(ori_ori_n875_), .Y(ori_ori_n926_));
  AO210      o0898(.A0(ori_ori_n862_), .A1(ori_ori_n852_), .B0(ori_ori_n926_), .Y(ori_ori_n927_));
  NOi31      o0899(.An(ori_ori_n554_), .B(ori_ori_n872_), .C(ori_ori_n296_), .Y(ori_ori_n928_));
  NO4        o0900(.A(ori_ori_n928_), .B(ori_ori_n927_), .C(ori_ori_n924_), .D(ori_ori_n922_), .Y(ori_ori_n929_));
  AO220      o0901(.A0(ori_ori_n463_), .A1(ori_ori_n753_), .B0(ori_ori_n177_), .B1(f), .Y(ori_ori_n930_));
  OAI210     o0902(.A0(ori_ori_n930_), .A1(ori_ori_n466_), .B0(ori_ori_n910_), .Y(ori_ori_n931_));
  NO2        o0903(.A(ori_ori_n450_), .B(ori_ori_n70_), .Y(ori_ori_n932_));
  OAI210     o0904(.A0(ori_ori_n855_), .A1(ori_ori_n932_), .B0(ori_ori_n716_), .Y(ori_ori_n933_));
  AN4        o0905(.A(ori_ori_n933_), .B(ori_ori_n931_), .C(ori_ori_n929_), .D(ori_ori_n919_), .Y(ori_ori_n934_));
  NA4        o0906(.A(ori_ori_n934_), .B(ori_ori_n918_), .C(ori_ori_n901_), .D(ori_ori_n850_), .Y(ori12));
  NO2        o0907(.A(ori_ori_n461_), .B(c), .Y(ori_ori_n936_));
  NO4        o0908(.A(ori_ori_n453_), .B(ori_ori_n257_), .C(ori_ori_n591_), .D(ori_ori_n217_), .Y(ori_ori_n937_));
  NA2        o0909(.A(ori_ori_n937_), .B(ori_ori_n936_), .Y(ori_ori_n938_));
  NA2        o0910(.A(ori_ori_n554_), .B(ori_ori_n932_), .Y(ori_ori_n939_));
  NO2        o0911(.A(ori_ori_n461_), .B(ori_ori_n115_), .Y(ori_ori_n940_));
  NO2        o0912(.A(ori_ori_n858_), .B(ori_ori_n363_), .Y(ori_ori_n941_));
  NO2        o0913(.A(ori_ori_n671_), .B(ori_ori_n390_), .Y(ori_ori_n942_));
  AOI220     o0914(.A0(ori_ori_n942_), .A1(ori_ori_n552_), .B0(ori_ori_n941_), .B1(ori_ori_n940_), .Y(ori_ori_n943_));
  NA4        o0915(.A(ori_ori_n943_), .B(ori_ori_n939_), .C(ori_ori_n938_), .D(ori_ori_n452_), .Y(ori_ori_n944_));
  AOI210     o0916(.A0(ori_ori_n237_), .A1(ori_ori_n346_), .B0(ori_ori_n203_), .Y(ori_ori_n945_));
  OR2        o0917(.A(ori_ori_n945_), .B(ori_ori_n937_), .Y(ori_ori_n946_));
  AOI210     o0918(.A0(ori_ori_n343_), .A1(ori_ori_n402_), .B0(ori_ori_n217_), .Y(ori_ori_n947_));
  OAI210     o0919(.A0(ori_ori_n947_), .A1(ori_ori_n946_), .B0(ori_ori_n416_), .Y(ori_ori_n948_));
  NO2        o0920(.A(ori_ori_n650_), .B(ori_ori_n267_), .Y(ori_ori_n949_));
  NO2        o0921(.A(ori_ori_n598_), .B(ori_ori_n851_), .Y(ori_ori_n950_));
  NO2        o0922(.A(ori_ori_n152_), .B(ori_ori_n241_), .Y(ori_ori_n951_));
  NA3        o0923(.A(ori_ori_n951_), .B(ori_ori_n244_), .C(i), .Y(ori_ori_n952_));
  NA2        o0924(.A(ori_ori_n952_), .B(ori_ori_n948_), .Y(ori_ori_n953_));
  OR2        o0925(.A(ori_ori_n331_), .B(ori_ori_n940_), .Y(ori_ori_n954_));
  NA2        o0926(.A(ori_ori_n954_), .B(ori_ori_n364_), .Y(ori_ori_n955_));
  NA4        o0927(.A(ori_ori_n454_), .B(ori_ori_n449_), .C(ori_ori_n183_), .D(o), .Y(ori_ori_n956_));
  NA2        o0928(.A(ori_ori_n956_), .B(ori_ori_n955_), .Y(ori_ori_n957_));
  NO3        o0929(.A(ori_ori_n676_), .B(ori_ori_n92_), .C(ori_ori_n45_), .Y(ori_ori_n958_));
  NO4        o0930(.A(ori_ori_n958_), .B(ori_ori_n957_), .C(ori_ori_n953_), .D(ori_ori_n944_), .Y(ori_ori_n959_));
  NO2        o0931(.A(ori_ori_n380_), .B(ori_ori_n379_), .Y(ori_ori_n960_));
  INV        o0932(.A(ori_ori_n72_), .Y(ori_ori_n961_));
  NA2        o0933(.A(ori_ori_n564_), .B(ori_ori_n145_), .Y(ori_ori_n962_));
  NOi21      o0934(.An(ori_ori_n34_), .B(ori_ori_n664_), .Y(ori_ori_n963_));
  AOI220     o0935(.A0(ori_ori_n963_), .A1(ori_ori_n962_), .B0(ori_ori_n961_), .B1(ori_ori_n960_), .Y(ori_ori_n964_));
  OAI210     o0936(.A0(ori_ori_n255_), .A1(ori_ori_n45_), .B0(ori_ori_n964_), .Y(ori_ori_n965_));
  NA2        o0937(.A(ori_ori_n448_), .B(ori_ori_n269_), .Y(ori_ori_n966_));
  NA2        o0938(.A(ori_ori_n966_), .B(ori_ori_n327_), .Y(ori_ori_n967_));
  NO2        o0939(.A(ori_ori_n49_), .B(ori_ori_n45_), .Y(ori_ori_n968_));
  NO2        o0940(.A(ori_ori_n515_), .B(ori_ori_n304_), .Y(ori_ori_n969_));
  INV        o0941(.A(ori_ori_n969_), .Y(ori_ori_n970_));
  NO2        o0942(.A(ori_ori_n970_), .B(ori_ori_n145_), .Y(ori_ori_n971_));
  INV        o0943(.A(ori_ori_n377_), .Y(ori_ori_n972_));
  NO4        o0944(.A(ori_ori_n972_), .B(ori_ori_n971_), .C(ori_ori_n967_), .D(ori_ori_n965_), .Y(ori_ori_n973_));
  NA2        o0945(.A(ori_ori_n356_), .B(o), .Y(ori_ori_n974_));
  NA2        o0946(.A(ori_ori_n164_), .B(i), .Y(ori_ori_n975_));
  NA2        o0947(.A(ori_ori_n46_), .B(i), .Y(ori_ori_n976_));
  OAI220     o0948(.A0(ori_ori_n976_), .A1(ori_ori_n202_), .B0(ori_ori_n975_), .B1(ori_ori_n92_), .Y(ori_ori_n977_));
  AOI210     o0949(.A0(ori_ori_n432_), .A1(ori_ori_n37_), .B0(ori_ori_n977_), .Y(ori_ori_n978_));
  NO2        o0950(.A(ori_ori_n145_), .B(ori_ori_n84_), .Y(ori_ori_n979_));
  OR2        o0951(.A(ori_ori_n979_), .B(ori_ori_n563_), .Y(ori_ori_n980_));
  NA2        o0952(.A(ori_ori_n564_), .B(ori_ori_n394_), .Y(ori_ori_n981_));
  AOI210     o0953(.A0(ori_ori_n981_), .A1(n), .B0(ori_ori_n980_), .Y(ori_ori_n982_));
  OAI220     o0954(.A0(ori_ori_n982_), .A1(ori_ori_n974_), .B0(ori_ori_n978_), .B1(ori_ori_n340_), .Y(ori_ori_n983_));
  NO2        o0955(.A(ori_ori_n671_), .B(ori_ori_n508_), .Y(ori_ori_n984_));
  NA3        o0956(.A(ori_ori_n351_), .B(ori_ori_n636_), .C(i), .Y(ori_ori_n985_));
  OAI210     o0957(.A0(ori_ori_n450_), .A1(ori_ori_n316_), .B0(ori_ori_n985_), .Y(ori_ori_n986_));
  OAI220     o0958(.A0(ori_ori_n986_), .A1(ori_ori_n984_), .B0(ori_ori_n690_), .B1(ori_ori_n765_), .Y(ori_ori_n987_));
  NA2        o0959(.A(ori_ori_n615_), .B(ori_ori_n113_), .Y(ori_ori_n988_));
  OR3        o0960(.A(ori_ori_n316_), .B(ori_ori_n447_), .C(f), .Y(ori_ori_n989_));
  NA3        o0961(.A(ori_ori_n636_), .B(ori_ori_n80_), .C(i), .Y(ori_ori_n990_));
  OA220      o0962(.A0(ori_ori_n990_), .A1(ori_ori_n988_), .B0(ori_ori_n989_), .B1(ori_ori_n597_), .Y(ori_ori_n991_));
  NA3        o0963(.A(ori_ori_n332_), .B(ori_ori_n117_), .C(o), .Y(ori_ori_n992_));
  AOI210     o0964(.A0(ori_ori_n687_), .A1(ori_ori_n992_), .B0(m), .Y(ori_ori_n993_));
  OAI210     o0965(.A0(ori_ori_n993_), .A1(ori_ori_n941_), .B0(ori_ori_n331_), .Y(ori_ori_n994_));
  NA2        o0966(.A(ori_ori_n705_), .B(ori_ori_n888_), .Y(ori_ori_n995_));
  NA2        o0967(.A(ori_ori_n853_), .B(ori_ori_n451_), .Y(ori_ori_n996_));
  NA2        o0968(.A(ori_ori_n225_), .B(ori_ori_n77_), .Y(ori_ori_n997_));
  NA2        o0969(.A(ori_ori_n997_), .B(ori_ori_n990_), .Y(ori_ori_n998_));
  AOI220     o0970(.A0(ori_ori_n998_), .A1(ori_ori_n263_), .B0(ori_ori_n996_), .B1(ori_ori_n995_), .Y(ori_ori_n999_));
  NA4        o0971(.A(ori_ori_n999_), .B(ori_ori_n994_), .C(ori_ori_n991_), .D(ori_ori_n987_), .Y(ori_ori_n1000_));
  NO2        o0972(.A(ori_ori_n390_), .B(ori_ori_n91_), .Y(ori_ori_n1001_));
  OAI210     o0973(.A0(ori_ori_n1001_), .A1(ori_ori_n949_), .B0(ori_ori_n242_), .Y(ori_ori_n1002_));
  NA2        o0974(.A(ori_ori_n675_), .B(ori_ori_n88_), .Y(ori_ori_n1003_));
  NO2        o0975(.A(ori_ori_n469_), .B(ori_ori_n217_), .Y(ori_ori_n1004_));
  AOI220     o0976(.A0(ori_ori_n1004_), .A1(ori_ori_n395_), .B0(ori_ori_n954_), .B1(ori_ori_n221_), .Y(ori_ori_n1005_));
  AOI220     o0977(.A0(ori_ori_n942_), .A1(ori_ori_n951_), .B0(ori_ori_n596_), .B1(ori_ori_n90_), .Y(ori_ori_n1006_));
  NA4        o0978(.A(ori_ori_n1006_), .B(ori_ori_n1005_), .C(ori_ori_n1003_), .D(ori_ori_n1002_), .Y(ori_ori_n1007_));
  OAI210     o0979(.A0(ori_ori_n996_), .A1(ori_ori_n950_), .B0(ori_ori_n552_), .Y(ori_ori_n1008_));
  AOI210     o0980(.A0(ori_ori_n433_), .A1(ori_ori_n425_), .B0(ori_ori_n830_), .Y(ori_ori_n1009_));
  INV        o0981(.A(ori_ori_n1009_), .Y(ori_ori_n1010_));
  NA2        o0982(.A(ori_ori_n993_), .B(ori_ori_n940_), .Y(ori_ori_n1011_));
  NO3        o0983(.A(ori_ori_n902_), .B(ori_ori_n49_), .C(ori_ori_n45_), .Y(ori_ori_n1012_));
  AOI220     o0984(.A0(ori_ori_n1012_), .A1(ori_ori_n634_), .B0(ori_ori_n655_), .B1(ori_ori_n541_), .Y(ori_ori_n1013_));
  NA4        o0985(.A(ori_ori_n1013_), .B(ori_ori_n1011_), .C(ori_ori_n1010_), .D(ori_ori_n1008_), .Y(ori_ori_n1014_));
  NO4        o0986(.A(ori_ori_n1014_), .B(ori_ori_n1007_), .C(ori_ori_n1000_), .D(ori_ori_n983_), .Y(ori_ori_n1015_));
  NAi31      o0987(.An(ori_ori_n141_), .B(ori_ori_n434_), .C(n), .Y(ori_ori_n1016_));
  NO3        o0988(.A(ori_ori_n124_), .B(ori_ori_n349_), .C(ori_ori_n859_), .Y(ori_ori_n1017_));
  NO2        o0989(.A(ori_ori_n1017_), .B(ori_ori_n1016_), .Y(ori_ori_n1018_));
  NO3        o0990(.A(ori_ori_n276_), .B(ori_ori_n141_), .C(ori_ori_n421_), .Y(ori_ori_n1019_));
  AOI210     o0991(.A0(ori_ori_n1019_), .A1(ori_ori_n509_), .B0(ori_ori_n1018_), .Y(ori_ori_n1020_));
  INV        o0992(.A(ori_ori_n1020_), .Y(ori_ori_n1021_));
  NA2        o0993(.A(ori_ori_n234_), .B(ori_ori_n173_), .Y(ori_ori_n1022_));
  NO3        o0994(.A(ori_ori_n313_), .B(ori_ori_n454_), .C(ori_ori_n177_), .Y(ori_ori_n1023_));
  NOi31      o0995(.An(ori_ori_n1022_), .B(ori_ori_n1023_), .C(ori_ori_n217_), .Y(ori_ori_n1024_));
  NAi21      o0996(.An(ori_ori_n564_), .B(ori_ori_n1004_), .Y(ori_ori_n1025_));
  NA2        o0997(.A(ori_ori_n492_), .B(o), .Y(ori_ori_n1026_));
  NA2        o0998(.A(ori_ori_n1026_), .B(ori_ori_n1025_), .Y(ori_ori_n1027_));
  OAI220     o0999(.A0(ori_ori_n1016_), .A1(ori_ori_n237_), .B0(ori_ori_n985_), .B1(ori_ori_n610_), .Y(ori_ori_n1028_));
  NO2        o1000(.A(ori_ori_n672_), .B(ori_ori_n390_), .Y(ori_ori_n1029_));
  NA2        o1001(.A(ori_ori_n945_), .B(ori_ori_n936_), .Y(ori_ori_n1030_));
  OAI220     o1002(.A0(ori_ori_n942_), .A1(ori_ori_n950_), .B0(ori_ori_n554_), .B1(ori_ori_n441_), .Y(ori_ori_n1031_));
  NA3        o1003(.A(ori_ori_n1031_), .B(ori_ori_n1030_), .C(ori_ori_n628_), .Y(ori_ori_n1032_));
  OAI210     o1004(.A0(ori_ori_n945_), .A1(ori_ori_n937_), .B0(ori_ori_n1022_), .Y(ori_ori_n1033_));
  NA3        o1005(.A(ori_ori_n981_), .B(ori_ori_n497_), .C(ori_ori_n46_), .Y(ori_ori_n1034_));
  AOI210     o1006(.A0(ori_ori_n393_), .A1(ori_ori_n391_), .B0(ori_ori_n339_), .Y(ori_ori_n1035_));
  NA4        o1007(.A(ori_ori_n1035_), .B(ori_ori_n1034_), .C(ori_ori_n1033_), .D(ori_ori_n277_), .Y(ori_ori_n1036_));
  OR4        o1008(.A(ori_ori_n1036_), .B(ori_ori_n1032_), .C(ori_ori_n1029_), .D(ori_ori_n1028_), .Y(ori_ori_n1037_));
  NO4        o1009(.A(ori_ori_n1037_), .B(ori_ori_n1027_), .C(ori_ori_n1024_), .D(ori_ori_n1021_), .Y(ori_ori_n1038_));
  NA4        o1010(.A(ori_ori_n1038_), .B(ori_ori_n1015_), .C(ori_ori_n973_), .D(ori_ori_n959_), .Y(ori13));
  AN2        o1011(.A(c), .B(b), .Y(ori_ori_n1040_));
  NAi32      o1012(.An(d), .Bn(c), .C(e), .Y(ori_ori_n1041_));
  NA2        o1013(.A(ori_ori_n140_), .B(ori_ori_n45_), .Y(ori_ori_n1042_));
  NA2        o1014(.A(ori_ori_n424_), .B(ori_ori_n216_), .Y(ori_ori_n1043_));
  AN2        o1015(.A(d), .B(c), .Y(ori_ori_n1044_));
  NA2        o1016(.A(ori_ori_n1044_), .B(ori_ori_n115_), .Y(ori_ori_n1045_));
  NA2        o1017(.A(ori_ori_n506_), .B(c), .Y(ori_ori_n1046_));
  NO4        o1018(.A(ori_ori_n1042_), .B(ori_ori_n594_), .C(ori_ori_n1046_), .D(ori_ori_n312_), .Y(ori_ori_n1047_));
  NAi32      o1019(.An(f), .Bn(e), .C(c), .Y(ori_ori_n1048_));
  NO2        o1020(.A(ori_ori_n1046_), .B(ori_ori_n312_), .Y(ori_ori_n1049_));
  NO2        o1021(.A(j), .B(ori_ori_n45_), .Y(ori_ori_n1050_));
  NA2        o1022(.A(ori_ori_n638_), .B(ori_ori_n1050_), .Y(ori_ori_n1051_));
  NOi21      o1023(.An(ori_ori_n1049_), .B(ori_ori_n1051_), .Y(ori_ori_n1052_));
  NO2        o1024(.A(ori_ori_n769_), .B(ori_ori_n112_), .Y(ori_ori_n1053_));
  NOi41      o1025(.An(n), .B(m), .C(i), .D(h), .Y(ori_ori_n1054_));
  NA3        o1026(.A(k), .B(j), .C(i), .Y(ori_ori_n1055_));
  NA3        o1027(.A(ori_ori_n477_), .B(ori_ori_n342_), .C(ori_ori_n56_), .Y(ori_ori_n1056_));
  NO2        o1028(.A(ori_ori_n1056_), .B(ori_ori_n1051_), .Y(ori_ori_n1057_));
  NO4        o1029(.A(ori_ori_n1056_), .B(ori_ori_n594_), .C(ori_ori_n460_), .D(ori_ori_n45_), .Y(ori_ori_n1058_));
  NO2        o1030(.A(f), .B(c), .Y(ori_ori_n1059_));
  NOi21      o1031(.An(ori_ori_n1059_), .B(ori_ori_n453_), .Y(ori_ori_n1060_));
  OR2        o1032(.A(ori_ori_n1058_), .B(ori_ori_n1057_), .Y(ori_ori_n1061_));
  OR3        o1033(.A(ori_ori_n1061_), .B(ori_ori_n1052_), .C(ori_ori_n1047_), .Y(ori02));
  OR3        o1034(.A(n), .B(m), .C(i), .Y(ori_ori_n1063_));
  NOi31      o1035(.An(e), .B(d), .C(c), .Y(ori_ori_n1064_));
  AN3        o1036(.A(o), .B(f), .C(c), .Y(ori_ori_n1065_));
  NA3        o1037(.A(ori_ori_n1065_), .B(ori_ori_n477_), .C(h), .Y(ori_ori_n1066_));
  OR2        o1038(.A(ori_ori_n1055_), .B(ori_ori_n312_), .Y(ori_ori_n1067_));
  OR2        o1039(.A(ori_ori_n1067_), .B(ori_ori_n1066_), .Y(ori_ori_n1068_));
  NO3        o1040(.A(ori_ori_n1056_), .B(ori_ori_n1042_), .C(ori_ori_n594_), .Y(ori_ori_n1069_));
  INV        o1041(.A(ori_ori_n1069_), .Y(ori_ori_n1070_));
  NA3        o1042(.A(l), .B(k), .C(j), .Y(ori_ori_n1071_));
  NA2        o1043(.A(i), .B(h), .Y(ori_ori_n1072_));
  NO3        o1044(.A(ori_ori_n1072_), .B(ori_ori_n1071_), .C(ori_ori_n131_), .Y(ori_ori_n1073_));
  NO3        o1045(.A(ori_ori_n142_), .B(ori_ori_n286_), .C(ori_ori_n217_), .Y(ori_ori_n1074_));
  AOI210     o1046(.A0(ori_ori_n1074_), .A1(ori_ori_n1073_), .B0(ori_ori_n1052_), .Y(ori_ori_n1075_));
  NA3        o1047(.A(c), .B(b), .C(a), .Y(ori_ori_n1076_));
  INV        o1048(.A(ori_ori_n1057_), .Y(ori_ori_n1077_));
  AN4        o1049(.A(ori_ori_n1077_), .B(ori_ori_n1075_), .C(ori_ori_n1070_), .D(ori_ori_n1068_), .Y(ori_ori_n1078_));
  INV        o1050(.A(ori_ori_n1078_), .Y(ori03));
  NO2        o1051(.A(ori_ori_n537_), .B(ori_ori_n606_), .Y(ori_ori_n1080_));
  NA4        o1052(.A(ori_ori_n88_), .B(ori_ori_n87_), .C(o), .D(ori_ori_n216_), .Y(ori_ori_n1081_));
  NA4        o1053(.A(ori_ori_n583_), .B(m), .C(ori_ori_n112_), .D(ori_ori_n216_), .Y(ori_ori_n1082_));
  NA3        o1054(.A(ori_ori_n1082_), .B(ori_ori_n381_), .C(ori_ori_n1081_), .Y(ori_ori_n1083_));
  NO2        o1055(.A(ori_ori_n1083_), .B(ori_ori_n1080_), .Y(ori_ori_n1084_));
  NOi31      o1056(.An(ori_ori_n815_), .B(ori_ori_n864_), .C(ori_ori_n854_), .Y(ori_ori_n1085_));
  OAI220     o1057(.A0(ori_ori_n1085_), .A1(ori_ori_n705_), .B0(ori_ori_n1084_), .B1(ori_ori_n595_), .Y(ori_ori_n1086_));
  NOi31      o1058(.An(i), .B(k), .C(j), .Y(ori_ori_n1087_));
  NA4        o1059(.A(ori_ori_n1087_), .B(ori_ori_n1064_), .C(ori_ori_n351_), .D(ori_ori_n342_), .Y(ori_ori_n1088_));
  OAI210     o1060(.A0(ori_ori_n830_), .A1(ori_ori_n435_), .B0(ori_ori_n1088_), .Y(ori_ori_n1089_));
  NOi31      o1061(.An(m), .B(n), .C(f), .Y(ori_ori_n1090_));
  NA2        o1062(.A(ori_ori_n1090_), .B(ori_ori_n51_), .Y(ori_ori_n1091_));
  AN2        o1063(.A(e), .B(c), .Y(ori_ori_n1092_));
  NA2        o1064(.A(ori_ori_n1092_), .B(a), .Y(ori_ori_n1093_));
  OAI220     o1065(.A0(ori_ori_n1093_), .A1(ori_ori_n1091_), .B0(ori_ori_n896_), .B1(ori_ori_n440_), .Y(ori_ori_n1094_));
  NA2        o1066(.A(ori_ori_n519_), .B(l), .Y(ori_ori_n1095_));
  NO3        o1067(.A(ori_ori_n1094_), .B(ori_ori_n1089_), .C(ori_ori_n1009_), .Y(ori_ori_n1096_));
  NO2        o1068(.A(ori_ori_n286_), .B(a), .Y(ori_ori_n1097_));
  NO2        o1069(.A(ori_ori_n87_), .B(o), .Y(ori_ori_n1098_));
  INV        o1070(.A(ori_ori_n1096_), .Y(ori_ori_n1099_));
  NO4        o1071(.A(ori_ori_n1099_), .B(ori_ori_n1086_), .C(ori_ori_n832_), .D(ori_ori_n573_), .Y(ori_ori_n1100_));
  NA2        o1072(.A(c), .B(b), .Y(ori_ori_n1101_));
  NO2        o1073(.A(ori_ori_n715_), .B(ori_ori_n1101_), .Y(ori_ori_n1102_));
  OAI210     o1074(.A0(ori_ori_n872_), .A1(ori_ori_n846_), .B0(ori_ori_n428_), .Y(ori_ori_n1103_));
  OAI210     o1075(.A0(ori_ori_n1103_), .A1(ori_ori_n873_), .B0(ori_ori_n1102_), .Y(ori_ori_n1104_));
  NAi21      o1076(.An(ori_ori_n436_), .B(ori_ori_n1102_), .Y(ori_ori_n1105_));
  NA3        o1077(.A(ori_ori_n441_), .B(ori_ori_n569_), .C(f), .Y(ori_ori_n1106_));
  OAI210     o1078(.A0(ori_ori_n558_), .A1(ori_ori_n39_), .B0(ori_ori_n1097_), .Y(ori_ori_n1107_));
  NA3        o1079(.A(ori_ori_n1107_), .B(ori_ori_n1106_), .C(ori_ori_n1105_), .Y(ori_ori_n1108_));
  NA2        o1080(.A(ori_ori_n266_), .B(ori_ori_n118_), .Y(ori_ori_n1109_));
  OAI210     o1081(.A0(ori_ori_n1109_), .A1(ori_ori_n290_), .B0(o), .Y(ori_ori_n1110_));
  NAi21      o1082(.An(f), .B(d), .Y(ori_ori_n1111_));
  NO2        o1083(.A(ori_ori_n1111_), .B(ori_ori_n1076_), .Y(ori_ori_n1112_));
  INV        o1084(.A(ori_ori_n1112_), .Y(ori_ori_n1113_));
  AOI210     o1085(.A0(ori_ori_n1110_), .A1(ori_ori_n296_), .B0(ori_ori_n1113_), .Y(ori_ori_n1114_));
  AOI210     o1086(.A0(ori_ori_n1114_), .A1(ori_ori_n113_), .B0(ori_ori_n1108_), .Y(ori_ori_n1115_));
  NA2        o1087(.A(ori_ori_n480_), .B(ori_ori_n479_), .Y(ori_ori_n1116_));
  NO2        o1088(.A(ori_ori_n184_), .B(ori_ori_n241_), .Y(ori_ori_n1117_));
  NA2        o1089(.A(ori_ori_n1117_), .B(m), .Y(ori_ori_n1118_));
  NA3        o1090(.A(ori_ori_n925_), .B(ori_ori_n1095_), .C(ori_ori_n483_), .Y(ori_ori_n1119_));
  NA2        o1091(.A(ori_ori_n1119_), .B(ori_ori_n481_), .Y(ori_ori_n1120_));
  AOI210     o1092(.A0(ori_ori_n1120_), .A1(ori_ori_n1116_), .B0(ori_ori_n1118_), .Y(ori_ori_n1121_));
  NA2        o1093(.A(ori_ori_n571_), .B(ori_ori_n423_), .Y(ori_ori_n1122_));
  NA2        o1094(.A(ori_ori_n457_), .B(ori_ori_n1112_), .Y(ori_ori_n1123_));
  NO2        o1095(.A(ori_ori_n384_), .B(ori_ori_n383_), .Y(ori_ori_n1124_));
  NA2        o1096(.A(ori_ori_n1117_), .B(ori_ori_n443_), .Y(ori_ori_n1125_));
  NAi41      o1097(.An(ori_ori_n1124_), .B(ori_ori_n1125_), .C(ori_ori_n1123_), .D(ori_ori_n1122_), .Y(ori_ori_n1126_));
  NO2        o1098(.A(ori_ori_n1126_), .B(ori_ori_n1121_), .Y(ori_ori_n1127_));
  NA4        o1099(.A(ori_ori_n1127_), .B(ori_ori_n1115_), .C(ori_ori_n1104_), .D(ori_ori_n1100_), .Y(ori00));
  AOI210     o1100(.A0(ori_ori_n906_), .A1(ori_ori_n951_), .B0(ori_ori_n1089_), .Y(ori_ori_n1129_));
  NO2        o1101(.A(ori_ori_n1069_), .B(ori_ori_n725_), .Y(ori_ori_n1130_));
  NA3        o1102(.A(ori_ori_n1130_), .B(ori_ori_n1129_), .C(ori_ori_n1010_), .Y(ori_ori_n1131_));
  NA2        o1103(.A(ori_ori_n521_), .B(f), .Y(ori_ori_n1132_));
  OAI210     o1104(.A0(ori_ori_n1017_), .A1(ori_ori_n40_), .B0(ori_ori_n657_), .Y(ori_ori_n1133_));
  NA3        o1105(.A(ori_ori_n1133_), .B(ori_ori_n262_), .C(n), .Y(ori_ori_n1134_));
  AOI210     o1106(.A0(ori_ori_n1134_), .A1(ori_ori_n1132_), .B0(ori_ori_n1045_), .Y(ori_ori_n1135_));
  NO3        o1107(.A(ori_ori_n1135_), .B(ori_ori_n1131_), .C(ori_ori_n1052_), .Y(ori_ori_n1136_));
  NA3        o1108(.A(ori_ori_n169_), .B(ori_ori_n46_), .C(ori_ori_n45_), .Y(ori_ori_n1137_));
  NA3        o1109(.A(d), .B(ori_ori_n56_), .C(b), .Y(ori_ori_n1138_));
  NO2        o1110(.A(ori_ori_n1138_), .B(ori_ori_n1137_), .Y(ori_ori_n1139_));
  INV        o1111(.A(ori_ori_n585_), .Y(ori_ori_n1140_));
  NO4        o1112(.A(ori_ori_n1140_), .B(ori_ori_n1139_), .C(ori_ori_n1124_), .D(ori_ori_n928_), .Y(ori_ori_n1141_));
  NO4        o1113(.A(ori_ori_n498_), .B(ori_ori_n366_), .C(ori_ori_n1101_), .D(ori_ori_n59_), .Y(ori_ori_n1142_));
  NA3        o1114(.A(ori_ori_n396_), .B(ori_ori_n224_), .C(o), .Y(ori_ori_n1143_));
  OA220      o1115(.A0(ori_ori_n1143_), .A1(ori_ori_n1138_), .B0(ori_ori_n397_), .B1(ori_ori_n134_), .Y(ori_ori_n1144_));
  NO2        o1116(.A(h), .B(o), .Y(ori_ori_n1145_));
  NA4        o1117(.A(ori_ori_n509_), .B(ori_ori_n477_), .C(ori_ori_n1145_), .D(ori_ori_n1040_), .Y(ori_ori_n1146_));
  OAI220     o1118(.A0(ori_ori_n537_), .A1(ori_ori_n606_), .B0(ori_ori_n92_), .B1(ori_ori_n91_), .Y(ori_ori_n1147_));
  NA2        o1119(.A(ori_ori_n1147_), .B(ori_ori_n545_), .Y(ori_ori_n1148_));
  AOI220     o1120(.A0(ori_ori_n324_), .A1(ori_ori_n251_), .B0(ori_ori_n179_), .B1(ori_ori_n149_), .Y(ori_ori_n1149_));
  NA4        o1121(.A(ori_ori_n1149_), .B(ori_ori_n1148_), .C(ori_ori_n1146_), .D(ori_ori_n1144_), .Y(ori_ori_n1150_));
  NO3        o1122(.A(ori_ori_n1150_), .B(ori_ori_n1142_), .C(ori_ori_n270_), .Y(ori_ori_n1151_));
  INV        o1123(.A(ori_ori_n329_), .Y(ori_ori_n1152_));
  AOI210     o1124(.A0(ori_ori_n251_), .A1(ori_ori_n356_), .B0(ori_ori_n587_), .Y(ori_ori_n1153_));
  NA3        o1125(.A(ori_ori_n1153_), .B(ori_ori_n1152_), .C(ori_ori_n155_), .Y(ori_ori_n1154_));
  NO2        o1126(.A(ori_ori_n243_), .B(ori_ori_n183_), .Y(ori_ori_n1155_));
  NA2        o1127(.A(ori_ori_n1155_), .B(ori_ori_n441_), .Y(ori_ori_n1156_));
  NA3        o1128(.A(ori_ori_n181_), .B(ori_ori_n112_), .C(o), .Y(ori_ori_n1157_));
  NA3        o1129(.A(ori_ori_n477_), .B(ori_ori_n40_), .C(f), .Y(ori_ori_n1158_));
  NOi31      o1130(.An(ori_ori_n882_), .B(ori_ori_n1158_), .C(ori_ori_n1157_), .Y(ori_ori_n1159_));
  NAi31      o1131(.An(ori_ori_n187_), .B(ori_ori_n870_), .C(ori_ori_n477_), .Y(ori_ori_n1160_));
  NAi31      o1132(.An(ori_ori_n1159_), .B(ori_ori_n1160_), .C(ori_ori_n1156_), .Y(ori_ori_n1161_));
  NO4        o1133(.A(ori_ori_n1047_), .B(ori_ori_n1161_), .C(ori_ori_n1154_), .D(ori_ori_n529_), .Y(ori_ori_n1162_));
  AN3        o1134(.A(ori_ori_n1162_), .B(ori_ori_n1151_), .C(ori_ori_n1141_), .Y(ori_ori_n1163_));
  NA3        o1135(.A(ori_ori_n1090_), .B(ori_ori_n615_), .C(ori_ori_n476_), .Y(ori_ori_n1164_));
  NA3        o1136(.A(ori_ori_n1164_), .B(ori_ori_n572_), .C(ori_ori_n245_), .Y(ori_ori_n1165_));
  NA2        o1137(.A(ori_ori_n1083_), .B(ori_ori_n545_), .Y(ori_ori_n1166_));
  NA4        o1138(.A(ori_ori_n660_), .B(ori_ori_n208_), .C(ori_ori_n224_), .D(ori_ori_n164_), .Y(ori_ori_n1167_));
  NA3        o1139(.A(ori_ori_n1167_), .B(ori_ori_n1166_), .C(ori_ori_n300_), .Y(ori_ori_n1168_));
  OAI210     o1140(.A0(ori_ori_n475_), .A1(ori_ori_n119_), .B0(ori_ori_n875_), .Y(ori_ori_n1169_));
  AOI220     o1141(.A0(ori_ori_n1169_), .A1(ori_ori_n1119_), .B0(ori_ori_n571_), .B1(ori_ori_n423_), .Y(ori_ori_n1170_));
  OR4        o1142(.A(ori_ori_n1045_), .B(ori_ori_n276_), .C(ori_ori_n226_), .D(e), .Y(ori_ori_n1171_));
  NA2        o1143(.A(n), .B(e), .Y(ori_ori_n1172_));
  NO2        o1144(.A(ori_ori_n1172_), .B(ori_ori_n147_), .Y(ori_ori_n1173_));
  NA2        o1145(.A(ori_ori_n1173_), .B(ori_ori_n278_), .Y(ori_ori_n1174_));
  OAI210     o1146(.A0(ori_ori_n367_), .A1(ori_ori_n318_), .B0(ori_ori_n459_), .Y(ori_ori_n1175_));
  NA4        o1147(.A(ori_ori_n1175_), .B(ori_ori_n1174_), .C(ori_ori_n1171_), .D(ori_ori_n1170_), .Y(ori_ori_n1176_));
  AOI210     o1148(.A0(ori_ori_n1173_), .A1(ori_ori_n861_), .B0(ori_ori_n831_), .Y(ori_ori_n1177_));
  AOI220     o1149(.A0(ori_ori_n963_), .A1(ori_ori_n584_), .B0(ori_ori_n660_), .B1(ori_ori_n248_), .Y(ori_ori_n1178_));
  NO2        o1150(.A(ori_ori_n68_), .B(h), .Y(ori_ori_n1179_));
  NA3        o1151(.A(ori_ori_n1178_), .B(ori_ori_n1177_), .C(ori_ori_n877_), .Y(ori_ori_n1180_));
  NO4        o1152(.A(ori_ori_n1180_), .B(ori_ori_n1176_), .C(ori_ori_n1168_), .D(ori_ori_n1165_), .Y(ori_ori_n1181_));
  NA2        o1153(.A(ori_ori_n847_), .B(ori_ori_n764_), .Y(ori_ori_n1182_));
  NA4        o1154(.A(ori_ori_n1182_), .B(ori_ori_n1181_), .C(ori_ori_n1163_), .D(ori_ori_n1136_), .Y(ori01));
  NO3        o1155(.A(ori_ori_n811_), .B(ori_ori_n803_), .C(ori_ori_n284_), .Y(ori_ori_n1184_));
  NA2        o1156(.A(ori_ori_n407_), .B(i), .Y(ori_ori_n1185_));
  NA3        o1157(.A(ori_ori_n1185_), .B(ori_ori_n1184_), .C(ori_ori_n1030_), .Y(ori_ori_n1186_));
  NA2        o1158(.A(ori_ori_n596_), .B(ori_ori_n90_), .Y(ori_ori_n1187_));
  NA2        o1159(.A(ori_ori_n564_), .B(ori_ori_n275_), .Y(ori_ori_n1188_));
  NA2        o1160(.A(ori_ori_n969_), .B(ori_ori_n1188_), .Y(ori_ori_n1189_));
  NA4        o1161(.A(ori_ori_n1189_), .B(ori_ori_n1187_), .C(ori_ori_n921_), .D(ori_ori_n341_), .Y(ori_ori_n1190_));
  NA2        o1162(.A(ori_ori_n45_), .B(f), .Y(ori_ori_n1191_));
  NA2        o1163(.A(ori_ori_n722_), .B(ori_ori_n97_), .Y(ori_ori_n1192_));
  NO2        o1164(.A(ori_ori_n1192_), .B(ori_ori_n1191_), .Y(ori_ori_n1193_));
  OAI210     o1165(.A0(ori_ori_n791_), .A1(ori_ori_n610_), .B0(ori_ori_n1167_), .Y(ori_ori_n1194_));
  AOI210     o1166(.A0(ori_ori_n1193_), .A1(ori_ori_n645_), .B0(ori_ori_n1194_), .Y(ori_ori_n1195_));
  INV        o1167(.A(ori_ori_n117_), .Y(ori_ori_n1196_));
  OR2        o1168(.A(ori_ori_n673_), .B(ori_ori_n381_), .Y(ori_ori_n1197_));
  NAi41      o1169(.An(ori_ori_n163_), .B(ori_ori_n1197_), .C(ori_ori_n1195_), .D(ori_ori_n905_), .Y(ori_ori_n1198_));
  NO2        o1170(.A(ori_ori_n689_), .B(ori_ori_n524_), .Y(ori_ori_n1199_));
  NA4        o1171(.A(ori_ori_n722_), .B(ori_ori_n97_), .C(ori_ori_n45_), .D(ori_ori_n216_), .Y(ori_ori_n1200_));
  OA220      o1172(.A0(ori_ori_n1200_), .A1(ori_ori_n682_), .B0(ori_ori_n197_), .B1(ori_ori_n195_), .Y(ori_ori_n1201_));
  NA3        o1173(.A(ori_ori_n1201_), .B(ori_ori_n1199_), .C(ori_ori_n137_), .Y(ori_ori_n1202_));
  NO4        o1174(.A(ori_ori_n1202_), .B(ori_ori_n1198_), .C(ori_ori_n1190_), .D(ori_ori_n1186_), .Y(ori_ori_n1203_));
  INV        o1175(.A(ori_ori_n1143_), .Y(ori_ori_n1204_));
  OAI210     o1176(.A0(ori_ori_n1204_), .A1(ori_ori_n306_), .B0(ori_ori_n541_), .Y(ori_ori_n1205_));
  AOI210     o1177(.A0(ori_ori_n206_), .A1(ori_ori_n89_), .B0(ori_ori_n216_), .Y(ori_ori_n1206_));
  OAI210     o1178(.A0(ori_ori_n818_), .A1(ori_ori_n441_), .B0(ori_ori_n1206_), .Y(ori_ori_n1207_));
  AN3        o1179(.A(m), .B(l), .C(k), .Y(ori_ori_n1208_));
  OAI210     o1180(.A0(ori_ori_n369_), .A1(ori_ori_n34_), .B0(ori_ori_n1208_), .Y(ori_ori_n1209_));
  NA2        o1181(.A(ori_ori_n205_), .B(ori_ori_n34_), .Y(ori_ori_n1210_));
  AO210      o1182(.A0(ori_ori_n1210_), .A1(ori_ori_n1209_), .B0(ori_ori_n340_), .Y(ori_ori_n1211_));
  NA3        o1183(.A(ori_ori_n1211_), .B(ori_ori_n1207_), .C(ori_ori_n1205_), .Y(ori_ori_n1212_));
  AOI210     o1184(.A0(ori_ori_n604_), .A1(ori_ori_n117_), .B0(ori_ori_n608_), .Y(ori_ori_n1213_));
  OAI210     o1185(.A0(ori_ori_n1196_), .A1(ori_ori_n601_), .B0(ori_ori_n1213_), .Y(ori_ori_n1214_));
  NA2        o1186(.A(ori_ori_n283_), .B(ori_ori_n197_), .Y(ori_ori_n1215_));
  NA2        o1187(.A(ori_ori_n1215_), .B(ori_ori_n678_), .Y(ori_ori_n1216_));
  NO3        o1188(.A(ori_ori_n830_), .B(ori_ori_n206_), .C(ori_ori_n421_), .Y(ori_ori_n1217_));
  INV        o1189(.A(ori_ori_n1217_), .Y(ori_ori_n1218_));
  OAI210     o1190(.A0(ori_ori_n1193_), .A1(ori_ori_n334_), .B0(ori_ori_n690_), .Y(ori_ori_n1219_));
  NA4        o1191(.A(ori_ori_n1219_), .B(ori_ori_n1218_), .C(ori_ori_n1216_), .D(ori_ori_n794_), .Y(ori_ori_n1220_));
  NO3        o1192(.A(ori_ori_n1220_), .B(ori_ori_n1214_), .C(ori_ori_n1212_), .Y(ori_ori_n1221_));
  NA3        o1193(.A(ori_ori_n611_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n1222_));
  NO2        o1194(.A(ori_ori_n1222_), .B(ori_ori_n206_), .Y(ori_ori_n1223_));
  AOI210     o1195(.A0(ori_ori_n516_), .A1(ori_ori_n58_), .B0(ori_ori_n1223_), .Y(ori_ori_n1224_));
  OR3        o1196(.A(ori_ori_n1192_), .B(ori_ori_n612_), .C(ori_ori_n1191_), .Y(ori_ori_n1225_));
  NO2        o1197(.A(ori_ori_n1200_), .B(ori_ori_n988_), .Y(ori_ori_n1226_));
  NO2        o1198(.A(ori_ori_n209_), .B(ori_ori_n111_), .Y(ori_ori_n1227_));
  NO3        o1199(.A(ori_ori_n1227_), .B(ori_ori_n1226_), .C(ori_ori_n1139_), .Y(ori_ori_n1228_));
  NA4        o1200(.A(ori_ori_n1228_), .B(ori_ori_n1225_), .C(ori_ori_n1224_), .D(ori_ori_n763_), .Y(ori_ori_n1229_));
  NO2        o1201(.A(ori_ori_n975_), .B(ori_ori_n236_), .Y(ori_ori_n1230_));
  NO2        o1202(.A(ori_ori_n976_), .B(ori_ori_n566_), .Y(ori_ori_n1231_));
  OAI210     o1203(.A0(ori_ori_n1231_), .A1(ori_ori_n1230_), .B0(ori_ori_n349_), .Y(ori_ori_n1232_));
  NO3        o1204(.A(ori_ori_n79_), .B(ori_ori_n304_), .C(ori_ori_n45_), .Y(ori_ori_n1233_));
  NA2        o1205(.A(ori_ori_n1233_), .B(ori_ori_n563_), .Y(ori_ori_n1234_));
  NA2        o1206(.A(ori_ori_n1234_), .B(ori_ori_n684_), .Y(ori_ori_n1235_));
  OR2        o1207(.A(ori_ori_n1143_), .B(ori_ori_n1138_), .Y(ori_ori_n1236_));
  NO2        o1208(.A(ori_ori_n381_), .B(ori_ori_n72_), .Y(ori_ori_n1237_));
  INV        o1209(.A(ori_ori_n1237_), .Y(ori_ori_n1238_));
  NA2        o1210(.A(ori_ori_n1233_), .B(ori_ori_n821_), .Y(ori_ori_n1239_));
  NA4        o1211(.A(ori_ori_n1239_), .B(ori_ori_n1238_), .C(ori_ori_n1236_), .D(ori_ori_n399_), .Y(ori_ori_n1240_));
  NOi41      o1212(.An(ori_ori_n1232_), .B(ori_ori_n1240_), .C(ori_ori_n1235_), .D(ori_ori_n1229_), .Y(ori_ori_n1241_));
  NO2        o1213(.A(ori_ori_n130_), .B(ori_ori_n45_), .Y(ori_ori_n1242_));
  NO2        o1214(.A(ori_ori_n45_), .B(ori_ori_n40_), .Y(ori_ori_n1243_));
  AO220      o1215(.A0(ori_ori_n1243_), .A1(ori_ori_n631_), .B0(ori_ori_n1242_), .B1(ori_ori_n720_), .Y(ori_ori_n1244_));
  NA2        o1216(.A(ori_ori_n1244_), .B(ori_ori_n349_), .Y(ori_ori_n1245_));
  INV        o1217(.A(ori_ori_n134_), .Y(ori_ori_n1246_));
  NO3        o1218(.A(ori_ori_n1072_), .B(ori_ori_n178_), .C(ori_ori_n87_), .Y(ori_ori_n1247_));
  AOI220     o1219(.A0(ori_ori_n1247_), .A1(ori_ori_n1246_), .B0(ori_ori_n1233_), .B1(ori_ori_n979_), .Y(ori_ori_n1248_));
  NA2        o1220(.A(ori_ori_n1248_), .B(ori_ori_n1245_), .Y(ori_ori_n1249_));
  NO2        o1221(.A(ori_ori_n623_), .B(ori_ori_n622_), .Y(ori_ori_n1250_));
  NO4        o1222(.A(ori_ori_n1072_), .B(ori_ori_n1250_), .C(ori_ori_n176_), .D(ori_ori_n87_), .Y(ori_ori_n1251_));
  NO3        o1223(.A(ori_ori_n1251_), .B(ori_ori_n1249_), .C(ori_ori_n649_), .Y(ori_ori_n1252_));
  NA4        o1224(.A(ori_ori_n1252_), .B(ori_ori_n1241_), .C(ori_ori_n1221_), .D(ori_ori_n1203_), .Y(ori06));
  NO2        o1225(.A(ori_ori_n422_), .B(ori_ori_n570_), .Y(ori_ori_n1254_));
  NA2        o1226(.A(ori_ori_n271_), .B(ori_ori_n1254_), .Y(ori_ori_n1255_));
  NO2        o1227(.A(ori_ori_n228_), .B(ori_ori_n103_), .Y(ori_ori_n1256_));
  OAI210     o1228(.A0(ori_ori_n1256_), .A1(ori_ori_n1247_), .B0(ori_ori_n395_), .Y(ori_ori_n1257_));
  NO3        o1229(.A(ori_ori_n607_), .B(ori_ori_n816_), .C(ori_ori_n609_), .Y(ori_ori_n1258_));
  OR2        o1230(.A(ori_ori_n1258_), .B(ori_ori_n896_), .Y(ori_ori_n1259_));
  NA4        o1231(.A(ori_ori_n1259_), .B(ori_ori_n1257_), .C(ori_ori_n1255_), .D(ori_ori_n1232_), .Y(ori_ori_n1260_));
  NO3        o1232(.A(ori_ori_n1260_), .B(ori_ori_n1235_), .C(ori_ori_n261_), .Y(ori_ori_n1261_));
  NO2        o1233(.A(ori_ori_n304_), .B(ori_ori_n45_), .Y(ori_ori_n1262_));
  AOI210     o1234(.A0(ori_ori_n1262_), .A1(ori_ori_n980_), .B0(ori_ori_n1230_), .Y(ori_ori_n1263_));
  AOI210     o1235(.A0(ori_ori_n1262_), .A1(ori_ori_n567_), .B0(ori_ori_n1244_), .Y(ori_ori_n1264_));
  AOI210     o1236(.A0(ori_ori_n1264_), .A1(ori_ori_n1263_), .B0(ori_ori_n346_), .Y(ori_ori_n1265_));
  OAI210     o1237(.A0(ori_ori_n89_), .A1(ori_ori_n40_), .B0(ori_ori_n688_), .Y(ori_ori_n1266_));
  NA2        o1238(.A(ori_ori_n1266_), .B(ori_ori_n653_), .Y(ori_ori_n1267_));
  NO2        o1239(.A(ori_ori_n526_), .B(ori_ori_n173_), .Y(ori_ori_n1268_));
  NOi21      o1240(.An(ori_ori_n136_), .B(ori_ori_n45_), .Y(ori_ori_n1269_));
  NO2        o1241(.A(ori_ori_n616_), .B(ori_ori_n1091_), .Y(ori_ori_n1270_));
  OAI210     o1242(.A0(ori_ori_n470_), .A1(ori_ori_n252_), .B0(ori_ori_n916_), .Y(ori_ori_n1271_));
  NO4        o1243(.A(ori_ori_n1271_), .B(ori_ori_n1270_), .C(ori_ori_n1269_), .D(ori_ori_n1268_), .Y(ori_ori_n1272_));
  NO2        o1244(.A(ori_ori_n380_), .B(ori_ori_n135_), .Y(ori_ori_n1273_));
  INV        o1245(.A(ori_ori_n608_), .Y(ori_ori_n1274_));
  NA3        o1246(.A(ori_ori_n1274_), .B(ori_ori_n1272_), .C(ori_ori_n1267_), .Y(ori_ori_n1275_));
  NO2        o1247(.A(ori_ori_n754_), .B(ori_ori_n379_), .Y(ori_ori_n1276_));
  AN2        o1248(.A(ori_ori_n963_), .B(ori_ori_n656_), .Y(ori_ori_n1277_));
  NO3        o1249(.A(ori_ori_n1277_), .B(ori_ori_n1275_), .C(ori_ori_n1265_), .Y(ori_ori_n1278_));
  NO2        o1250(.A(ori_ori_n810_), .B(ori_ori_n280_), .Y(ori_ori_n1279_));
  OAI220     o1251(.A0(ori_ori_n744_), .A1(ori_ori_n47_), .B0(ori_ori_n228_), .B1(ori_ori_n625_), .Y(ori_ori_n1280_));
  AOI220     o1252(.A0(ori_ori_n372_), .A1(ori_ori_n1280_), .B0(ori_ori_n1279_), .B1(ori_ori_n271_), .Y(ori_ori_n1281_));
  NO3        o1253(.A(ori_ori_n247_), .B(ori_ori_n103_), .C(ori_ori_n286_), .Y(ori_ori_n1282_));
  OAI220     o1254(.A0(ori_ori_n712_), .A1(ori_ori_n252_), .B0(ori_ori_n523_), .B1(ori_ori_n526_), .Y(ori_ori_n1283_));
  INV        o1255(.A(k), .Y(ori_ori_n1284_));
  NO3        o1256(.A(ori_ori_n1284_), .B(ori_ori_n606_), .C(j), .Y(ori_ori_n1285_));
  NO3        o1257(.A(ori_ori_n1283_), .B(ori_ori_n1282_), .C(ori_ori_n1094_), .Y(ori_ori_n1286_));
  NA2        o1258(.A(ori_ori_n801_), .B(ori_ori_n800_), .Y(ori_ori_n1287_));
  NAi31      o1259(.An(ori_ori_n754_), .B(ori_ori_n1287_), .C(ori_ori_n205_), .Y(ori_ori_n1288_));
  NA4        o1260(.A(ori_ori_n1288_), .B(ori_ori_n1286_), .C(ori_ori_n1281_), .D(ori_ori_n1178_), .Y(ori_ori_n1289_));
  NOi31      o1261(.An(ori_ori_n1258_), .B(ori_ori_n474_), .C(ori_ori_n408_), .Y(ori_ori_n1290_));
  OR3        o1262(.A(ori_ori_n1290_), .B(ori_ori_n791_), .C(ori_ori_n550_), .Y(ori_ori_n1291_));
  AOI210     o1263(.A0(ori_ori_n579_), .A1(ori_ori_n459_), .B0(ori_ori_n385_), .Y(ori_ori_n1292_));
  NA2        o1264(.A(ori_ori_n1285_), .B(ori_ori_n797_), .Y(ori_ori_n1293_));
  NA3        o1265(.A(ori_ori_n1293_), .B(ori_ori_n1292_), .C(ori_ori_n1291_), .Y(ori_ori_n1294_));
  AOI220     o1266(.A0(ori_ori_n1276_), .A1(ori_ori_n764_), .B0(ori_ori_n1273_), .B1(ori_ori_n242_), .Y(ori_ori_n1295_));
  AN2        o1267(.A(ori_ori_n937_), .B(ori_ori_n936_), .Y(ori_ori_n1296_));
  NO3        o1268(.A(ori_ori_n1296_), .B(ori_ori_n512_), .C(ori_ori_n492_), .Y(ori_ori_n1297_));
  NA3        o1269(.A(ori_ori_n1297_), .B(ori_ori_n1295_), .C(ori_ori_n1239_), .Y(ori_ori_n1298_));
  NAi21      o1270(.An(j), .B(i), .Y(ori_ori_n1299_));
  NO4        o1271(.A(ori_ori_n1250_), .B(ori_ori_n1299_), .C(ori_ori_n453_), .D(ori_ori_n239_), .Y(ori_ori_n1300_));
  NO4        o1272(.A(ori_ori_n1300_), .B(ori_ori_n1298_), .C(ori_ori_n1294_), .D(ori_ori_n1289_), .Y(ori_ori_n1301_));
  NA4        o1273(.A(ori_ori_n1301_), .B(ori_ori_n1278_), .C(ori_ori_n1261_), .D(ori_ori_n1252_), .Y(ori07));
  NOi21      o1274(.An(j), .B(k), .Y(ori_ori_n1303_));
  NA4        o1275(.A(ori_ori_n181_), .B(ori_ori_n109_), .C(ori_ori_n1303_), .D(f), .Y(ori_ori_n1304_));
  NAi32      o1276(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1305_));
  NO3        o1277(.A(ori_ori_n1305_), .B(o), .C(f), .Y(ori_ori_n1306_));
  INV        o1278(.A(ori_ori_n1306_), .Y(ori_ori_n1307_));
  NAi21      o1279(.An(f), .B(c), .Y(ori_ori_n1308_));
  OR2        o1280(.A(e), .B(d), .Y(ori_ori_n1309_));
  NO2        o1281(.A(ori_ori_n637_), .B(ori_ori_n330_), .Y(ori_ori_n1310_));
  NA3        o1282(.A(ori_ori_n1310_), .B(ori_ori_n1050_), .C(ori_ori_n181_), .Y(ori_ori_n1311_));
  NOi31      o1283(.An(n), .B(m), .C(b), .Y(ori_ori_n1312_));
  NA3        o1284(.A(ori_ori_n1311_), .B(ori_ori_n1307_), .C(ori_ori_n1304_), .Y(ori_ori_n1313_));
  NOi41      o1285(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1314_));
  NA3        o1286(.A(ori_ori_n1314_), .B(ori_ori_n879_), .C(ori_ori_n424_), .Y(ori_ori_n1315_));
  NO2        o1287(.A(ori_ori_n1315_), .B(ori_ori_n56_), .Y(ori_ori_n1316_));
  NO2        o1288(.A(k), .B(i), .Y(ori_ori_n1317_));
  NA3        o1289(.A(ori_ori_n1317_), .B(ori_ori_n904_), .C(ori_ori_n181_), .Y(ori_ori_n1318_));
  NA2        o1290(.A(ori_ori_n87_), .B(ori_ori_n45_), .Y(ori_ori_n1319_));
  NO2        o1291(.A(ori_ori_n1048_), .B(ori_ori_n453_), .Y(ori_ori_n1320_));
  NA3        o1292(.A(ori_ori_n1320_), .B(ori_ori_n1319_), .C(ori_ori_n217_), .Y(ori_ori_n1321_));
  NO2        o1293(.A(ori_ori_n1055_), .B(ori_ori_n312_), .Y(ori_ori_n1322_));
  NA2        o1294(.A(ori_ori_n551_), .B(ori_ori_n80_), .Y(ori_ori_n1323_));
  NA2        o1295(.A(ori_ori_n1179_), .B(ori_ori_n294_), .Y(ori_ori_n1324_));
  NA4        o1296(.A(ori_ori_n1324_), .B(ori_ori_n1323_), .C(ori_ori_n1321_), .D(ori_ori_n1318_), .Y(ori_ori_n1325_));
  NO3        o1297(.A(ori_ori_n1325_), .B(ori_ori_n1316_), .C(ori_ori_n1313_), .Y(ori_ori_n1326_));
  NO3        o1298(.A(e), .B(d), .C(c), .Y(ori_ori_n1327_));
  NO2        o1299(.A(ori_ori_n131_), .B(ori_ori_n217_), .Y(ori_ori_n1328_));
  NA2        o1300(.A(ori_ori_n1328_), .B(ori_ori_n1327_), .Y(ori_ori_n1329_));
  INV        o1301(.A(ori_ori_n1329_), .Y(ori_ori_n1330_));
  OR2        o1302(.A(h), .B(f), .Y(ori_ori_n1331_));
  NO3        o1303(.A(n), .B(m), .C(i), .Y(ori_ori_n1332_));
  NA2        o1304(.A(ori_ori_n1092_), .B(ori_ori_n1332_), .Y(ori_ori_n1333_));
  NO2        o1305(.A(ori_ori_n1333_), .B(ori_ori_n1331_), .Y(ori_ori_n1334_));
  NA3        o1306(.A(ori_ori_n709_), .B(ori_ori_n697_), .C(ori_ori_n112_), .Y(ori_ori_n1335_));
  NA3        o1307(.A(ori_ori_n1312_), .B(ori_ori_n1053_), .C(ori_ori_n686_), .Y(ori_ori_n1336_));
  AOI210     o1308(.A0(ori_ori_n1336_), .A1(ori_ori_n1335_), .B0(ori_ori_n45_), .Y(ori_ori_n1337_));
  NA2        o1309(.A(ori_ori_n1332_), .B(ori_ori_n651_), .Y(ori_ori_n1338_));
  NO2        o1310(.A(l), .B(k), .Y(ori_ori_n1339_));
  NOi41      o1311(.An(ori_ori_n556_), .B(ori_ori_n1339_), .C(ori_ori_n489_), .D(ori_ori_n453_), .Y(ori_ori_n1340_));
  NO3        o1312(.A(ori_ori_n453_), .B(d), .C(c), .Y(ori_ori_n1341_));
  NO4        o1313(.A(ori_ori_n1340_), .B(ori_ori_n1337_), .C(ori_ori_n1334_), .D(ori_ori_n1330_), .Y(ori_ori_n1342_));
  NO2        o1314(.A(ori_ori_n148_), .B(h), .Y(ori_ori_n1343_));
  NO2        o1315(.A(o), .B(c), .Y(ori_ori_n1344_));
  NO2        o1316(.A(ori_ori_n461_), .B(a), .Y(ori_ori_n1345_));
  NA2        o1317(.A(ori_ori_n1345_), .B(ori_ori_n113_), .Y(ori_ori_n1346_));
  NO2        o1318(.A(i), .B(h), .Y(ori_ori_n1347_));
  NA2        o1319(.A(ori_ori_n138_), .B(ori_ori_n224_), .Y(ori_ori_n1348_));
  NO2        o1320(.A(ori_ori_n1348_), .B(ori_ori_n1478_), .Y(ori_ori_n1349_));
  NO2        o1321(.A(ori_ori_n761_), .B(ori_ori_n189_), .Y(ori_ori_n1350_));
  NOi31      o1322(.An(m), .B(n), .C(b), .Y(ori_ori_n1351_));
  NOi31      o1323(.An(f), .B(d), .C(c), .Y(ori_ori_n1352_));
  NA2        o1324(.A(ori_ori_n1352_), .B(ori_ori_n1351_), .Y(ori_ori_n1353_));
  INV        o1325(.A(ori_ori_n1353_), .Y(ori_ori_n1354_));
  NO3        o1326(.A(ori_ori_n1354_), .B(ori_ori_n1350_), .C(ori_ori_n1349_), .Y(ori_ori_n1355_));
  NA2        o1327(.A(ori_ori_n1065_), .B(ori_ori_n477_), .Y(ori_ori_n1356_));
  NO4        o1328(.A(ori_ori_n1356_), .B(ori_ori_n1053_), .C(ori_ori_n453_), .D(ori_ori_n45_), .Y(ori_ori_n1357_));
  NO3        o1329(.A(ori_ori_n41_), .B(i), .C(h), .Y(ori_ori_n1358_));
  NO2        o1330(.A(ori_ori_n1054_), .B(ori_ori_n1357_), .Y(ori_ori_n1359_));
  AN3        o1331(.A(ori_ori_n1359_), .B(ori_ori_n1355_), .C(ori_ori_n1346_), .Y(ori_ori_n1360_));
  NA2        o1332(.A(ori_ori_n1312_), .B(ori_ori_n392_), .Y(ori_ori_n1361_));
  INV        o1333(.A(ori_ori_n1361_), .Y(ori_ori_n1362_));
  NA2        o1334(.A(ori_ori_n1341_), .B(ori_ori_n218_), .Y(ori_ori_n1363_));
  NA2        o1335(.A(ori_ori_n1073_), .B(ori_ori_n1356_), .Y(ori_ori_n1364_));
  NAi31      o1336(.An(ori_ori_n1362_), .B(ori_ori_n1364_), .C(ori_ori_n1363_), .Y(ori_ori_n1365_));
  NO4        o1337(.A(ori_ori_n131_), .B(o), .C(f), .D(e), .Y(ori_ori_n1366_));
  NA2        o1338(.A(ori_ori_n196_), .B(ori_ori_n99_), .Y(ori_ori_n1367_));
  NA2        o1339(.A(ori_ori_n1314_), .B(ori_ori_n1339_), .Y(ori_ori_n1368_));
  INV        o1340(.A(ori_ori_n1368_), .Y(ori_ori_n1369_));
  OR3        o1341(.A(ori_ori_n550_), .B(ori_ori_n549_), .C(ori_ori_n112_), .Y(ori_ori_n1370_));
  NA2        o1342(.A(ori_ori_n1090_), .B(ori_ori_n421_), .Y(ori_ori_n1371_));
  NO2        o1343(.A(ori_ori_n1371_), .B(ori_ori_n449_), .Y(ori_ori_n1372_));
  AO210      o1344(.A0(ori_ori_n1372_), .A1(ori_ori_n115_), .B0(ori_ori_n1369_), .Y(ori_ori_n1373_));
  NO2        o1345(.A(ori_ori_n1373_), .B(ori_ori_n1365_), .Y(ori_ori_n1374_));
  NA4        o1346(.A(ori_ori_n1374_), .B(ori_ori_n1360_), .C(ori_ori_n1342_), .D(ori_ori_n1326_), .Y(ori_ori_n1375_));
  NO2        o1347(.A(ori_ori_n1101_), .B(ori_ori_n110_), .Y(ori_ori_n1376_));
  NA2        o1348(.A(ori_ori_n392_), .B(ori_ori_n56_), .Y(ori_ori_n1377_));
  AOI210     o1349(.A0(ori_ori_n1377_), .A1(ori_ori_n1048_), .B0(ori_ori_n1338_), .Y(ori_ori_n1378_));
  NA2        o1350(.A(ori_ori_n218_), .B(ori_ori_n181_), .Y(ori_ori_n1379_));
  AOI210     o1351(.A0(ori_ori_n1379_), .A1(ori_ori_n1157_), .B0(ori_ori_n1377_), .Y(ori_ori_n1380_));
  NO2        o1352(.A(ori_ori_n1066_), .B(ori_ori_n1063_), .Y(ori_ori_n1381_));
  NO3        o1353(.A(ori_ori_n1381_), .B(ori_ori_n1380_), .C(ori_ori_n1378_), .Y(ori_ori_n1382_));
  NO2        o1354(.A(ori_ori_n404_), .B(j), .Y(ori_ori_n1383_));
  NA2        o1355(.A(ori_ori_n1358_), .B(ori_ori_n1090_), .Y(ori_ori_n1384_));
  NAi41      o1356(.An(ori_ori_n1347_), .B(ori_ori_n1060_), .C(ori_ori_n170_), .D(ori_ori_n151_), .Y(ori_ori_n1385_));
  NA2        o1357(.A(ori_ori_n1385_), .B(ori_ori_n1384_), .Y(ori_ori_n1386_));
  NA3        o1358(.A(o), .B(ori_ori_n1383_), .C(ori_ori_n160_), .Y(ori_ori_n1387_));
  INV        o1359(.A(ori_ori_n1387_), .Y(ori_ori_n1388_));
  NO3        o1360(.A(ori_ori_n754_), .B(ori_ori_n176_), .C(ori_ori_n424_), .Y(ori_ori_n1389_));
  NO3        o1361(.A(ori_ori_n1389_), .B(ori_ori_n1388_), .C(ori_ori_n1386_), .Y(ori_ori_n1390_));
  NO3        o1362(.A(ori_ori_n1063_), .B(ori_ori_n591_), .C(o), .Y(ori_ori_n1391_));
  NOi21      o1363(.An(ori_ori_n1379_), .B(ori_ori_n1391_), .Y(ori_ori_n1392_));
  AOI210     o1364(.A0(ori_ori_n1392_), .A1(ori_ori_n1367_), .B0(ori_ori_n1048_), .Y(ori_ori_n1393_));
  OR2        o1365(.A(n), .B(i), .Y(ori_ori_n1394_));
  NA2        o1366(.A(ori_ori_n1394_), .B(ori_ori_n49_), .Y(ori_ori_n1395_));
  AOI220     o1367(.A0(ori_ori_n1395_), .A1(ori_ori_n1145_), .B0(ori_ori_n834_), .B1(ori_ori_n196_), .Y(ori_ori_n1396_));
  INV        o1368(.A(ori_ori_n1396_), .Y(ori_ori_n1397_));
  NO2        o1369(.A(ori_ori_n679_), .B(ori_ori_n178_), .Y(ori_ori_n1398_));
  NO3        o1370(.A(ori_ori_n1398_), .B(ori_ori_n1397_), .C(ori_ori_n1393_), .Y(ori_ori_n1399_));
  NO3        o1371(.A(ori_ori_n1076_), .B(ori_ori_n1309_), .C(ori_ori_n49_), .Y(ori_ori_n1400_));
  NO2        o1372(.A(ori_ori_n1063_), .B(h), .Y(ori_ori_n1401_));
  NA2        o1373(.A(ori_ori_n1401_), .B(ori_ori_n1043_), .Y(ori_ori_n1402_));
  NO2        o1374(.A(ori_ori_n1402_), .B(c), .Y(ori_ori_n1403_));
  NA3        o1375(.A(ori_ori_n1376_), .B(ori_ori_n477_), .C(f), .Y(ori_ori_n1404_));
  NA2        o1376(.A(ori_ori_n181_), .B(ori_ori_n112_), .Y(ori_ori_n1405_));
  NO2        o1377(.A(ori_ori_n1476_), .B(ori_ori_n1404_), .Y(ori_ori_n1406_));
  NO2        o1378(.A(ori_ori_n1299_), .B(ori_ori_n176_), .Y(ori_ori_n1407_));
  NOi21      o1379(.An(d), .B(f), .Y(ori_ori_n1408_));
  NO3        o1380(.A(ori_ori_n1352_), .B(ori_ori_n1408_), .C(ori_ori_n40_), .Y(ori_ori_n1409_));
  NA2        o1381(.A(ori_ori_n1409_), .B(ori_ori_n1407_), .Y(ori_ori_n1410_));
  INV        o1382(.A(ori_ori_n1410_), .Y(ori_ori_n1411_));
  NO3        o1383(.A(ori_ori_n1411_), .B(ori_ori_n1406_), .C(ori_ori_n1403_), .Y(ori_ori_n1412_));
  NA4        o1384(.A(ori_ori_n1412_), .B(ori_ori_n1399_), .C(ori_ori_n1390_), .D(ori_ori_n1382_), .Y(ori_ori_n1413_));
  NO2        o1385(.A(ori_ori_n1065_), .B(ori_ori_n40_), .Y(ori_ori_n1414_));
  NO2        o1386(.A(ori_ori_n477_), .B(ori_ori_n304_), .Y(ori_ori_n1415_));
  OAI210     o1387(.A0(ori_ori_n1415_), .A1(ori_ori_n1414_), .B0(ori_ori_n1322_), .Y(ori_ori_n1416_));
  OAI210     o1388(.A0(ori_ori_n1366_), .A1(ori_ori_n1312_), .B0(ori_ori_n893_), .Y(ori_ori_n1417_));
  NO2        o1389(.A(ori_ori_n1041_), .B(ori_ori_n131_), .Y(ori_ori_n1418_));
  NA2        o1390(.A(ori_ori_n1418_), .B(ori_ori_n630_), .Y(ori_ori_n1419_));
  NA3        o1391(.A(ori_ori_n1419_), .B(ori_ori_n1417_), .C(ori_ori_n1416_), .Y(ori_ori_n1420_));
  NA2        o1392(.A(ori_ori_n1344_), .B(ori_ori_n1408_), .Y(ori_ori_n1421_));
  NO2        o1393(.A(ori_ori_n1421_), .B(m), .Y(ori_ori_n1422_));
  NA3        o1394(.A(ori_ori_n1074_), .B(ori_ori_n109_), .C(ori_ori_n224_), .Y(ori_ori_n1423_));
  NO2        o1395(.A(ori_ori_n152_), .B(ori_ori_n183_), .Y(ori_ori_n1424_));
  OAI210     o1396(.A0(ori_ori_n1424_), .A1(ori_ori_n110_), .B0(ori_ori_n1351_), .Y(ori_ori_n1425_));
  NA2        o1397(.A(ori_ori_n1425_), .B(ori_ori_n1423_), .Y(ori_ori_n1426_));
  NO3        o1398(.A(ori_ori_n1426_), .B(ori_ori_n1422_), .C(ori_ori_n1420_), .Y(ori_ori_n1427_));
  NO2        o1399(.A(ori_ori_n1308_), .B(e), .Y(ori_ori_n1428_));
  NA2        o1400(.A(ori_ori_n1428_), .B(ori_ori_n419_), .Y(ori_ori_n1429_));
  BUFFER     o1401(.A(ori_ori_n131_), .Y(ori_ori_n1430_));
  NO2        o1402(.A(ori_ori_n1430_), .B(ori_ori_n1429_), .Y(ori_ori_n1431_));
  NO2        o1403(.A(ori_ori_n1370_), .B(ori_ori_n363_), .Y(ori_ori_n1432_));
  NO2        o1404(.A(ori_ori_n1432_), .B(ori_ori_n1431_), .Y(ori_ori_n1433_));
  NO2        o1405(.A(ori_ori_n183_), .B(c), .Y(ori_ori_n1434_));
  OAI210     o1406(.A0(ori_ori_n1434_), .A1(ori_ori_n1428_), .B0(ori_ori_n181_), .Y(ori_ori_n1435_));
  AOI210     o1407(.A0(ori_ori_n542_), .A1(ori_ori_n379_), .B0(ori_ori_n1435_), .Y(ori_ori_n1436_));
  AOI210     o1408(.A0(j), .A1(ori_ori_n1341_), .B0(ori_ori_n1400_), .Y(ori_ori_n1437_));
  INV        o1409(.A(ori_ori_n1098_), .Y(ori_ori_n1438_));
  OAI210     o1410(.A0(ori_ori_n1438_), .A1(ori_ori_n69_), .B0(ori_ori_n1437_), .Y(ori_ori_n1439_));
  AOI210     o1411(.A0(ori_ori_n909_), .A1(ori_ori_n431_), .B0(ori_ori_n105_), .Y(ori_ori_n1440_));
  OR2        o1412(.A(ori_ori_n1440_), .B(ori_ori_n549_), .Y(ori_ori_n1441_));
  NO2        o1413(.A(ori_ori_n1441_), .B(ori_ori_n176_), .Y(ori_ori_n1442_));
  NA3        o1414(.A(ori_ori_n1074_), .B(ori_ori_n1071_), .C(ori_ori_n224_), .Y(ori_ori_n1443_));
  NO2        o1415(.A(ori_ori_n49_), .B(l), .Y(ori_ori_n1444_));
  INV        o1416(.A(ori_ori_n494_), .Y(ori_ori_n1445_));
  NA2        o1417(.A(ori_ori_n1445_), .B(ori_ori_n1444_), .Y(ori_ori_n1446_));
  NO2        o1418(.A(m), .B(i), .Y(ori_ori_n1447_));
  BUFFER     o1419(.A(ori_ori_n1447_), .Y(ori_ori_n1448_));
  NA2        o1420(.A(ori_ori_n1448_), .B(ori_ori_n1343_), .Y(ori_ori_n1449_));
  NA3        o1421(.A(ori_ori_n1449_), .B(ori_ori_n1446_), .C(ori_ori_n1443_), .Y(ori_ori_n1450_));
  NO4        o1422(.A(ori_ori_n1450_), .B(ori_ori_n1442_), .C(ori_ori_n1439_), .D(ori_ori_n1436_), .Y(ori_ori_n1451_));
  NA3        o1423(.A(ori_ori_n1451_), .B(ori_ori_n1433_), .C(ori_ori_n1427_), .Y(ori_ori_n1452_));
  NA3        o1424(.A(ori_ori_n968_), .B(ori_ori_n138_), .C(ori_ori_n46_), .Y(ori_ori_n1453_));
  INV        o1425(.A(ori_ori_n1453_), .Y(ori_ori_n1454_));
  INV        o1426(.A(d), .Y(ori_ori_n1455_));
  NA2        o1427(.A(ori_ori_n1455_), .B(ori_ori_n1401_), .Y(ori_ori_n1456_));
  NO2        o1428(.A(ori_ori_n71_), .B(c), .Y(ori_ori_n1457_));
  NA2        o1429(.A(ori_ori_n1407_), .B(ori_ori_n1457_), .Y(ori_ori_n1458_));
  NA2        o1430(.A(ori_ori_n1458_), .B(ori_ori_n1456_), .Y(ori_ori_n1459_));
  NO2        o1431(.A(ori_ori_n1459_), .B(ori_ori_n1454_), .Y(ori_ori_n1460_));
  AOI210     o1432(.A0(ori_ori_n158_), .A1(ori_ori_n56_), .B0(ori_ori_n1428_), .Y(ori_ori_n1461_));
  NO2        o1433(.A(ori_ori_n1461_), .B(ori_ori_n1405_), .Y(ori_ori_n1462_));
  INV        o1434(.A(ori_ori_n1462_), .Y(ori_ori_n1463_));
  NOi31      o1435(.An(ori_ori_n30_), .B(ori_ori_n1479_), .C(n), .Y(ori_ori_n1464_));
  INV        o1436(.A(ori_ori_n1464_), .Y(ori_ori_n1465_));
  NO2        o1437(.A(ori_ori_n1371_), .B(d), .Y(ori_ori_n1466_));
  NA4        o1438(.A(ori_ori_n1477_), .B(ori_ori_n1465_), .C(ori_ori_n1463_), .D(ori_ori_n1460_), .Y(ori_ori_n1467_));
  OR4        o1439(.A(ori_ori_n1467_), .B(ori_ori_n1452_), .C(ori_ori_n1413_), .D(ori_ori_n1375_), .Y(ori04));
  NO3        o1440(.A(ori_ori_n1319_), .B(ori_ori_n91_), .C(k), .Y(ori_ori_n1469_));
  AOI210     o1441(.A0(ori_ori_n1469_), .A1(ori_ori_n1049_), .B0(ori_ori_n1159_), .Y(ori_ori_n1470_));
  INV        o1442(.A(ori_ori_n1470_), .Y(ori_ori_n1471_));
  NO3        o1443(.A(ori_ori_n1471_), .B(ori_ori_n1058_), .C(ori_ori_n1047_), .Y(ori_ori_n1472_));
  NA3        o1444(.A(ori_ori_n1472_), .B(ori_ori_n1088_), .C(ori_ori_n1078_), .Y(ori05));
  INV        o1445(.A(ori_ori_n113_), .Y(ori_ori_n1476_));
  INV        o1446(.A(ori_ori_n1466_), .Y(ori_ori_n1477_));
  INV        o1447(.A(h), .Y(ori_ori_n1478_));
  INV        o1448(.A(ori_ori_n161_), .Y(ori_ori_n1479_));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(m), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(m), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(m), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(m), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(m), .Y(mai_mai_n51_));
  INV        m0023(.A(mai_mai_n51_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO3        m0025(.A(mai_mai_n53_), .B(mai_mai_n48_), .C(mai_mai_n39_), .Y(mai_mai_n54_));
  AOI210     m0026(.A0(mai_mai_n54_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NAi21      m0031(.An(i), .B(h), .Y(mai_mai_n60_));
  NAi31      m0032(.An(i), .B(l), .C(j), .Y(mai_mai_n61_));
  NAi41      m0033(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n62_));
  NA2        m0034(.A(m), .B(f), .Y(mai_mai_n63_));
  NO2        m0035(.A(mai_mai_n63_), .B(mai_mai_n62_), .Y(mai_mai_n64_));
  NAi21      m0036(.An(i), .B(j), .Y(mai_mai_n65_));
  NAi32      m0037(.An(n), .Bn(k), .C(m), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi31      m0039(.An(l), .B(m), .C(k), .Y(mai_mai_n68_));
  NAi21      m0040(.An(e), .B(h), .Y(mai_mai_n69_));
  NAi41      m0041(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n70_));
  NA2        m0042(.A(mai_mai_n67_), .B(mai_mai_n64_), .Y(mai_mai_n71_));
  INV        m0043(.A(m), .Y(mai_mai_n72_));
  NOi21      m0044(.An(k), .B(l), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  AN4        m0046(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n75_));
  NOi31      m0047(.An(h), .B(m), .C(f), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n77_));
  NAi32      m0049(.An(m), .Bn(k), .C(j), .Y(mai_mai_n78_));
  NOi32      m0050(.An(h), .Bn(m), .C(f), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n79_), .B(mai_mai_n75_), .Y(mai_mai_n80_));
  OA220      m0052(.A0(mai_mai_n80_), .A1(mai_mai_n78_), .B0(mai_mai_n77_), .B1(mai_mai_n74_), .Y(mai_mai_n81_));
  NA2        m0053(.A(mai_mai_n81_), .B(mai_mai_n71_), .Y(mai_mai_n82_));
  INV        m0054(.A(n), .Y(mai_mai_n83_));
  NOi32      m0055(.An(e), .Bn(b), .C(d), .Y(mai_mai_n84_));
  NA2        m0056(.A(mai_mai_n84_), .B(mai_mai_n83_), .Y(mai_mai_n85_));
  INV        m0057(.A(j), .Y(mai_mai_n86_));
  AN3        m0058(.A(m), .B(k), .C(i), .Y(mai_mai_n87_));
  NA3        m0059(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(m), .Y(mai_mai_n88_));
  NO2        m0060(.A(mai_mai_n88_), .B(f), .Y(mai_mai_n89_));
  NAi32      m0061(.An(m), .Bn(f), .C(h), .Y(mai_mai_n90_));
  NAi31      m0062(.An(j), .B(m), .C(l), .Y(mai_mai_n91_));
  NO2        m0063(.A(mai_mai_n91_), .B(mai_mai_n90_), .Y(mai_mai_n92_));
  NA2        m0064(.A(m), .B(l), .Y(mai_mai_n93_));
  NAi31      m0065(.An(k), .B(j), .C(m), .Y(mai_mai_n94_));
  NO3        m0066(.A(mai_mai_n94_), .B(mai_mai_n93_), .C(f), .Y(mai_mai_n95_));
  AN2        m0067(.A(j), .B(m), .Y(mai_mai_n96_));
  NOi32      m0068(.An(m), .Bn(l), .C(i), .Y(mai_mai_n97_));
  NOi21      m0069(.An(m), .B(i), .Y(mai_mai_n98_));
  NOi32      m0070(.An(m), .Bn(j), .C(k), .Y(mai_mai_n99_));
  AOI220     m0071(.A0(mai_mai_n99_), .A1(mai_mai_n98_), .B0(mai_mai_n97_), .B1(mai_mai_n96_), .Y(mai_mai_n100_));
  NO2        m0072(.A(mai_mai_n100_), .B(f), .Y(mai_mai_n101_));
  NO4        m0073(.A(mai_mai_n101_), .B(mai_mai_n95_), .C(mai_mai_n92_), .D(mai_mai_n89_), .Y(mai_mai_n102_));
  NAi41      m0074(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n103_));
  AN2        m0075(.A(e), .B(b), .Y(mai_mai_n104_));
  NOi31      m0076(.An(c), .B(h), .C(f), .Y(mai_mai_n105_));
  NA2        m0077(.A(mai_mai_n105_), .B(mai_mai_n104_), .Y(mai_mai_n106_));
  NO2        m0078(.A(mai_mai_n106_), .B(mai_mai_n103_), .Y(mai_mai_n107_));
  NOi21      m0079(.An(m), .B(f), .Y(mai_mai_n108_));
  NOi21      m0080(.An(i), .B(h), .Y(mai_mai_n109_));
  NA3        m0081(.A(mai_mai_n109_), .B(mai_mai_n108_), .C(mai_mai_n36_), .Y(mai_mai_n110_));
  INV        m0082(.A(a), .Y(mai_mai_n111_));
  NA2        m0083(.A(mai_mai_n104_), .B(mai_mai_n111_), .Y(mai_mai_n112_));
  INV        m0084(.A(l), .Y(mai_mai_n113_));
  NOi21      m0085(.An(m), .B(n), .Y(mai_mai_n114_));
  AN2        m0086(.A(k), .B(h), .Y(mai_mai_n115_));
  NO2        m0087(.A(mai_mai_n110_), .B(mai_mai_n85_), .Y(mai_mai_n116_));
  INV        m0088(.A(b), .Y(mai_mai_n117_));
  NA2        m0089(.A(l), .B(j), .Y(mai_mai_n118_));
  AN2        m0090(.A(k), .B(i), .Y(mai_mai_n119_));
  NA2        m0091(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n120_));
  NA2        m0092(.A(m), .B(e), .Y(mai_mai_n121_));
  NOi32      m0093(.An(c), .Bn(a), .C(d), .Y(mai_mai_n122_));
  NA2        m0094(.A(mai_mai_n122_), .B(mai_mai_n114_), .Y(mai_mai_n123_));
  NO4        m0095(.A(mai_mai_n123_), .B(mai_mai_n121_), .C(mai_mai_n120_), .D(mai_mai_n117_), .Y(mai_mai_n124_));
  NO3        m0096(.A(mai_mai_n124_), .B(mai_mai_n116_), .C(mai_mai_n107_), .Y(mai_mai_n125_));
  OAI210     m0097(.A0(mai_mai_n102_), .A1(mai_mai_n85_), .B0(mai_mai_n125_), .Y(mai_mai_n126_));
  NOi31      m0098(.An(k), .B(m), .C(j), .Y(mai_mai_n127_));
  NOi31      m0099(.An(k), .B(m), .C(i), .Y(mai_mai_n128_));
  NOi32      m0100(.An(f), .Bn(b), .C(e), .Y(mai_mai_n129_));
  NAi21      m0101(.An(m), .B(h), .Y(mai_mai_n130_));
  NAi21      m0102(.An(m), .B(n), .Y(mai_mai_n131_));
  NAi21      m0103(.An(j), .B(k), .Y(mai_mai_n132_));
  NO3        m0104(.A(mai_mai_n132_), .B(mai_mai_n131_), .C(mai_mai_n130_), .Y(mai_mai_n133_));
  NAi41      m0105(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n134_));
  NAi31      m0106(.An(j), .B(k), .C(h), .Y(mai_mai_n135_));
  NA2        m0107(.A(mai_mai_n133_), .B(mai_mai_n129_), .Y(mai_mai_n136_));
  NO2        m0108(.A(k), .B(j), .Y(mai_mai_n137_));
  NO2        m0109(.A(mai_mai_n137_), .B(mai_mai_n131_), .Y(mai_mai_n138_));
  AN2        m0110(.A(k), .B(j), .Y(mai_mai_n139_));
  NAi21      m0111(.An(c), .B(b), .Y(mai_mai_n140_));
  NA2        m0112(.A(f), .B(d), .Y(mai_mai_n141_));
  NO4        m0113(.A(mai_mai_n141_), .B(mai_mai_n140_), .C(mai_mai_n139_), .D(mai_mai_n130_), .Y(mai_mai_n142_));
  NA2        m0114(.A(h), .B(c), .Y(mai_mai_n143_));
  NAi31      m0115(.An(f), .B(e), .C(b), .Y(mai_mai_n144_));
  NA2        m0116(.A(mai_mai_n142_), .B(mai_mai_n138_), .Y(mai_mai_n145_));
  NA2        m0117(.A(d), .B(b), .Y(mai_mai_n146_));
  NAi21      m0118(.An(e), .B(f), .Y(mai_mai_n147_));
  NO2        m0119(.A(mai_mai_n147_), .B(mai_mai_n146_), .Y(mai_mai_n148_));
  NA2        m0120(.A(b), .B(a), .Y(mai_mai_n149_));
  NAi21      m0121(.An(e), .B(m), .Y(mai_mai_n150_));
  NAi21      m0122(.An(c), .B(d), .Y(mai_mai_n151_));
  NAi31      m0123(.An(l), .B(k), .C(h), .Y(mai_mai_n152_));
  NO2        m0124(.A(mai_mai_n131_), .B(mai_mai_n152_), .Y(mai_mai_n153_));
  NA2        m0125(.A(mai_mai_n145_), .B(mai_mai_n136_), .Y(mai_mai_n154_));
  NAi31      m0126(.An(e), .B(f), .C(b), .Y(mai_mai_n155_));
  NOi21      m0127(.An(m), .B(d), .Y(mai_mai_n156_));
  NO2        m0128(.A(mai_mai_n156_), .B(mai_mai_n155_), .Y(mai_mai_n157_));
  NOi21      m0129(.An(h), .B(i), .Y(mai_mai_n158_));
  NOi21      m0130(.An(k), .B(m), .Y(mai_mai_n159_));
  NA3        m0131(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(n), .Y(mai_mai_n160_));
  NOi21      m0132(.An(mai_mai_n157_), .B(mai_mai_n160_), .Y(mai_mai_n161_));
  NOi21      m0133(.An(h), .B(m), .Y(mai_mai_n162_));
  NO2        m0134(.A(mai_mai_n141_), .B(mai_mai_n140_), .Y(mai_mai_n163_));
  NA2        m0135(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  NAi31      m0136(.An(l), .B(j), .C(h), .Y(mai_mai_n165_));
  NO2        m0137(.A(mai_mai_n165_), .B(mai_mai_n49_), .Y(mai_mai_n166_));
  NA2        m0138(.A(mai_mai_n166_), .B(mai_mai_n64_), .Y(mai_mai_n167_));
  NOi32      m0139(.An(n), .Bn(k), .C(m), .Y(mai_mai_n168_));
  NA2        m0140(.A(l), .B(i), .Y(mai_mai_n169_));
  NA2        m0141(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  OAI210     m0142(.A0(mai_mai_n170_), .A1(mai_mai_n164_), .B0(mai_mai_n167_), .Y(mai_mai_n171_));
  NAi31      m0143(.An(d), .B(f), .C(c), .Y(mai_mai_n172_));
  NAi31      m0144(.An(e), .B(f), .C(c), .Y(mai_mai_n173_));
  NA2        m0145(.A(mai_mai_n173_), .B(mai_mai_n172_), .Y(mai_mai_n174_));
  NA2        m0146(.A(j), .B(h), .Y(mai_mai_n175_));
  OR3        m0147(.A(n), .B(m), .C(k), .Y(mai_mai_n176_));
  NO2        m0148(.A(mai_mai_n176_), .B(mai_mai_n175_), .Y(mai_mai_n177_));
  NAi32      m0149(.An(m), .Bn(k), .C(n), .Y(mai_mai_n178_));
  NO2        m0150(.A(mai_mai_n178_), .B(mai_mai_n175_), .Y(mai_mai_n179_));
  AOI220     m0151(.A0(mai_mai_n179_), .A1(mai_mai_n157_), .B0(mai_mai_n177_), .B1(mai_mai_n174_), .Y(mai_mai_n180_));
  NO2        m0152(.A(n), .B(m), .Y(mai_mai_n181_));
  NA2        m0153(.A(mai_mai_n181_), .B(mai_mai_n50_), .Y(mai_mai_n182_));
  NAi21      m0154(.An(f), .B(e), .Y(mai_mai_n183_));
  NA2        m0155(.A(d), .B(c), .Y(mai_mai_n184_));
  NO2        m0156(.A(mai_mai_n184_), .B(mai_mai_n183_), .Y(mai_mai_n185_));
  NOi21      m0157(.An(mai_mai_n185_), .B(mai_mai_n182_), .Y(mai_mai_n186_));
  NAi21      m0158(.An(d), .B(c), .Y(mai_mai_n187_));
  NAi31      m0159(.An(m), .B(n), .C(b), .Y(mai_mai_n188_));
  NA2        m0160(.A(k), .B(i), .Y(mai_mai_n189_));
  NAi21      m0161(.An(h), .B(f), .Y(mai_mai_n190_));
  NO2        m0162(.A(mai_mai_n190_), .B(mai_mai_n189_), .Y(mai_mai_n191_));
  NO2        m0163(.A(mai_mai_n188_), .B(mai_mai_n151_), .Y(mai_mai_n192_));
  NA2        m0164(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n193_));
  NOi32      m0165(.An(f), .Bn(c), .C(d), .Y(mai_mai_n194_));
  NOi32      m0166(.An(f), .Bn(c), .C(e), .Y(mai_mai_n195_));
  NO2        m0167(.A(mai_mai_n195_), .B(mai_mai_n194_), .Y(mai_mai_n196_));
  NO3        m0168(.A(n), .B(m), .C(j), .Y(mai_mai_n197_));
  NA2        m0169(.A(mai_mai_n197_), .B(mai_mai_n115_), .Y(mai_mai_n198_));
  AO210      m0170(.A0(mai_mai_n198_), .A1(mai_mai_n182_), .B0(mai_mai_n196_), .Y(mai_mai_n199_));
  NAi41      m0171(.An(mai_mai_n186_), .B(mai_mai_n199_), .C(mai_mai_n193_), .D(mai_mai_n180_), .Y(mai_mai_n200_));
  OR4        m0172(.A(mai_mai_n200_), .B(mai_mai_n171_), .C(mai_mai_n161_), .D(mai_mai_n154_), .Y(mai_mai_n201_));
  NO4        m0173(.A(mai_mai_n201_), .B(mai_mai_n126_), .C(mai_mai_n82_), .D(mai_mai_n55_), .Y(mai_mai_n202_));
  NA3        m0174(.A(m), .B(mai_mai_n113_), .C(j), .Y(mai_mai_n203_));
  NAi31      m0175(.An(n), .B(h), .C(m), .Y(mai_mai_n204_));
  NO2        m0176(.A(mai_mai_n204_), .B(mai_mai_n203_), .Y(mai_mai_n205_));
  NOi32      m0177(.An(m), .Bn(k), .C(l), .Y(mai_mai_n206_));
  NA3        m0178(.A(mai_mai_n206_), .B(mai_mai_n86_), .C(m), .Y(mai_mai_n207_));
  NO2        m0179(.A(mai_mai_n207_), .B(n), .Y(mai_mai_n208_));
  NOi21      m0180(.An(k), .B(j), .Y(mai_mai_n209_));
  AN2        m0181(.A(i), .B(m), .Y(mai_mai_n210_));
  NA3        m0182(.A(mai_mai_n73_), .B(mai_mai_n210_), .C(mai_mai_n114_), .Y(mai_mai_n211_));
  INV        m0183(.A(mai_mai_n211_), .Y(mai_mai_n212_));
  NO2        m0184(.A(mai_mai_n208_), .B(mai_mai_n205_), .Y(mai_mai_n213_));
  NAi41      m0185(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n214_));
  INV        m0186(.A(mai_mai_n214_), .Y(mai_mai_n215_));
  INV        m0187(.A(f), .Y(mai_mai_n216_));
  INV        m0188(.A(m), .Y(mai_mai_n217_));
  NOi31      m0189(.An(i), .B(j), .C(h), .Y(mai_mai_n218_));
  NOi21      m0190(.An(l), .B(m), .Y(mai_mai_n219_));
  NA2        m0191(.A(mai_mai_n219_), .B(mai_mai_n218_), .Y(mai_mai_n220_));
  NO3        m0192(.A(mai_mai_n220_), .B(mai_mai_n217_), .C(mai_mai_n216_), .Y(mai_mai_n221_));
  NA2        m0193(.A(mai_mai_n221_), .B(mai_mai_n215_), .Y(mai_mai_n222_));
  OAI210     m0194(.A0(mai_mai_n213_), .A1(mai_mai_n32_), .B0(mai_mai_n222_), .Y(mai_mai_n223_));
  NOi21      m0195(.An(n), .B(m), .Y(mai_mai_n224_));
  NOi32      m0196(.An(l), .Bn(i), .C(j), .Y(mai_mai_n225_));
  NA2        m0197(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n226_));
  OA220      m0198(.A0(mai_mai_n226_), .A1(mai_mai_n106_), .B0(mai_mai_n78_), .B1(mai_mai_n77_), .Y(mai_mai_n227_));
  NAi21      m0199(.An(j), .B(h), .Y(mai_mai_n228_));
  XN2        m0200(.A(i), .B(h), .Y(mai_mai_n229_));
  NA2        m0201(.A(mai_mai_n229_), .B(mai_mai_n228_), .Y(mai_mai_n230_));
  NOi31      m0202(.An(k), .B(n), .C(m), .Y(mai_mai_n231_));
  NOi31      m0203(.An(mai_mai_n231_), .B(mai_mai_n184_), .C(mai_mai_n183_), .Y(mai_mai_n232_));
  NA2        m0204(.A(mai_mai_n232_), .B(mai_mai_n230_), .Y(mai_mai_n233_));
  NAi31      m0205(.An(f), .B(e), .C(c), .Y(mai_mai_n234_));
  NO4        m0206(.A(mai_mai_n234_), .B(mai_mai_n176_), .C(mai_mai_n175_), .D(mai_mai_n59_), .Y(mai_mai_n235_));
  NA4        m0207(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n236_));
  NAi32      m0208(.An(m), .Bn(i), .C(k), .Y(mai_mai_n237_));
  NO3        m0209(.A(mai_mai_n237_), .B(mai_mai_n90_), .C(mai_mai_n236_), .Y(mai_mai_n238_));
  INV        m0210(.A(k), .Y(mai_mai_n239_));
  NO2        m0211(.A(mai_mai_n238_), .B(mai_mai_n235_), .Y(mai_mai_n240_));
  NAi21      m0212(.An(n), .B(a), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n241_), .B(mai_mai_n146_), .Y(mai_mai_n242_));
  NAi41      m0214(.An(m), .B(m), .C(k), .D(h), .Y(mai_mai_n243_));
  NO2        m0215(.A(mai_mai_n243_), .B(e), .Y(mai_mai_n244_));
  NO3        m0216(.A(mai_mai_n147_), .B(mai_mai_n94_), .C(mai_mai_n93_), .Y(mai_mai_n245_));
  OAI210     m0217(.A0(mai_mai_n245_), .A1(mai_mai_n244_), .B0(mai_mai_n242_), .Y(mai_mai_n246_));
  AN4        m0218(.A(mai_mai_n246_), .B(mai_mai_n240_), .C(mai_mai_n233_), .D(mai_mai_n227_), .Y(mai_mai_n247_));
  OR2        m0219(.A(h), .B(m), .Y(mai_mai_n248_));
  NO2        m0220(.A(mai_mai_n248_), .B(mai_mai_n103_), .Y(mai_mai_n249_));
  NA2        m0221(.A(mai_mai_n249_), .B(mai_mai_n129_), .Y(mai_mai_n250_));
  NAi41      m0222(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n251_));
  NO2        m0223(.A(mai_mai_n251_), .B(mai_mai_n216_), .Y(mai_mai_n252_));
  NA2        m0224(.A(mai_mai_n159_), .B(mai_mai_n109_), .Y(mai_mai_n253_));
  NAi21      m0225(.An(mai_mai_n253_), .B(mai_mai_n252_), .Y(mai_mai_n254_));
  NO2        m0226(.A(n), .B(a), .Y(mai_mai_n255_));
  NAi31      m0227(.An(mai_mai_n243_), .B(mai_mai_n255_), .C(mai_mai_n104_), .Y(mai_mai_n256_));
  AN2        m0228(.A(mai_mai_n256_), .B(mai_mai_n254_), .Y(mai_mai_n257_));
  NAi21      m0229(.An(h), .B(i), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n181_), .B(k), .Y(mai_mai_n259_));
  NO2        m0231(.A(mai_mai_n259_), .B(mai_mai_n258_), .Y(mai_mai_n260_));
  NA2        m0232(.A(mai_mai_n260_), .B(mai_mai_n194_), .Y(mai_mai_n261_));
  NA3        m0233(.A(mai_mai_n261_), .B(mai_mai_n257_), .C(mai_mai_n250_), .Y(mai_mai_n262_));
  NOi21      m0234(.An(m), .B(e), .Y(mai_mai_n263_));
  NO2        m0235(.A(mai_mai_n70_), .B(mai_mai_n72_), .Y(mai_mai_n264_));
  NA2        m0236(.A(mai_mai_n264_), .B(mai_mai_n263_), .Y(mai_mai_n265_));
  NOi32      m0237(.An(l), .Bn(j), .C(i), .Y(mai_mai_n266_));
  AOI210     m0238(.A0(mai_mai_n73_), .A1(mai_mai_n86_), .B0(mai_mai_n266_), .Y(mai_mai_n267_));
  NO2        m0239(.A(mai_mai_n258_), .B(mai_mai_n44_), .Y(mai_mai_n268_));
  NAi21      m0240(.An(f), .B(m), .Y(mai_mai_n269_));
  NO2        m0241(.A(mai_mai_n269_), .B(mai_mai_n62_), .Y(mai_mai_n270_));
  NO2        m0242(.A(mai_mai_n66_), .B(mai_mai_n118_), .Y(mai_mai_n271_));
  AOI220     m0243(.A0(mai_mai_n271_), .A1(mai_mai_n270_), .B0(mai_mai_n268_), .B1(mai_mai_n64_), .Y(mai_mai_n272_));
  OAI210     m0244(.A0(mai_mai_n267_), .A1(mai_mai_n265_), .B0(mai_mai_n272_), .Y(mai_mai_n273_));
  NOi41      m0245(.An(mai_mai_n247_), .B(mai_mai_n273_), .C(mai_mai_n262_), .D(mai_mai_n223_), .Y(mai_mai_n274_));
  NO4        m0246(.A(mai_mai_n205_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n275_));
  NO2        m0247(.A(mai_mai_n275_), .B(mai_mai_n112_), .Y(mai_mai_n276_));
  NA3        m0248(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n277_));
  NAi21      m0249(.An(h), .B(m), .Y(mai_mai_n278_));
  NO2        m0250(.A(mai_mai_n253_), .B(mai_mai_n269_), .Y(mai_mai_n279_));
  NAi31      m0251(.An(m), .B(k), .C(h), .Y(mai_mai_n280_));
  NO3        m0252(.A(mai_mai_n131_), .B(mai_mai_n280_), .C(l), .Y(mai_mai_n281_));
  NAi31      m0253(.An(e), .B(d), .C(a), .Y(mai_mai_n282_));
  NA2        m0254(.A(mai_mai_n281_), .B(mai_mai_n129_), .Y(mai_mai_n283_));
  INV        m0255(.A(mai_mai_n283_), .Y(mai_mai_n284_));
  NA4        m0256(.A(mai_mai_n159_), .B(mai_mai_n79_), .C(mai_mai_n75_), .D(mai_mai_n118_), .Y(mai_mai_n285_));
  NA3        m0257(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(mai_mai_n83_), .Y(mai_mai_n286_));
  NO2        m0258(.A(mai_mai_n286_), .B(mai_mai_n196_), .Y(mai_mai_n287_));
  NOi21      m0259(.An(mai_mai_n285_), .B(mai_mai_n287_), .Y(mai_mai_n288_));
  NA3        m0260(.A(e), .B(c), .C(b), .Y(mai_mai_n289_));
  NAi21      m0261(.An(l), .B(k), .Y(mai_mai_n290_));
  NO2        m0262(.A(mai_mai_n290_), .B(mai_mai_n49_), .Y(mai_mai_n291_));
  NOi21      m0263(.An(l), .B(j), .Y(mai_mai_n292_));
  NA2        m0264(.A(mai_mai_n162_), .B(mai_mai_n292_), .Y(mai_mai_n293_));
  NA3        m0265(.A(mai_mai_n119_), .B(mai_mai_n118_), .C(m), .Y(mai_mai_n294_));
  OR3        m0266(.A(mai_mai_n70_), .B(mai_mai_n72_), .C(e), .Y(mai_mai_n295_));
  AOI210     m0267(.A0(mai_mai_n294_), .A1(mai_mai_n293_), .B0(mai_mai_n295_), .Y(mai_mai_n296_));
  INV        m0268(.A(mai_mai_n296_), .Y(mai_mai_n297_));
  NAi32      m0269(.An(j), .Bn(h), .C(i), .Y(mai_mai_n298_));
  NAi21      m0270(.An(m), .B(l), .Y(mai_mai_n299_));
  NO3        m0271(.A(mai_mai_n299_), .B(mai_mai_n298_), .C(mai_mai_n83_), .Y(mai_mai_n300_));
  NA2        m0272(.A(h), .B(m), .Y(mai_mai_n301_));
  NA2        m0273(.A(mai_mai_n300_), .B(mai_mai_n163_), .Y(mai_mai_n302_));
  NA3        m0274(.A(mai_mai_n302_), .B(mai_mai_n297_), .C(mai_mai_n288_), .Y(mai_mai_n303_));
  NO2        m0275(.A(mai_mai_n144_), .B(d), .Y(mai_mai_n304_));
  NA2        m0276(.A(mai_mai_n304_), .B(mai_mai_n53_), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n106_), .B(mai_mai_n103_), .Y(mai_mai_n306_));
  NAi32      m0278(.An(n), .Bn(m), .C(l), .Y(mai_mai_n307_));
  NO2        m0279(.A(mai_mai_n307_), .B(mai_mai_n298_), .Y(mai_mai_n308_));
  NA2        m0280(.A(mai_mai_n308_), .B(mai_mai_n185_), .Y(mai_mai_n309_));
  NAi31      m0281(.An(k), .B(l), .C(j), .Y(mai_mai_n310_));
  OAI210     m0282(.A0(mai_mai_n290_), .A1(j), .B0(mai_mai_n310_), .Y(mai_mai_n311_));
  NOi21      m0283(.An(mai_mai_n311_), .B(mai_mai_n121_), .Y(mai_mai_n312_));
  NA2        m0284(.A(mai_mai_n309_), .B(mai_mai_n305_), .Y(mai_mai_n313_));
  NO4        m0285(.A(mai_mai_n313_), .B(mai_mai_n303_), .C(mai_mai_n284_), .D(mai_mai_n276_), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n260_), .B(mai_mai_n195_), .Y(mai_mai_n315_));
  NAi21      m0287(.An(m), .B(k), .Y(mai_mai_n316_));
  NO2        m0288(.A(mai_mai_n229_), .B(mai_mai_n316_), .Y(mai_mai_n317_));
  NAi41      m0289(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n318_));
  NO2        m0290(.A(mai_mai_n318_), .B(mai_mai_n150_), .Y(mai_mai_n319_));
  NA2        m0291(.A(mai_mai_n319_), .B(mai_mai_n317_), .Y(mai_mai_n320_));
  NAi31      m0292(.An(i), .B(l), .C(h), .Y(mai_mai_n321_));
  NO4        m0293(.A(mai_mai_n321_), .B(mai_mai_n150_), .C(mai_mai_n70_), .D(mai_mai_n72_), .Y(mai_mai_n322_));
  NA2        m0294(.A(e), .B(c), .Y(mai_mai_n323_));
  NO3        m0295(.A(mai_mai_n323_), .B(n), .C(d), .Y(mai_mai_n324_));
  NOi21      m0296(.An(f), .B(h), .Y(mai_mai_n325_));
  NA2        m0297(.A(mai_mai_n325_), .B(mai_mai_n119_), .Y(mai_mai_n326_));
  NO2        m0298(.A(mai_mai_n326_), .B(mai_mai_n217_), .Y(mai_mai_n327_));
  NAi31      m0299(.An(d), .B(e), .C(b), .Y(mai_mai_n328_));
  NO2        m0300(.A(mai_mai_n131_), .B(mai_mai_n328_), .Y(mai_mai_n329_));
  NA2        m0301(.A(mai_mai_n329_), .B(mai_mai_n327_), .Y(mai_mai_n330_));
  NAi41      m0302(.An(mai_mai_n322_), .B(mai_mai_n330_), .C(mai_mai_n320_), .D(mai_mai_n315_), .Y(mai_mai_n331_));
  NO4        m0303(.A(mai_mai_n318_), .B(mai_mai_n78_), .C(mai_mai_n69_), .D(mai_mai_n217_), .Y(mai_mai_n332_));
  NA2        m0304(.A(mai_mai_n255_), .B(mai_mai_n104_), .Y(mai_mai_n333_));
  OR2        m0305(.A(mai_mai_n333_), .B(mai_mai_n207_), .Y(mai_mai_n334_));
  NOi31      m0306(.An(l), .B(n), .C(m), .Y(mai_mai_n335_));
  NA2        m0307(.A(mai_mai_n335_), .B(mai_mai_n218_), .Y(mai_mai_n336_));
  NO2        m0308(.A(mai_mai_n336_), .B(mai_mai_n196_), .Y(mai_mai_n337_));
  NAi32      m0309(.An(mai_mai_n337_), .Bn(mai_mai_n332_), .C(mai_mai_n334_), .Y(mai_mai_n338_));
  NAi32      m0310(.An(m), .Bn(j), .C(k), .Y(mai_mai_n339_));
  NAi41      m0311(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n340_));
  OAI210     m0312(.A0(mai_mai_n214_), .A1(mai_mai_n339_), .B0(mai_mai_n340_), .Y(mai_mai_n341_));
  NOi31      m0313(.An(j), .B(m), .C(k), .Y(mai_mai_n342_));
  NO2        m0314(.A(mai_mai_n127_), .B(mai_mai_n342_), .Y(mai_mai_n343_));
  AN3        m0315(.A(h), .B(m), .C(f), .Y(mai_mai_n344_));
  NAi31      m0316(.An(mai_mai_n343_), .B(mai_mai_n344_), .C(mai_mai_n341_), .Y(mai_mai_n345_));
  NOi32      m0317(.An(m), .Bn(j), .C(l), .Y(mai_mai_n346_));
  NO2        m0318(.A(mai_mai_n346_), .B(mai_mai_n97_), .Y(mai_mai_n347_));
  NAi32      m0319(.An(mai_mai_n347_), .Bn(mai_mai_n204_), .C(mai_mai_n304_), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n299_), .B(mai_mai_n298_), .Y(mai_mai_n349_));
  NO2        m0321(.A(mai_mai_n220_), .B(m), .Y(mai_mai_n350_));
  NA2        m0322(.A(mai_mai_n252_), .B(mai_mai_n349_), .Y(mai_mai_n351_));
  NA2        m0323(.A(mai_mai_n237_), .B(mai_mai_n78_), .Y(mai_mai_n352_));
  NA3        m0324(.A(mai_mai_n352_), .B(mai_mai_n344_), .C(mai_mai_n215_), .Y(mai_mai_n353_));
  NA4        m0325(.A(mai_mai_n353_), .B(mai_mai_n351_), .C(mai_mai_n348_), .D(mai_mai_n345_), .Y(mai_mai_n354_));
  NA3        m0326(.A(h), .B(m), .C(f), .Y(mai_mai_n355_));
  NO2        m0327(.A(mai_mai_n355_), .B(mai_mai_n74_), .Y(mai_mai_n356_));
  NA2        m0328(.A(mai_mai_n340_), .B(mai_mai_n214_), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n162_), .B(e), .Y(mai_mai_n358_));
  NO2        m0330(.A(mai_mai_n358_), .B(mai_mai_n41_), .Y(mai_mai_n359_));
  NA2        m0331(.A(mai_mai_n357_), .B(mai_mai_n356_), .Y(mai_mai_n360_));
  NOi32      m0332(.An(j), .Bn(m), .C(i), .Y(mai_mai_n361_));
  NA3        m0333(.A(mai_mai_n361_), .B(mai_mai_n290_), .C(mai_mai_n114_), .Y(mai_mai_n362_));
  AO210      m0334(.A0(mai_mai_n112_), .A1(mai_mai_n32_), .B0(mai_mai_n362_), .Y(mai_mai_n363_));
  NOi32      m0335(.An(e), .Bn(b), .C(a), .Y(mai_mai_n364_));
  AN2        m0336(.A(l), .B(j), .Y(mai_mai_n365_));
  NO2        m0337(.A(mai_mai_n316_), .B(mai_mai_n365_), .Y(mai_mai_n366_));
  NO3        m0338(.A(mai_mai_n318_), .B(mai_mai_n69_), .C(mai_mai_n217_), .Y(mai_mai_n367_));
  NA2        m0339(.A(mai_mai_n211_), .B(mai_mai_n35_), .Y(mai_mai_n368_));
  AOI220     m0340(.A0(mai_mai_n368_), .A1(mai_mai_n364_), .B0(mai_mai_n367_), .B1(mai_mai_n366_), .Y(mai_mai_n369_));
  NA2        m0341(.A(mai_mai_n210_), .B(k), .Y(mai_mai_n370_));
  NA3        m0342(.A(m), .B(mai_mai_n113_), .C(mai_mai_n216_), .Y(mai_mai_n371_));
  NA4        m0343(.A(mai_mai_n206_), .B(mai_mai_n86_), .C(m), .D(mai_mai_n216_), .Y(mai_mai_n372_));
  NAi41      m0344(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n373_));
  NA2        m0345(.A(mai_mai_n51_), .B(mai_mai_n114_), .Y(mai_mai_n374_));
  NA3        m0346(.A(mai_mai_n369_), .B(mai_mai_n363_), .C(mai_mai_n360_), .Y(mai_mai_n375_));
  NO4        m0347(.A(mai_mai_n375_), .B(mai_mai_n354_), .C(mai_mai_n338_), .D(mai_mai_n331_), .Y(mai_mai_n376_));
  NA4        m0348(.A(mai_mai_n376_), .B(mai_mai_n314_), .C(mai_mai_n274_), .D(mai_mai_n202_), .Y(mai10));
  NA3        m0349(.A(m), .B(k), .C(i), .Y(mai_mai_n378_));
  NO3        m0350(.A(mai_mai_n378_), .B(j), .C(mai_mai_n217_), .Y(mai_mai_n379_));
  NOi21      m0351(.An(e), .B(f), .Y(mai_mai_n380_));
  NO4        m0352(.A(mai_mai_n151_), .B(mai_mai_n380_), .C(n), .D(mai_mai_n111_), .Y(mai_mai_n381_));
  NAi31      m0353(.An(b), .B(f), .C(c), .Y(mai_mai_n382_));
  INV        m0354(.A(mai_mai_n382_), .Y(mai_mai_n383_));
  NOi32      m0355(.An(k), .Bn(h), .C(j), .Y(mai_mai_n384_));
  NA2        m0356(.A(mai_mai_n384_), .B(mai_mai_n224_), .Y(mai_mai_n385_));
  NA2        m0357(.A(mai_mai_n160_), .B(mai_mai_n385_), .Y(mai_mai_n386_));
  AOI220     m0358(.A0(mai_mai_n386_), .A1(mai_mai_n383_), .B0(mai_mai_n381_), .B1(mai_mai_n379_), .Y(mai_mai_n387_));
  AN2        m0359(.A(j), .B(h), .Y(mai_mai_n388_));
  NO3        m0360(.A(n), .B(m), .C(k), .Y(mai_mai_n389_));
  NA2        m0361(.A(mai_mai_n389_), .B(mai_mai_n388_), .Y(mai_mai_n390_));
  NO3        m0362(.A(mai_mai_n390_), .B(mai_mai_n151_), .C(mai_mai_n216_), .Y(mai_mai_n391_));
  OR2        m0363(.A(m), .B(k), .Y(mai_mai_n392_));
  NO2        m0364(.A(mai_mai_n175_), .B(mai_mai_n392_), .Y(mai_mai_n393_));
  NA4        m0365(.A(n), .B(f), .C(c), .D(mai_mai_n117_), .Y(mai_mai_n394_));
  NOi21      m0366(.An(mai_mai_n393_), .B(mai_mai_n394_), .Y(mai_mai_n395_));
  NOi32      m0367(.An(d), .Bn(a), .C(c), .Y(mai_mai_n396_));
  NA2        m0368(.A(mai_mai_n396_), .B(mai_mai_n183_), .Y(mai_mai_n397_));
  NAi21      m0369(.An(i), .B(m), .Y(mai_mai_n398_));
  NAi31      m0370(.An(k), .B(m), .C(j), .Y(mai_mai_n399_));
  NO3        m0371(.A(mai_mai_n399_), .B(mai_mai_n398_), .C(n), .Y(mai_mai_n400_));
  NO2        m0372(.A(mai_mai_n395_), .B(mai_mai_n391_), .Y(mai_mai_n401_));
  NO2        m0373(.A(mai_mai_n394_), .B(mai_mai_n299_), .Y(mai_mai_n402_));
  NOi32      m0374(.An(f), .Bn(d), .C(c), .Y(mai_mai_n403_));
  AOI220     m0375(.A0(mai_mai_n403_), .A1(mai_mai_n308_), .B0(mai_mai_n402_), .B1(mai_mai_n218_), .Y(mai_mai_n404_));
  NA3        m0376(.A(mai_mai_n404_), .B(mai_mai_n401_), .C(mai_mai_n387_), .Y(mai_mai_n405_));
  NO2        m0377(.A(mai_mai_n59_), .B(mai_mai_n117_), .Y(mai_mai_n406_));
  NA2        m0378(.A(mai_mai_n255_), .B(mai_mai_n406_), .Y(mai_mai_n407_));
  INV        m0379(.A(e), .Y(mai_mai_n408_));
  NA2        m0380(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n409_));
  OAI220     m0381(.A0(mai_mai_n409_), .A1(mai_mai_n203_), .B0(mai_mai_n207_), .B1(mai_mai_n408_), .Y(mai_mai_n410_));
  AN2        m0382(.A(m), .B(e), .Y(mai_mai_n411_));
  NA3        m0383(.A(mai_mai_n411_), .B(mai_mai_n206_), .C(i), .Y(mai_mai_n412_));
  INV        m0384(.A(mai_mai_n412_), .Y(mai_mai_n413_));
  NO2        m0385(.A(mai_mai_n100_), .B(mai_mai_n408_), .Y(mai_mai_n414_));
  NO3        m0386(.A(mai_mai_n414_), .B(mai_mai_n413_), .C(mai_mai_n410_), .Y(mai_mai_n415_));
  NOi32      m0387(.An(h), .Bn(e), .C(m), .Y(mai_mai_n416_));
  NA3        m0388(.A(mai_mai_n416_), .B(mai_mai_n292_), .C(m), .Y(mai_mai_n417_));
  NOi21      m0389(.An(m), .B(h), .Y(mai_mai_n418_));
  AN3        m0390(.A(m), .B(l), .C(i), .Y(mai_mai_n419_));
  NA3        m0391(.A(mai_mai_n419_), .B(mai_mai_n418_), .C(e), .Y(mai_mai_n420_));
  AN3        m0392(.A(h), .B(m), .C(e), .Y(mai_mai_n421_));
  NA2        m0393(.A(mai_mai_n421_), .B(mai_mai_n97_), .Y(mai_mai_n422_));
  AN3        m0394(.A(mai_mai_n422_), .B(mai_mai_n420_), .C(mai_mai_n417_), .Y(mai_mai_n423_));
  AOI210     m0395(.A0(mai_mai_n423_), .A1(mai_mai_n415_), .B0(mai_mai_n407_), .Y(mai_mai_n424_));
  NA3        m0396(.A(mai_mai_n396_), .B(mai_mai_n183_), .C(mai_mai_n83_), .Y(mai_mai_n425_));
  NAi31      m0397(.An(b), .B(c), .C(a), .Y(mai_mai_n426_));
  NO2        m0398(.A(mai_mai_n426_), .B(n), .Y(mai_mai_n427_));
  NA2        m0399(.A(mai_mai_n51_), .B(m), .Y(mai_mai_n428_));
  NO2        m0400(.A(mai_mai_n428_), .B(mai_mai_n147_), .Y(mai_mai_n429_));
  NA2        m0401(.A(mai_mai_n429_), .B(mai_mai_n427_), .Y(mai_mai_n430_));
  INV        m0402(.A(mai_mai_n430_), .Y(mai_mai_n431_));
  NO3        m0403(.A(mai_mai_n431_), .B(mai_mai_n424_), .C(mai_mai_n405_), .Y(mai_mai_n432_));
  NA2        m0404(.A(i), .B(m), .Y(mai_mai_n433_));
  NOi21      m0405(.An(a), .B(n), .Y(mai_mai_n434_));
  NOi21      m0406(.An(d), .B(c), .Y(mai_mai_n435_));
  NA2        m0407(.A(mai_mai_n435_), .B(mai_mai_n434_), .Y(mai_mai_n436_));
  NA3        m0408(.A(i), .B(m), .C(f), .Y(mai_mai_n437_));
  OR2        m0409(.A(mai_mai_n437_), .B(mai_mai_n68_), .Y(mai_mai_n438_));
  NA3        m0410(.A(mai_mai_n419_), .B(mai_mai_n418_), .C(mai_mai_n183_), .Y(mai_mai_n439_));
  AOI210     m0411(.A0(mai_mai_n439_), .A1(mai_mai_n438_), .B0(mai_mai_n436_), .Y(mai_mai_n440_));
  INV        m0412(.A(mai_mai_n440_), .Y(mai_mai_n441_));
  OR2        m0413(.A(n), .B(m), .Y(mai_mai_n442_));
  NO2        m0414(.A(mai_mai_n442_), .B(mai_mai_n152_), .Y(mai_mai_n443_));
  NO2        m0415(.A(mai_mai_n184_), .B(mai_mai_n147_), .Y(mai_mai_n444_));
  OAI210     m0416(.A0(mai_mai_n443_), .A1(mai_mai_n177_), .B0(mai_mai_n444_), .Y(mai_mai_n445_));
  INV        m0417(.A(mai_mai_n374_), .Y(mai_mai_n446_));
  NA3        m0418(.A(mai_mai_n446_), .B(mai_mai_n364_), .C(d), .Y(mai_mai_n447_));
  NO2        m0419(.A(mai_mai_n426_), .B(mai_mai_n49_), .Y(mai_mai_n448_));
  NO3        m0420(.A(mai_mai_n63_), .B(mai_mai_n113_), .C(e), .Y(mai_mai_n449_));
  NAi21      m0421(.An(k), .B(j), .Y(mai_mai_n450_));
  NA2        m0422(.A(mai_mai_n258_), .B(mai_mai_n450_), .Y(mai_mai_n451_));
  NA3        m0423(.A(mai_mai_n451_), .B(mai_mai_n449_), .C(mai_mai_n448_), .Y(mai_mai_n452_));
  NAi21      m0424(.An(e), .B(d), .Y(mai_mai_n453_));
  INV        m0425(.A(mai_mai_n453_), .Y(mai_mai_n454_));
  NO2        m0426(.A(mai_mai_n259_), .B(mai_mai_n216_), .Y(mai_mai_n455_));
  NA3        m0427(.A(mai_mai_n455_), .B(mai_mai_n454_), .C(mai_mai_n230_), .Y(mai_mai_n456_));
  NA4        m0428(.A(mai_mai_n456_), .B(mai_mai_n452_), .C(mai_mai_n447_), .D(mai_mai_n445_), .Y(mai_mai_n457_));
  NO2        m0429(.A(mai_mai_n336_), .B(mai_mai_n216_), .Y(mai_mai_n458_));
  NA2        m0430(.A(mai_mai_n458_), .B(mai_mai_n454_), .Y(mai_mai_n459_));
  NOi31      m0431(.An(n), .B(m), .C(k), .Y(mai_mai_n460_));
  AOI220     m0432(.A0(mai_mai_n460_), .A1(mai_mai_n388_), .B0(mai_mai_n224_), .B1(mai_mai_n50_), .Y(mai_mai_n461_));
  NAi31      m0433(.An(m), .B(f), .C(c), .Y(mai_mai_n462_));
  OR3        m0434(.A(mai_mai_n462_), .B(mai_mai_n461_), .C(e), .Y(mai_mai_n463_));
  NA3        m0435(.A(mai_mai_n463_), .B(mai_mai_n459_), .C(mai_mai_n309_), .Y(mai_mai_n464_));
  NOi41      m0436(.An(mai_mai_n441_), .B(mai_mai_n464_), .C(mai_mai_n457_), .D(mai_mai_n273_), .Y(mai_mai_n465_));
  NOi32      m0437(.An(c), .Bn(a), .C(b), .Y(mai_mai_n466_));
  NA2        m0438(.A(mai_mai_n466_), .B(mai_mai_n114_), .Y(mai_mai_n467_));
  INV        m0439(.A(mai_mai_n280_), .Y(mai_mai_n468_));
  AN2        m0440(.A(e), .B(d), .Y(mai_mai_n469_));
  NA2        m0441(.A(mai_mai_n469_), .B(mai_mai_n468_), .Y(mai_mai_n470_));
  INV        m0442(.A(mai_mai_n147_), .Y(mai_mai_n471_));
  NO2        m0443(.A(mai_mai_n130_), .B(mai_mai_n41_), .Y(mai_mai_n472_));
  NO2        m0444(.A(mai_mai_n63_), .B(e), .Y(mai_mai_n473_));
  NA4        m0445(.A(mai_mai_n321_), .B(mai_mai_n165_), .C(mai_mai_n267_), .D(mai_mai_n120_), .Y(mai_mai_n474_));
  AOI220     m0446(.A0(mai_mai_n474_), .A1(mai_mai_n473_), .B0(mai_mai_n472_), .B1(mai_mai_n471_), .Y(mai_mai_n475_));
  AOI210     m0447(.A0(mai_mai_n475_), .A1(mai_mai_n470_), .B0(mai_mai_n467_), .Y(mai_mai_n476_));
  NO2        m0448(.A(mai_mai_n212_), .B(mai_mai_n208_), .Y(mai_mai_n477_));
  NOi21      m0449(.An(a), .B(b), .Y(mai_mai_n478_));
  NA3        m0450(.A(e), .B(d), .C(c), .Y(mai_mai_n479_));
  NAi21      m0451(.An(mai_mai_n479_), .B(mai_mai_n478_), .Y(mai_mai_n480_));
  NO2        m0452(.A(mai_mai_n425_), .B(mai_mai_n207_), .Y(mai_mai_n481_));
  NOi21      m0453(.An(mai_mai_n480_), .B(mai_mai_n481_), .Y(mai_mai_n482_));
  AOI210     m0454(.A0(mai_mai_n275_), .A1(mai_mai_n477_), .B0(mai_mai_n482_), .Y(mai_mai_n483_));
  NO4        m0455(.A(mai_mai_n190_), .B(mai_mai_n103_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n484_));
  NA2        m0456(.A(mai_mai_n383_), .B(mai_mai_n153_), .Y(mai_mai_n485_));
  OR2        m0457(.A(k), .B(j), .Y(mai_mai_n486_));
  NA2        m0458(.A(l), .B(k), .Y(mai_mai_n487_));
  NA3        m0459(.A(mai_mai_n487_), .B(mai_mai_n486_), .C(mai_mai_n224_), .Y(mai_mai_n488_));
  AOI210     m0460(.A0(mai_mai_n237_), .A1(mai_mai_n339_), .B0(mai_mai_n83_), .Y(mai_mai_n489_));
  NOi21      m0461(.An(mai_mai_n488_), .B(mai_mai_n489_), .Y(mai_mai_n490_));
  OR3        m0462(.A(mai_mai_n490_), .B(mai_mai_n143_), .C(mai_mai_n134_), .Y(mai_mai_n491_));
  INV        m0463(.A(mai_mai_n285_), .Y(mai_mai_n492_));
  NO3        m0464(.A(mai_mai_n425_), .B(mai_mai_n91_), .C(mai_mai_n130_), .Y(mai_mai_n493_));
  NO3        m0465(.A(mai_mai_n493_), .B(mai_mai_n492_), .C(mai_mai_n322_), .Y(mai_mai_n494_));
  NA3        m0466(.A(mai_mai_n494_), .B(mai_mai_n491_), .C(mai_mai_n485_), .Y(mai_mai_n495_));
  NO4        m0467(.A(mai_mai_n495_), .B(mai_mai_n484_), .C(mai_mai_n483_), .D(mai_mai_n476_), .Y(mai_mai_n496_));
  NA2        m0468(.A(mai_mai_n67_), .B(mai_mai_n64_), .Y(mai_mai_n497_));
  NOi21      m0469(.An(d), .B(e), .Y(mai_mai_n498_));
  NO2        m0470(.A(mai_mai_n190_), .B(mai_mai_n56_), .Y(mai_mai_n499_));
  NAi31      m0471(.An(j), .B(l), .C(i), .Y(mai_mai_n500_));
  OAI210     m0472(.A0(mai_mai_n500_), .A1(mai_mai_n131_), .B0(mai_mai_n103_), .Y(mai_mai_n501_));
  NA3        m0473(.A(mai_mai_n501_), .B(mai_mai_n499_), .C(mai_mai_n498_), .Y(mai_mai_n502_));
  NO3        m0474(.A(mai_mai_n397_), .B(mai_mai_n347_), .C(mai_mai_n204_), .Y(mai_mai_n503_));
  NO2        m0475(.A(mai_mai_n397_), .B(mai_mai_n374_), .Y(mai_mai_n504_));
  NO4        m0476(.A(mai_mai_n504_), .B(mai_mai_n503_), .C(mai_mai_n186_), .D(mai_mai_n306_), .Y(mai_mai_n505_));
  NA4        m0477(.A(mai_mai_n505_), .B(mai_mai_n502_), .C(mai_mai_n497_), .D(mai_mai_n247_), .Y(mai_mai_n506_));
  OAI210     m0478(.A0(mai_mai_n128_), .A1(mai_mai_n127_), .B0(n), .Y(mai_mai_n507_));
  NO2        m0479(.A(mai_mai_n507_), .B(mai_mai_n130_), .Y(mai_mai_n508_));
  BUFFER     m0480(.A(mai_mai_n249_), .Y(mai_mai_n509_));
  OA210      m0481(.A0(mai_mai_n509_), .A1(mai_mai_n508_), .B0(mai_mai_n195_), .Y(mai_mai_n510_));
  XO2        m0482(.A(i), .B(h), .Y(mai_mai_n511_));
  NA3        m0483(.A(mai_mai_n511_), .B(mai_mai_n159_), .C(n), .Y(mai_mai_n512_));
  NAi41      m0484(.An(mai_mai_n300_), .B(mai_mai_n512_), .C(mai_mai_n461_), .D(mai_mai_n385_), .Y(mai_mai_n513_));
  NOi32      m0485(.An(mai_mai_n513_), .Bn(mai_mai_n473_), .C(mai_mai_n277_), .Y(mai_mai_n514_));
  NAi31      m0486(.An(c), .B(f), .C(d), .Y(mai_mai_n515_));
  AOI210     m0487(.A0(mai_mai_n286_), .A1(mai_mai_n198_), .B0(mai_mai_n515_), .Y(mai_mai_n516_));
  NOi21      m0488(.An(mai_mai_n81_), .B(mai_mai_n516_), .Y(mai_mai_n517_));
  NA3        m0489(.A(mai_mai_n381_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n518_));
  NA2        m0490(.A(mai_mai_n231_), .B(mai_mai_n109_), .Y(mai_mai_n519_));
  AOI210     m0491(.A0(mai_mai_n519_), .A1(mai_mai_n182_), .B0(mai_mai_n515_), .Y(mai_mai_n520_));
  AOI210     m0492(.A0(mai_mai_n362_), .A1(mai_mai_n35_), .B0(mai_mai_n480_), .Y(mai_mai_n521_));
  NOi31      m0493(.An(mai_mai_n518_), .B(mai_mai_n521_), .C(mai_mai_n520_), .Y(mai_mai_n522_));
  AN2        m0494(.A(mai_mai_n166_), .B(mai_mai_n64_), .Y(mai_mai_n523_));
  NA3        m0495(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n524_));
  NO2        m0496(.A(mai_mai_n524_), .B(mai_mai_n436_), .Y(mai_mai_n525_));
  NO2        m0497(.A(mai_mai_n525_), .B(mai_mai_n296_), .Y(mai_mai_n526_));
  NAi41      m0498(.An(mai_mai_n523_), .B(mai_mai_n526_), .C(mai_mai_n522_), .D(mai_mai_n517_), .Y(mai_mai_n527_));
  NO4        m0499(.A(mai_mai_n527_), .B(mai_mai_n514_), .C(mai_mai_n510_), .D(mai_mai_n506_), .Y(mai_mai_n528_));
  NA4        m0500(.A(mai_mai_n528_), .B(mai_mai_n496_), .C(mai_mai_n465_), .D(mai_mai_n432_), .Y(mai11));
  NO2        m0501(.A(mai_mai_n70_), .B(f), .Y(mai_mai_n530_));
  NA2        m0502(.A(j), .B(m), .Y(mai_mai_n531_));
  NAi31      m0503(.An(i), .B(m), .C(l), .Y(mai_mai_n532_));
  NA3        m0504(.A(m), .B(k), .C(j), .Y(mai_mai_n533_));
  OAI220     m0505(.A0(mai_mai_n533_), .A1(mai_mai_n130_), .B0(mai_mai_n532_), .B1(mai_mai_n531_), .Y(mai_mai_n534_));
  NA2        m0506(.A(mai_mai_n534_), .B(mai_mai_n530_), .Y(mai_mai_n535_));
  NOi32      m0507(.An(e), .Bn(b), .C(f), .Y(mai_mai_n536_));
  NA2        m0508(.A(mai_mai_n266_), .B(mai_mai_n114_), .Y(mai_mai_n537_));
  NA2        m0509(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n538_));
  NAi31      m0510(.An(d), .B(e), .C(a), .Y(mai_mai_n539_));
  NO2        m0511(.A(mai_mai_n539_), .B(n), .Y(mai_mai_n540_));
  NA2        m0512(.A(mai_mai_n540_), .B(mai_mai_n101_), .Y(mai_mai_n541_));
  NAi41      m0513(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n542_));
  AN2        m0514(.A(mai_mai_n542_), .B(mai_mai_n373_), .Y(mai_mai_n543_));
  AOI210     m0515(.A0(mai_mai_n543_), .A1(mai_mai_n397_), .B0(mai_mai_n278_), .Y(mai_mai_n544_));
  NA2        m0516(.A(j), .B(i), .Y(mai_mai_n545_));
  NAi31      m0517(.An(n), .B(m), .C(k), .Y(mai_mai_n546_));
  NO3        m0518(.A(mai_mai_n546_), .B(mai_mai_n545_), .C(mai_mai_n113_), .Y(mai_mai_n547_));
  NO4        m0519(.A(n), .B(d), .C(mai_mai_n117_), .D(a), .Y(mai_mai_n548_));
  OR2        m0520(.A(n), .B(c), .Y(mai_mai_n549_));
  NO2        m0521(.A(mai_mai_n549_), .B(mai_mai_n149_), .Y(mai_mai_n550_));
  NO2        m0522(.A(mai_mai_n550_), .B(mai_mai_n548_), .Y(mai_mai_n551_));
  NOi32      m0523(.An(m), .Bn(f), .C(i), .Y(mai_mai_n552_));
  NA2        m0524(.A(mai_mai_n534_), .B(f), .Y(mai_mai_n553_));
  NO2        m0525(.A(mai_mai_n280_), .B(mai_mai_n49_), .Y(mai_mai_n554_));
  NO2        m0526(.A(mai_mai_n553_), .B(mai_mai_n551_), .Y(mai_mai_n555_));
  AOI210     m0527(.A0(mai_mai_n547_), .A1(mai_mai_n544_), .B0(mai_mai_n555_), .Y(mai_mai_n556_));
  NA2        m0528(.A(mai_mai_n139_), .B(mai_mai_n34_), .Y(mai_mai_n557_));
  OAI220     m0529(.A0(mai_mai_n557_), .A1(m), .B0(mai_mai_n538_), .B1(mai_mai_n237_), .Y(mai_mai_n558_));
  NOi41      m0530(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n559_));
  NAi32      m0531(.An(e), .Bn(b), .C(c), .Y(mai_mai_n560_));
  OR2        m0532(.A(mai_mai_n560_), .B(mai_mai_n83_), .Y(mai_mai_n561_));
  AN2        m0533(.A(mai_mai_n340_), .B(mai_mai_n318_), .Y(mai_mai_n562_));
  NA2        m0534(.A(mai_mai_n562_), .B(mai_mai_n561_), .Y(mai_mai_n563_));
  OA210      m0535(.A0(mai_mai_n563_), .A1(mai_mai_n559_), .B0(mai_mai_n558_), .Y(mai_mai_n564_));
  OAI220     m0536(.A0(mai_mai_n399_), .A1(mai_mai_n398_), .B0(mai_mai_n532_), .B1(mai_mai_n531_), .Y(mai_mai_n565_));
  NO3        m0537(.A(mai_mai_n61_), .B(mai_mai_n49_), .C(mai_mai_n217_), .Y(mai_mai_n566_));
  NO2        m0538(.A(mai_mai_n234_), .B(mai_mai_n111_), .Y(mai_mai_n567_));
  OAI210     m0539(.A0(mai_mai_n566_), .A1(mai_mai_n400_), .B0(mai_mai_n567_), .Y(mai_mai_n568_));
  INV        m0540(.A(mai_mai_n568_), .Y(mai_mai_n569_));
  NO2        m0541(.A(mai_mai_n282_), .B(n), .Y(mai_mai_n570_));
  NO2        m0542(.A(mai_mai_n427_), .B(mai_mai_n570_), .Y(mai_mai_n571_));
  NA2        m0543(.A(mai_mai_n565_), .B(f), .Y(mai_mai_n572_));
  NAi32      m0544(.An(d), .Bn(a), .C(b), .Y(mai_mai_n573_));
  NO2        m0545(.A(mai_mai_n573_), .B(mai_mai_n49_), .Y(mai_mai_n574_));
  NA2        m0546(.A(h), .B(f), .Y(mai_mai_n575_));
  NO2        m0547(.A(mai_mai_n575_), .B(mai_mai_n94_), .Y(mai_mai_n576_));
  NO3        m0548(.A(mai_mai_n178_), .B(mai_mai_n175_), .C(m), .Y(mai_mai_n577_));
  AOI220     m0549(.A0(mai_mai_n577_), .A1(mai_mai_n58_), .B0(mai_mai_n576_), .B1(mai_mai_n574_), .Y(mai_mai_n578_));
  OAI210     m0550(.A0(mai_mai_n572_), .A1(mai_mai_n571_), .B0(mai_mai_n578_), .Y(mai_mai_n579_));
  AN3        m0551(.A(j), .B(h), .C(m), .Y(mai_mai_n580_));
  NO2        m0552(.A(mai_mai_n146_), .B(c), .Y(mai_mai_n581_));
  NA3        m0553(.A(mai_mai_n581_), .B(mai_mai_n580_), .C(mai_mai_n460_), .Y(mai_mai_n582_));
  NA3        m0554(.A(f), .B(d), .C(b), .Y(mai_mai_n583_));
  NO4        m0555(.A(mai_mai_n583_), .B(mai_mai_n178_), .C(mai_mai_n175_), .D(m), .Y(mai_mai_n584_));
  NAi21      m0556(.An(mai_mai_n584_), .B(mai_mai_n582_), .Y(mai_mai_n585_));
  NO4        m0557(.A(mai_mai_n585_), .B(mai_mai_n579_), .C(mai_mai_n569_), .D(mai_mai_n564_), .Y(mai_mai_n586_));
  AN4        m0558(.A(mai_mai_n586_), .B(mai_mai_n556_), .C(mai_mai_n541_), .D(mai_mai_n535_), .Y(mai_mai_n587_));
  INV        m0559(.A(k), .Y(mai_mai_n588_));
  NA3        m0560(.A(l), .B(mai_mai_n588_), .C(i), .Y(mai_mai_n589_));
  INV        m0561(.A(mai_mai_n589_), .Y(mai_mai_n590_));
  NA4        m0562(.A(mai_mai_n396_), .B(mai_mai_n418_), .C(mai_mai_n183_), .D(mai_mai_n114_), .Y(mai_mai_n591_));
  NAi32      m0563(.An(h), .Bn(f), .C(m), .Y(mai_mai_n592_));
  NAi41      m0564(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n593_));
  OAI210     m0565(.A0(mai_mai_n539_), .A1(n), .B0(mai_mai_n593_), .Y(mai_mai_n594_));
  NA2        m0566(.A(mai_mai_n594_), .B(m), .Y(mai_mai_n595_));
  NAi31      m0567(.An(h), .B(m), .C(f), .Y(mai_mai_n596_));
  OR3        m0568(.A(mai_mai_n596_), .B(mai_mai_n282_), .C(mai_mai_n49_), .Y(mai_mai_n597_));
  NA4        m0569(.A(mai_mai_n418_), .B(mai_mai_n122_), .C(mai_mai_n114_), .D(e), .Y(mai_mai_n598_));
  AN2        m0570(.A(mai_mai_n598_), .B(mai_mai_n597_), .Y(mai_mai_n599_));
  OA210      m0571(.A0(mai_mai_n595_), .A1(mai_mai_n592_), .B0(mai_mai_n599_), .Y(mai_mai_n600_));
  NO3        m0572(.A(mai_mai_n592_), .B(mai_mai_n70_), .C(mai_mai_n72_), .Y(mai_mai_n601_));
  NO4        m0573(.A(mai_mai_n596_), .B(mai_mai_n549_), .C(mai_mai_n149_), .D(mai_mai_n72_), .Y(mai_mai_n602_));
  OR2        m0574(.A(mai_mai_n602_), .B(mai_mai_n601_), .Y(mai_mai_n603_));
  NAi31      m0575(.An(mai_mai_n603_), .B(mai_mai_n600_), .C(mai_mai_n591_), .Y(mai_mai_n604_));
  NAi31      m0576(.An(f), .B(h), .C(m), .Y(mai_mai_n605_));
  NO4        m0577(.A(mai_mai_n310_), .B(mai_mai_n605_), .C(mai_mai_n70_), .D(mai_mai_n72_), .Y(mai_mai_n606_));
  NOi32      m0578(.An(b), .Bn(a), .C(c), .Y(mai_mai_n607_));
  NOi41      m0579(.An(mai_mai_n607_), .B(mai_mai_n355_), .C(mai_mai_n66_), .D(mai_mai_n118_), .Y(mai_mai_n608_));
  OR2        m0580(.A(mai_mai_n608_), .B(mai_mai_n606_), .Y(mai_mai_n609_));
  NOi32      m0581(.An(d), .Bn(a), .C(e), .Y(mai_mai_n610_));
  NA2        m0582(.A(mai_mai_n610_), .B(mai_mai_n114_), .Y(mai_mai_n611_));
  NO2        m0583(.A(n), .B(c), .Y(mai_mai_n612_));
  NA3        m0584(.A(mai_mai_n612_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n613_));
  NAi32      m0585(.An(n), .Bn(f), .C(m), .Y(mai_mai_n614_));
  NA3        m0586(.A(mai_mai_n614_), .B(mai_mai_n613_), .C(mai_mai_n611_), .Y(mai_mai_n615_));
  NOi32      m0587(.An(e), .Bn(a), .C(d), .Y(mai_mai_n616_));
  AOI210     m0588(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n616_), .Y(mai_mai_n617_));
  AOI210     m0589(.A0(mai_mai_n617_), .A1(mai_mai_n216_), .B0(mai_mai_n557_), .Y(mai_mai_n618_));
  AOI210     m0590(.A0(mai_mai_n618_), .A1(mai_mai_n615_), .B0(mai_mai_n609_), .Y(mai_mai_n619_));
  OAI210     m0591(.A0(mai_mai_n254_), .A1(mai_mai_n86_), .B0(mai_mai_n619_), .Y(mai_mai_n620_));
  AOI210     m0592(.A0(mai_mai_n604_), .A1(mai_mai_n590_), .B0(mai_mai_n620_), .Y(mai_mai_n621_));
  NO3        m0593(.A(mai_mai_n316_), .B(mai_mai_n60_), .C(n), .Y(mai_mai_n622_));
  NA3        m0594(.A(mai_mai_n515_), .B(mai_mai_n173_), .C(mai_mai_n172_), .Y(mai_mai_n623_));
  NA2        m0595(.A(mai_mai_n462_), .B(mai_mai_n234_), .Y(mai_mai_n624_));
  OR2        m0596(.A(mai_mai_n624_), .B(mai_mai_n623_), .Y(mai_mai_n625_));
  NA2        m0597(.A(mai_mai_n73_), .B(mai_mai_n114_), .Y(mai_mai_n626_));
  NO2        m0598(.A(mai_mai_n626_), .B(mai_mai_n45_), .Y(mai_mai_n627_));
  AOI220     m0599(.A0(mai_mai_n627_), .A1(mai_mai_n544_), .B0(mai_mai_n625_), .B1(mai_mai_n622_), .Y(mai_mai_n628_));
  NO2        m0600(.A(mai_mai_n628_), .B(mai_mai_n86_), .Y(mai_mai_n629_));
  NA3        m0601(.A(mai_mai_n559_), .B(mai_mai_n342_), .C(mai_mai_n46_), .Y(mai_mai_n630_));
  NOi32      m0602(.An(e), .Bn(c), .C(f), .Y(mai_mai_n631_));
  NOi21      m0603(.An(f), .B(m), .Y(mai_mai_n632_));
  NO2        m0604(.A(mai_mai_n632_), .B(mai_mai_n214_), .Y(mai_mai_n633_));
  AOI220     m0605(.A0(mai_mai_n633_), .A1(mai_mai_n393_), .B0(mai_mai_n631_), .B1(mai_mai_n177_), .Y(mai_mai_n634_));
  NA3        m0606(.A(mai_mai_n634_), .B(mai_mai_n630_), .C(mai_mai_n180_), .Y(mai_mai_n635_));
  NOi21      m0607(.An(j), .B(l), .Y(mai_mai_n636_));
  NAi21      m0608(.An(k), .B(h), .Y(mai_mai_n637_));
  NO2        m0609(.A(mai_mai_n637_), .B(mai_mai_n269_), .Y(mai_mai_n638_));
  NA2        m0610(.A(mai_mai_n638_), .B(mai_mai_n636_), .Y(mai_mai_n639_));
  OR2        m0611(.A(mai_mai_n639_), .B(mai_mai_n595_), .Y(mai_mai_n640_));
  NOi31      m0612(.An(m), .B(n), .C(k), .Y(mai_mai_n641_));
  NA2        m0613(.A(mai_mai_n636_), .B(mai_mai_n641_), .Y(mai_mai_n642_));
  NO2        m0614(.A(mai_mai_n282_), .B(mai_mai_n49_), .Y(mai_mai_n643_));
  NO2        m0615(.A(mai_mai_n310_), .B(mai_mai_n605_), .Y(mai_mai_n644_));
  NO2        m0616(.A(mai_mai_n539_), .B(mai_mai_n49_), .Y(mai_mai_n645_));
  AOI220     m0617(.A0(mai_mai_n645_), .A1(mai_mai_n644_), .B0(mai_mai_n643_), .B1(mai_mai_n576_), .Y(mai_mai_n646_));
  NA2        m0618(.A(mai_mai_n646_), .B(mai_mai_n640_), .Y(mai_mai_n647_));
  NA2        m0619(.A(mai_mai_n109_), .B(mai_mai_n36_), .Y(mai_mai_n648_));
  NO2        m0620(.A(k), .B(mai_mai_n217_), .Y(mai_mai_n649_));
  INV        m0621(.A(mai_mai_n364_), .Y(mai_mai_n650_));
  NO2        m0622(.A(mai_mai_n650_), .B(n), .Y(mai_mai_n651_));
  NAi31      m0623(.An(mai_mai_n648_), .B(mai_mai_n651_), .C(mai_mai_n649_), .Y(mai_mai_n652_));
  NO2        m0624(.A(mai_mai_n538_), .B(mai_mai_n178_), .Y(mai_mai_n653_));
  NA3        m0625(.A(mai_mai_n560_), .B(mai_mai_n277_), .C(mai_mai_n144_), .Y(mai_mai_n654_));
  NA2        m0626(.A(mai_mai_n511_), .B(mai_mai_n159_), .Y(mai_mai_n655_));
  NO3        m0627(.A(mai_mai_n394_), .B(mai_mai_n655_), .C(mai_mai_n86_), .Y(mai_mai_n656_));
  AOI210     m0628(.A0(mai_mai_n654_), .A1(mai_mai_n653_), .B0(mai_mai_n656_), .Y(mai_mai_n657_));
  AN3        m0629(.A(f), .B(d), .C(b), .Y(mai_mai_n658_));
  OAI210     m0630(.A0(mai_mai_n658_), .A1(mai_mai_n129_), .B0(n), .Y(mai_mai_n659_));
  NA3        m0631(.A(mai_mai_n511_), .B(mai_mai_n159_), .C(mai_mai_n217_), .Y(mai_mai_n660_));
  AOI210     m0632(.A0(mai_mai_n659_), .A1(mai_mai_n236_), .B0(mai_mai_n660_), .Y(mai_mai_n661_));
  NAi31      m0633(.An(m), .B(n), .C(k), .Y(mai_mai_n662_));
  INV        m0634(.A(mai_mai_n256_), .Y(mai_mai_n663_));
  OAI210     m0635(.A0(mai_mai_n663_), .A1(mai_mai_n661_), .B0(j), .Y(mai_mai_n664_));
  NA3        m0636(.A(mai_mai_n664_), .B(mai_mai_n657_), .C(mai_mai_n652_), .Y(mai_mai_n665_));
  NO4        m0637(.A(mai_mai_n665_), .B(mai_mai_n647_), .C(mai_mai_n635_), .D(mai_mai_n629_), .Y(mai_mai_n666_));
  NA2        m0638(.A(mai_mai_n381_), .B(mai_mai_n162_), .Y(mai_mai_n667_));
  NAi31      m0639(.An(m), .B(h), .C(f), .Y(mai_mai_n668_));
  OA210      m0640(.A0(mai_mai_n539_), .A1(n), .B0(mai_mai_n593_), .Y(mai_mai_n669_));
  NO2        m0641(.A(mai_mai_n669_), .B(mai_mai_n90_), .Y(mai_mai_n670_));
  INV        m0642(.A(mai_mai_n670_), .Y(mai_mai_n671_));
  AOI210     m0643(.A0(mai_mai_n671_), .A1(mai_mai_n667_), .B0(mai_mai_n533_), .Y(mai_mai_n672_));
  NO3        m0644(.A(m), .B(mai_mai_n216_), .C(mai_mai_n56_), .Y(mai_mai_n673_));
  NAi21      m0645(.An(h), .B(j), .Y(mai_mai_n674_));
  NO2        m0646(.A(mai_mai_n519_), .B(mai_mai_n86_), .Y(mai_mai_n675_));
  OAI210     m0647(.A0(mai_mai_n675_), .A1(mai_mai_n393_), .B0(mai_mai_n673_), .Y(mai_mai_n676_));
  OR2        m0648(.A(mai_mai_n70_), .B(mai_mai_n72_), .Y(mai_mai_n677_));
  NA2        m0649(.A(mai_mai_n607_), .B(mai_mai_n344_), .Y(mai_mai_n678_));
  OA220      m0650(.A0(mai_mai_n642_), .A1(mai_mai_n678_), .B0(mai_mai_n639_), .B1(mai_mai_n677_), .Y(mai_mai_n679_));
  AN2        m0651(.A(h), .B(f), .Y(mai_mai_n680_));
  NA2        m0652(.A(mai_mai_n680_), .B(mai_mai_n37_), .Y(mai_mai_n681_));
  NA2        m0653(.A(mai_mai_n99_), .B(mai_mai_n46_), .Y(mai_mai_n682_));
  OAI220     m0654(.A0(mai_mai_n682_), .A1(mai_mai_n333_), .B0(mai_mai_n681_), .B1(mai_mai_n467_), .Y(mai_mai_n683_));
  AOI210     m0655(.A0(mai_mai_n573_), .A1(mai_mai_n426_), .B0(mai_mai_n49_), .Y(mai_mai_n684_));
  OAI220     m0656(.A0(mai_mai_n596_), .A1(mai_mai_n589_), .B0(mai_mai_n326_), .B1(mai_mai_n531_), .Y(mai_mai_n685_));
  AOI210     m0657(.A0(mai_mai_n685_), .A1(mai_mai_n684_), .B0(mai_mai_n683_), .Y(mai_mai_n686_));
  NA3        m0658(.A(mai_mai_n686_), .B(mai_mai_n679_), .C(mai_mai_n676_), .Y(mai_mai_n687_));
  NO2        m0659(.A(mai_mai_n258_), .B(f), .Y(mai_mai_n688_));
  NO2        m0660(.A(mai_mai_n632_), .B(mai_mai_n60_), .Y(mai_mai_n689_));
  NO3        m0661(.A(mai_mai_n689_), .B(mai_mai_n688_), .C(mai_mai_n34_), .Y(mai_mai_n690_));
  NA2        m0662(.A(mai_mai_n329_), .B(mai_mai_n139_), .Y(mai_mai_n691_));
  NA2        m0663(.A(mai_mai_n131_), .B(mai_mai_n49_), .Y(mai_mai_n692_));
  AOI220     m0664(.A0(mai_mai_n692_), .A1(mai_mai_n536_), .B0(mai_mai_n364_), .B1(mai_mai_n114_), .Y(mai_mai_n693_));
  OA220      m0665(.A0(mai_mai_n693_), .A1(mai_mai_n557_), .B0(mai_mai_n362_), .B1(mai_mai_n112_), .Y(mai_mai_n694_));
  OAI210     m0666(.A0(mai_mai_n691_), .A1(mai_mai_n690_), .B0(mai_mai_n694_), .Y(mai_mai_n695_));
  NO3        m0667(.A(mai_mai_n403_), .B(mai_mai_n195_), .C(mai_mai_n194_), .Y(mai_mai_n696_));
  NA2        m0668(.A(mai_mai_n696_), .B(mai_mai_n234_), .Y(mai_mai_n697_));
  NA3        m0669(.A(mai_mai_n697_), .B(mai_mai_n260_), .C(j), .Y(mai_mai_n698_));
  NO3        m0670(.A(mai_mai_n462_), .B(mai_mai_n175_), .C(i), .Y(mai_mai_n699_));
  NA2        m0671(.A(mai_mai_n466_), .B(mai_mai_n83_), .Y(mai_mai_n700_));
  NO4        m0672(.A(mai_mai_n533_), .B(mai_mai_n700_), .C(mai_mai_n130_), .D(mai_mai_n216_), .Y(mai_mai_n701_));
  INV        m0673(.A(mai_mai_n701_), .Y(mai_mai_n702_));
  NA4        m0674(.A(mai_mai_n702_), .B(mai_mai_n698_), .C(mai_mai_n518_), .D(mai_mai_n401_), .Y(mai_mai_n703_));
  NO4        m0675(.A(mai_mai_n703_), .B(mai_mai_n695_), .C(mai_mai_n687_), .D(mai_mai_n672_), .Y(mai_mai_n704_));
  NA4        m0676(.A(mai_mai_n704_), .B(mai_mai_n666_), .C(mai_mai_n621_), .D(mai_mai_n587_), .Y(mai08));
  NO2        m0677(.A(k), .B(h), .Y(mai_mai_n706_));
  AO210      m0678(.A0(mai_mai_n258_), .A1(mai_mai_n450_), .B0(mai_mai_n706_), .Y(mai_mai_n707_));
  NO2        m0679(.A(mai_mai_n707_), .B(mai_mai_n299_), .Y(mai_mai_n708_));
  NA2        m0680(.A(mai_mai_n631_), .B(mai_mai_n83_), .Y(mai_mai_n709_));
  NA2        m0681(.A(mai_mai_n709_), .B(mai_mai_n462_), .Y(mai_mai_n710_));
  AOI210     m0682(.A0(mai_mai_n710_), .A1(mai_mai_n708_), .B0(mai_mai_n493_), .Y(mai_mai_n711_));
  NA2        m0683(.A(mai_mai_n83_), .B(mai_mai_n111_), .Y(mai_mai_n712_));
  NO2        m0684(.A(mai_mai_n712_), .B(mai_mai_n57_), .Y(mai_mai_n713_));
  NO4        m0685(.A(mai_mai_n378_), .B(mai_mai_n113_), .C(j), .D(mai_mai_n217_), .Y(mai_mai_n714_));
  NA2        m0686(.A(mai_mai_n583_), .B(mai_mai_n236_), .Y(mai_mai_n715_));
  AOI220     m0687(.A0(mai_mai_n715_), .A1(mai_mai_n350_), .B0(mai_mai_n714_), .B1(mai_mai_n713_), .Y(mai_mai_n716_));
  AOI210     m0688(.A0(mai_mai_n583_), .A1(mai_mai_n155_), .B0(mai_mai_n83_), .Y(mai_mai_n717_));
  NA4        m0689(.A(mai_mai_n219_), .B(mai_mai_n139_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n718_));
  AN2        m0690(.A(l), .B(k), .Y(mai_mai_n719_));
  NA4        m0691(.A(mai_mai_n719_), .B(mai_mai_n109_), .C(mai_mai_n72_), .D(mai_mai_n217_), .Y(mai_mai_n720_));
  OAI210     m0692(.A0(mai_mai_n718_), .A1(m), .B0(mai_mai_n720_), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n721_), .B(mai_mai_n717_), .Y(mai_mai_n722_));
  NA4        m0694(.A(mai_mai_n722_), .B(mai_mai_n716_), .C(mai_mai_n711_), .D(mai_mai_n351_), .Y(mai_mai_n723_));
  AN2        m0695(.A(mai_mai_n540_), .B(mai_mai_n95_), .Y(mai_mai_n724_));
  NO4        m0696(.A(mai_mai_n175_), .B(mai_mai_n392_), .C(mai_mai_n113_), .D(m), .Y(mai_mai_n725_));
  AOI210     m0697(.A0(mai_mai_n725_), .A1(mai_mai_n715_), .B0(mai_mai_n525_), .Y(mai_mai_n726_));
  NO2        m0698(.A(mai_mai_n38_), .B(mai_mai_n216_), .Y(mai_mai_n727_));
  AOI220     m0699(.A0(mai_mai_n633_), .A1(mai_mai_n349_), .B0(mai_mai_n727_), .B1(mai_mai_n570_), .Y(mai_mai_n728_));
  NAi31      m0700(.An(mai_mai_n724_), .B(mai_mai_n728_), .C(mai_mai_n726_), .Y(mai_mai_n729_));
  NO2        m0701(.A(mai_mai_n543_), .B(mai_mai_n35_), .Y(mai_mai_n730_));
  INV        m0702(.A(mai_mai_n730_), .Y(mai_mai_n731_));
  NO3        m0703(.A(mai_mai_n316_), .B(mai_mai_n130_), .C(mai_mai_n41_), .Y(mai_mai_n732_));
  NA2        m0704(.A(mai_mai_n707_), .B(mai_mai_n135_), .Y(mai_mai_n733_));
  AOI220     m0705(.A0(mai_mai_n733_), .A1(mai_mai_n402_), .B0(mai_mai_n732_), .B1(mai_mai_n75_), .Y(mai_mai_n734_));
  OAI210     m0706(.A0(mai_mai_n731_), .A1(mai_mai_n86_), .B0(mai_mai_n734_), .Y(mai_mai_n735_));
  NA2        m0707(.A(mai_mai_n364_), .B(mai_mai_n43_), .Y(mai_mai_n736_));
  NA3        m0708(.A(mai_mai_n697_), .B(mai_mai_n335_), .C(mai_mai_n384_), .Y(mai_mai_n737_));
  NA2        m0709(.A(mai_mai_n719_), .B(mai_mai_n224_), .Y(mai_mai_n738_));
  NO2        m0710(.A(mai_mai_n738_), .B(mai_mai_n328_), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n739_), .B(mai_mai_n688_), .Y(mai_mai_n740_));
  NA3        m0712(.A(m), .B(l), .C(k), .Y(mai_mai_n741_));
  NO2        m0713(.A(mai_mai_n542_), .B(mai_mai_n278_), .Y(mai_mai_n742_));
  NOi21      m0714(.An(mai_mai_n742_), .B(mai_mai_n537_), .Y(mai_mai_n743_));
  NA4        m0715(.A(mai_mai_n114_), .B(l), .C(k), .D(mai_mai_n86_), .Y(mai_mai_n744_));
  NA3        m0716(.A(mai_mai_n122_), .B(mai_mai_n411_), .C(i), .Y(mai_mai_n745_));
  NO2        m0717(.A(mai_mai_n745_), .B(mai_mai_n744_), .Y(mai_mai_n746_));
  NO2        m0718(.A(mai_mai_n746_), .B(mai_mai_n743_), .Y(mai_mai_n747_));
  NA4        m0719(.A(mai_mai_n747_), .B(mai_mai_n740_), .C(mai_mai_n737_), .D(mai_mai_n736_), .Y(mai_mai_n748_));
  NO4        m0720(.A(mai_mai_n748_), .B(mai_mai_n735_), .C(mai_mai_n729_), .D(mai_mai_n723_), .Y(mai_mai_n749_));
  NA2        m0721(.A(mai_mai_n633_), .B(mai_mai_n393_), .Y(mai_mai_n750_));
  NOi31      m0722(.An(m), .B(h), .C(f), .Y(mai_mai_n751_));
  NA2        m0723(.A(mai_mai_n645_), .B(mai_mai_n751_), .Y(mai_mai_n752_));
  AO210      m0724(.A0(mai_mai_n752_), .A1(mai_mai_n597_), .B0(mai_mai_n545_), .Y(mai_mai_n753_));
  NO3        m0725(.A(mai_mai_n397_), .B(mai_mai_n531_), .C(h), .Y(mai_mai_n754_));
  AOI210     m0726(.A0(mai_mai_n754_), .A1(mai_mai_n114_), .B0(mai_mai_n504_), .Y(mai_mai_n755_));
  NA4        m0727(.A(mai_mai_n755_), .B(mai_mai_n753_), .C(mai_mai_n750_), .D(mai_mai_n257_), .Y(mai_mai_n756_));
  NA2        m0728(.A(mai_mai_n719_), .B(mai_mai_n72_), .Y(mai_mai_n757_));
  NO4        m0729(.A(mai_mai_n696_), .B(mai_mai_n175_), .C(n), .D(i), .Y(mai_mai_n758_));
  NOi21      m0730(.An(h), .B(j), .Y(mai_mai_n759_));
  NA2        m0731(.A(mai_mai_n759_), .B(f), .Y(mai_mai_n760_));
  NO2        m0732(.A(mai_mai_n760_), .B(mai_mai_n251_), .Y(mai_mai_n761_));
  NO3        m0733(.A(mai_mai_n761_), .B(mai_mai_n758_), .C(mai_mai_n699_), .Y(mai_mai_n762_));
  NO2        m0734(.A(mai_mai_n762_), .B(mai_mai_n757_), .Y(mai_mai_n763_));
  AOI210     m0735(.A0(mai_mai_n756_), .A1(l), .B0(mai_mai_n763_), .Y(mai_mai_n764_));
  NO2        m0736(.A(j), .B(i), .Y(mai_mai_n765_));
  NA3        m0737(.A(mai_mai_n765_), .B(mai_mai_n79_), .C(l), .Y(mai_mai_n766_));
  NA2        m0738(.A(mai_mai_n765_), .B(mai_mai_n33_), .Y(mai_mai_n767_));
  OR2        m0739(.A(mai_mai_n766_), .B(mai_mai_n595_), .Y(mai_mai_n768_));
  NO3        m0740(.A(mai_mai_n151_), .B(mai_mai_n49_), .C(mai_mai_n111_), .Y(mai_mai_n769_));
  NO3        m0741(.A(mai_mai_n549_), .B(mai_mai_n149_), .C(mai_mai_n72_), .Y(mai_mai_n770_));
  NO3        m0742(.A(mai_mai_n487_), .B(mai_mai_n437_), .C(j), .Y(mai_mai_n771_));
  OAI210     m0743(.A0(mai_mai_n770_), .A1(mai_mai_n769_), .B0(mai_mai_n771_), .Y(mai_mai_n772_));
  OAI210     m0744(.A0(mai_mai_n752_), .A1(mai_mai_n61_), .B0(mai_mai_n772_), .Y(mai_mai_n773_));
  NA2        m0745(.A(k), .B(j), .Y(mai_mai_n774_));
  NO3        m0746(.A(mai_mai_n299_), .B(mai_mai_n774_), .C(mai_mai_n40_), .Y(mai_mai_n775_));
  AOI210     m0747(.A0(mai_mai_n536_), .A1(n), .B0(mai_mai_n559_), .Y(mai_mai_n776_));
  NA2        m0748(.A(mai_mai_n776_), .B(mai_mai_n562_), .Y(mai_mai_n777_));
  AN3        m0749(.A(mai_mai_n777_), .B(mai_mai_n775_), .C(mai_mai_n98_), .Y(mai_mai_n778_));
  NO3        m0750(.A(mai_mai_n175_), .B(mai_mai_n392_), .C(mai_mai_n113_), .Y(mai_mai_n779_));
  AOI220     m0751(.A0(mai_mai_n779_), .A1(mai_mai_n252_), .B0(mai_mai_n624_), .B1(mai_mai_n308_), .Y(mai_mai_n780_));
  NAi31      m0752(.An(mai_mai_n617_), .B(mai_mai_n92_), .C(mai_mai_n83_), .Y(mai_mai_n781_));
  NA2        m0753(.A(mai_mai_n781_), .B(mai_mai_n780_), .Y(mai_mai_n782_));
  NO2        m0754(.A(mai_mai_n299_), .B(mai_mai_n135_), .Y(mai_mai_n783_));
  AOI220     m0755(.A0(mai_mai_n783_), .A1(mai_mai_n633_), .B0(mai_mai_n732_), .B1(mai_mai_n717_), .Y(mai_mai_n784_));
  NO2        m0756(.A(mai_mai_n741_), .B(mai_mai_n90_), .Y(mai_mai_n785_));
  NA2        m0757(.A(mai_mai_n785_), .B(mai_mai_n594_), .Y(mai_mai_n786_));
  NO2        m0758(.A(mai_mai_n596_), .B(mai_mai_n118_), .Y(mai_mai_n787_));
  OAI210     m0759(.A0(mai_mai_n787_), .A1(mai_mai_n771_), .B0(mai_mai_n684_), .Y(mai_mai_n788_));
  NA3        m0760(.A(mai_mai_n788_), .B(mai_mai_n786_), .C(mai_mai_n784_), .Y(mai_mai_n789_));
  OR4        m0761(.A(mai_mai_n789_), .B(mai_mai_n782_), .C(mai_mai_n778_), .D(mai_mai_n773_), .Y(mai_mai_n790_));
  NA3        m0762(.A(mai_mai_n776_), .B(mai_mai_n562_), .C(mai_mai_n561_), .Y(mai_mai_n791_));
  NA4        m0763(.A(mai_mai_n791_), .B(mai_mai_n219_), .C(mai_mai_n450_), .D(mai_mai_n34_), .Y(mai_mai_n792_));
  NO4        m0764(.A(mai_mai_n487_), .B(mai_mai_n433_), .C(j), .D(f), .Y(mai_mai_n793_));
  OAI220     m0765(.A0(mai_mai_n718_), .A1(mai_mai_n709_), .B0(mai_mai_n333_), .B1(mai_mai_n38_), .Y(mai_mai_n794_));
  AOI210     m0766(.A0(mai_mai_n793_), .A1(mai_mai_n264_), .B0(mai_mai_n794_), .Y(mai_mai_n795_));
  NA3        m0767(.A(mai_mai_n552_), .B(mai_mai_n292_), .C(h), .Y(mai_mai_n796_));
  NOi21      m0768(.An(mai_mai_n684_), .B(mai_mai_n796_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n91_), .B(mai_mai_n47_), .Y(mai_mai_n798_));
  OAI220     m0770(.A0(mai_mai_n796_), .A1(mai_mai_n613_), .B0(mai_mai_n766_), .B1(mai_mai_n677_), .Y(mai_mai_n799_));
  AOI210     m0771(.A0(mai_mai_n798_), .A1(mai_mai_n651_), .B0(mai_mai_n799_), .Y(mai_mai_n800_));
  NAi41      m0772(.An(mai_mai_n797_), .B(mai_mai_n800_), .C(mai_mai_n795_), .D(mai_mai_n792_), .Y(mai_mai_n801_));
  OR2        m0773(.A(mai_mai_n785_), .B(mai_mai_n95_), .Y(mai_mai_n802_));
  AOI220     m0774(.A0(mai_mai_n802_), .A1(mai_mai_n242_), .B0(mai_mai_n771_), .B1(mai_mai_n643_), .Y(mai_mai_n803_));
  NO2        m0775(.A(mai_mai_n669_), .B(mai_mai_n72_), .Y(mai_mai_n804_));
  AOI210     m0776(.A0(mai_mai_n793_), .A1(mai_mai_n804_), .B0(mai_mai_n337_), .Y(mai_mai_n805_));
  OAI210     m0777(.A0(mai_mai_n741_), .A1(mai_mai_n668_), .B0(mai_mai_n524_), .Y(mai_mai_n806_));
  NA3        m0778(.A(mai_mai_n255_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n807_));
  AOI220     m0779(.A0(mai_mai_n612_), .A1(mai_mai_n29_), .B0(mai_mai_n466_), .B1(mai_mai_n83_), .Y(mai_mai_n808_));
  NA2        m0780(.A(mai_mai_n808_), .B(mai_mai_n807_), .Y(mai_mai_n809_));
  NA2        m0781(.A(mai_mai_n809_), .B(mai_mai_n806_), .Y(mai_mai_n810_));
  NA3        m0782(.A(mai_mai_n810_), .B(mai_mai_n805_), .C(mai_mai_n803_), .Y(mai_mai_n811_));
  NOi41      m0783(.An(mai_mai_n768_), .B(mai_mai_n811_), .C(mai_mai_n801_), .D(mai_mai_n790_), .Y(mai_mai_n812_));
  OR3        m0784(.A(mai_mai_n718_), .B(mai_mai_n236_), .C(m), .Y(mai_mai_n813_));
  NO3        m0785(.A(mai_mai_n343_), .B(mai_mai_n301_), .C(mai_mai_n113_), .Y(mai_mai_n814_));
  NA2        m0786(.A(mai_mai_n814_), .B(mai_mai_n777_), .Y(mai_mai_n815_));
  NO3        m0787(.A(mai_mai_n531_), .B(mai_mai_n93_), .C(h), .Y(mai_mai_n816_));
  NA2        m0788(.A(mai_mai_n816_), .B(mai_mai_n713_), .Y(mai_mai_n817_));
  NA4        m0789(.A(mai_mai_n817_), .B(mai_mai_n815_), .C(mai_mai_n813_), .D(mai_mai_n404_), .Y(mai_mai_n818_));
  OR2        m0790(.A(mai_mai_n668_), .B(mai_mai_n91_), .Y(mai_mai_n819_));
  NOi31      m0791(.An(b), .B(d), .C(a), .Y(mai_mai_n820_));
  NO2        m0792(.A(mai_mai_n820_), .B(mai_mai_n610_), .Y(mai_mai_n821_));
  NO2        m0793(.A(mai_mai_n821_), .B(n), .Y(mai_mai_n822_));
  NOi21      m0794(.An(mai_mai_n808_), .B(mai_mai_n822_), .Y(mai_mai_n823_));
  OAI220     m0795(.A0(mai_mai_n823_), .A1(mai_mai_n819_), .B0(mai_mai_n796_), .B1(mai_mai_n611_), .Y(mai_mai_n824_));
  NO2        m0796(.A(mai_mai_n560_), .B(mai_mai_n83_), .Y(mai_mai_n825_));
  NO3        m0797(.A(mai_mai_n632_), .B(mai_mai_n328_), .C(mai_mai_n118_), .Y(mai_mai_n826_));
  NOi21      m0798(.An(mai_mai_n826_), .B(mai_mai_n160_), .Y(mai_mai_n827_));
  AOI210     m0799(.A0(mai_mai_n814_), .A1(mai_mai_n825_), .B0(mai_mai_n827_), .Y(mai_mai_n828_));
  OAI210     m0800(.A0(mai_mai_n718_), .A1(mai_mai_n394_), .B0(mai_mai_n828_), .Y(mai_mai_n829_));
  NO2        m0801(.A(mai_mai_n696_), .B(n), .Y(mai_mai_n830_));
  AOI220     m0802(.A0(mai_mai_n783_), .A1(mai_mai_n673_), .B0(mai_mai_n830_), .B1(mai_mai_n708_), .Y(mai_mai_n831_));
  NO2        m0803(.A(mai_mai_n323_), .B(mai_mai_n241_), .Y(mai_mai_n832_));
  OAI210     m0804(.A0(mai_mai_n95_), .A1(mai_mai_n92_), .B0(mai_mai_n832_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n122_), .B(mai_mai_n83_), .Y(mai_mai_n834_));
  INV        m0806(.A(mai_mai_n833_), .Y(mai_mai_n835_));
  NA2        m0807(.A(mai_mai_n739_), .B(mai_mai_n34_), .Y(mai_mai_n836_));
  NO2        m0808(.A(mai_mai_n278_), .B(i), .Y(mai_mai_n837_));
  OAI210     m0809(.A0(mai_mai_n602_), .A1(mai_mai_n601_), .B0(mai_mai_n365_), .Y(mai_mai_n838_));
  NAi41      m0810(.An(mai_mai_n835_), .B(mai_mai_n838_), .C(mai_mai_n836_), .D(mai_mai_n831_), .Y(mai_mai_n839_));
  NO4        m0811(.A(mai_mai_n839_), .B(mai_mai_n829_), .C(mai_mai_n824_), .D(mai_mai_n818_), .Y(mai_mai_n840_));
  NA4        m0812(.A(mai_mai_n840_), .B(mai_mai_n812_), .C(mai_mai_n764_), .D(mai_mai_n749_), .Y(mai09));
  INV        m0813(.A(mai_mai_n123_), .Y(mai_mai_n842_));
  NA2        m0814(.A(f), .B(e), .Y(mai_mai_n843_));
  NO2        m0815(.A(mai_mai_n229_), .B(mai_mai_n113_), .Y(mai_mai_n844_));
  NA2        m0816(.A(mai_mai_n844_), .B(m), .Y(mai_mai_n845_));
  NA4        m0817(.A(mai_mai_n310_), .B(mai_mai_n165_), .C(mai_mai_n267_), .D(mai_mai_n120_), .Y(mai_mai_n846_));
  AOI210     m0818(.A0(mai_mai_n846_), .A1(m), .B0(mai_mai_n472_), .Y(mai_mai_n847_));
  AOI210     m0819(.A0(mai_mai_n847_), .A1(mai_mai_n845_), .B0(mai_mai_n843_), .Y(mai_mai_n848_));
  NA2        m0820(.A(mai_mai_n443_), .B(e), .Y(mai_mai_n849_));
  NO2        m0821(.A(mai_mai_n849_), .B(mai_mai_n515_), .Y(mai_mai_n850_));
  AOI210     m0822(.A0(mai_mai_n848_), .A1(mai_mai_n842_), .B0(mai_mai_n850_), .Y(mai_mai_n851_));
  NO2        m0823(.A(mai_mai_n207_), .B(mai_mai_n216_), .Y(mai_mai_n852_));
  NA3        m0824(.A(m), .B(l), .C(i), .Y(mai_mai_n853_));
  OAI220     m0825(.A0(mai_mai_n596_), .A1(mai_mai_n853_), .B0(mai_mai_n355_), .B1(mai_mai_n532_), .Y(mai_mai_n854_));
  NAi21      m0826(.An(mai_mai_n854_), .B(mai_mai_n438_), .Y(mai_mai_n855_));
  OR2        m0827(.A(mai_mai_n855_), .B(mai_mai_n852_), .Y(mai_mai_n856_));
  NA3        m0828(.A(mai_mai_n819_), .B(mai_mai_n572_), .C(mai_mai_n524_), .Y(mai_mai_n857_));
  OA210      m0829(.A0(mai_mai_n857_), .A1(mai_mai_n856_), .B0(mai_mai_n822_), .Y(mai_mai_n858_));
  INV        m0830(.A(mai_mai_n340_), .Y(mai_mai_n859_));
  NO2        m0831(.A(mai_mai_n128_), .B(mai_mai_n127_), .Y(mai_mai_n860_));
  NOi31      m0832(.An(k), .B(m), .C(l), .Y(mai_mai_n861_));
  NO2        m0833(.A(mai_mai_n342_), .B(mai_mai_n861_), .Y(mai_mai_n862_));
  AOI210     m0834(.A0(mai_mai_n862_), .A1(mai_mai_n860_), .B0(mai_mai_n605_), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n807_), .B(mai_mai_n333_), .Y(mai_mai_n864_));
  NA2        m0836(.A(mai_mai_n344_), .B(mai_mai_n346_), .Y(mai_mai_n865_));
  OAI210     m0837(.A0(mai_mai_n207_), .A1(mai_mai_n216_), .B0(mai_mai_n865_), .Y(mai_mai_n866_));
  AOI220     m0838(.A0(mai_mai_n866_), .A1(mai_mai_n864_), .B0(mai_mai_n863_), .B1(mai_mai_n859_), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n169_), .B(mai_mai_n115_), .Y(mai_mai_n868_));
  NA3        m0840(.A(mai_mai_n868_), .B(mai_mai_n707_), .C(mai_mai_n135_), .Y(mai_mai_n869_));
  NA3        m0841(.A(mai_mai_n869_), .B(mai_mai_n192_), .C(mai_mai_n31_), .Y(mai_mai_n870_));
  NA4        m0842(.A(mai_mai_n870_), .B(mai_mai_n867_), .C(mai_mai_n634_), .D(mai_mai_n81_), .Y(mai_mai_n871_));
  NO2        m0843(.A(mai_mai_n592_), .B(mai_mai_n500_), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n872_), .B(mai_mai_n192_), .Y(mai_mai_n873_));
  NOi21      m0845(.An(f), .B(d), .Y(mai_mai_n874_));
  NA2        m0846(.A(mai_mai_n874_), .B(m), .Y(mai_mai_n875_));
  NO2        m0847(.A(mai_mai_n875_), .B(mai_mai_n52_), .Y(mai_mai_n876_));
  NOi32      m0848(.An(m), .Bn(f), .C(d), .Y(mai_mai_n877_));
  NA4        m0849(.A(mai_mai_n877_), .B(mai_mai_n612_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n878_));
  NOi21      m0850(.An(mai_mai_n311_), .B(mai_mai_n878_), .Y(mai_mai_n879_));
  AOI210     m0851(.A0(mai_mai_n876_), .A1(mai_mai_n550_), .B0(mai_mai_n879_), .Y(mai_mai_n880_));
  NA3        m0852(.A(mai_mai_n310_), .B(mai_mai_n267_), .C(mai_mai_n120_), .Y(mai_mai_n881_));
  AN2        m0853(.A(f), .B(d), .Y(mai_mai_n882_));
  NA3        m0854(.A(mai_mai_n478_), .B(mai_mai_n882_), .C(mai_mai_n83_), .Y(mai_mai_n883_));
  NO3        m0855(.A(mai_mai_n883_), .B(mai_mai_n72_), .C(mai_mai_n217_), .Y(mai_mai_n884_));
  NA2        m0856(.A(mai_mai_n881_), .B(mai_mai_n884_), .Y(mai_mai_n885_));
  NAi41      m0857(.An(mai_mai_n492_), .B(mai_mai_n885_), .C(mai_mai_n880_), .D(mai_mai_n873_), .Y(mai_mai_n886_));
  NO4        m0858(.A(mai_mai_n632_), .B(mai_mai_n131_), .C(mai_mai_n328_), .D(mai_mai_n152_), .Y(mai_mai_n887_));
  NO2        m0859(.A(mai_mai_n662_), .B(mai_mai_n328_), .Y(mai_mai_n888_));
  AN2        m0860(.A(mai_mai_n888_), .B(mai_mai_n688_), .Y(mai_mai_n889_));
  NO3        m0861(.A(mai_mai_n889_), .B(mai_mai_n887_), .C(mai_mai_n238_), .Y(mai_mai_n890_));
  NA2        m0862(.A(mai_mai_n610_), .B(mai_mai_n83_), .Y(mai_mai_n891_));
  NO2        m0863(.A(mai_mai_n865_), .B(mai_mai_n891_), .Y(mai_mai_n892_));
  NA3        m0864(.A(mai_mai_n159_), .B(mai_mai_n109_), .C(mai_mai_n108_), .Y(mai_mai_n893_));
  OAI220     m0865(.A0(mai_mai_n883_), .A1(mai_mai_n428_), .B0(mai_mai_n340_), .B1(mai_mai_n893_), .Y(mai_mai_n894_));
  NOi41      m0866(.An(mai_mai_n227_), .B(mai_mai_n894_), .C(mai_mai_n892_), .D(mai_mai_n306_), .Y(mai_mai_n895_));
  NA2        m0867(.A(c), .B(mai_mai_n117_), .Y(mai_mai_n896_));
  NO2        m0868(.A(mai_mai_n896_), .B(mai_mai_n408_), .Y(mai_mai_n897_));
  NA3        m0869(.A(mai_mai_n897_), .B(mai_mai_n513_), .C(f), .Y(mai_mai_n898_));
  OR2        m0870(.A(mai_mai_n668_), .B(mai_mai_n546_), .Y(mai_mai_n899_));
  INV        m0871(.A(mai_mai_n899_), .Y(mai_mai_n900_));
  NA2        m0872(.A(mai_mai_n821_), .B(mai_mai_n112_), .Y(mai_mai_n901_));
  NA2        m0873(.A(mai_mai_n901_), .B(mai_mai_n900_), .Y(mai_mai_n902_));
  NA4        m0874(.A(mai_mai_n902_), .B(mai_mai_n898_), .C(mai_mai_n895_), .D(mai_mai_n890_), .Y(mai_mai_n903_));
  NO4        m0875(.A(mai_mai_n903_), .B(mai_mai_n886_), .C(mai_mai_n871_), .D(mai_mai_n858_), .Y(mai_mai_n904_));
  OR2        m0876(.A(mai_mai_n883_), .B(mai_mai_n72_), .Y(mai_mai_n905_));
  NA2        m0877(.A(mai_mai_n844_), .B(m), .Y(mai_mai_n906_));
  AOI210     m0878(.A0(mai_mai_n906_), .A1(mai_mai_n293_), .B0(mai_mai_n905_), .Y(mai_mai_n907_));
  NO2        m0879(.A(mai_mai_n135_), .B(mai_mai_n131_), .Y(mai_mai_n908_));
  NO2        m0880(.A(mai_mai_n234_), .B(mai_mai_n228_), .Y(mai_mai_n909_));
  AOI220     m0881(.A0(mai_mai_n909_), .A1(mai_mai_n231_), .B0(mai_mai_n304_), .B1(mai_mai_n908_), .Y(mai_mai_n910_));
  NO2        m0882(.A(mai_mai_n428_), .B(mai_mai_n843_), .Y(mai_mai_n911_));
  INV        m0883(.A(mai_mai_n910_), .Y(mai_mai_n912_));
  NA2        m0884(.A(e), .B(d), .Y(mai_mai_n913_));
  OAI220     m0885(.A0(mai_mai_n913_), .A1(c), .B0(mai_mai_n323_), .B1(d), .Y(mai_mai_n914_));
  NA3        m0886(.A(mai_mai_n914_), .B(mai_mai_n455_), .C(mai_mai_n511_), .Y(mai_mai_n915_));
  AOI210     m0887(.A0(mai_mai_n519_), .A1(mai_mai_n182_), .B0(mai_mai_n234_), .Y(mai_mai_n916_));
  AOI210     m0888(.A0(mai_mai_n633_), .A1(mai_mai_n349_), .B0(mai_mai_n916_), .Y(mai_mai_n917_));
  INV        m0889(.A(mai_mai_n165_), .Y(mai_mai_n918_));
  NA2        m0890(.A(mai_mai_n884_), .B(mai_mai_n918_), .Y(mai_mai_n919_));
  NA3        m0891(.A(mai_mai_n168_), .B(mai_mai_n84_), .C(mai_mai_n34_), .Y(mai_mai_n920_));
  NA4        m0892(.A(mai_mai_n920_), .B(mai_mai_n919_), .C(mai_mai_n917_), .D(mai_mai_n915_), .Y(mai_mai_n921_));
  NO3        m0893(.A(mai_mai_n921_), .B(mai_mai_n912_), .C(mai_mai_n907_), .Y(mai_mai_n922_));
  NA2        m0894(.A(mai_mai_n859_), .B(mai_mai_n31_), .Y(mai_mai_n923_));
  AO210      m0895(.A0(mai_mai_n923_), .A1(mai_mai_n709_), .B0(mai_mai_n220_), .Y(mai_mai_n924_));
  OAI220     m0896(.A0(mai_mai_n632_), .A1(mai_mai_n60_), .B0(mai_mai_n301_), .B1(j), .Y(mai_mai_n925_));
  AOI220     m0897(.A0(mai_mai_n925_), .A1(mai_mai_n888_), .B0(mai_mai_n622_), .B1(mai_mai_n631_), .Y(mai_mai_n926_));
  OAI210     m0898(.A0(mai_mai_n849_), .A1(mai_mai_n172_), .B0(mai_mai_n926_), .Y(mai_mai_n927_));
  OAI210     m0899(.A0(mai_mai_n844_), .A1(mai_mai_n918_), .B0(mai_mai_n877_), .Y(mai_mai_n928_));
  NO2        m0900(.A(mai_mai_n928_), .B(mai_mai_n613_), .Y(mai_mai_n929_));
  AOI210     m0901(.A0(mai_mai_n119_), .A1(mai_mai_n118_), .B0(mai_mai_n266_), .Y(mai_mai_n930_));
  NO2        m0902(.A(mai_mai_n930_), .B(mai_mai_n878_), .Y(mai_mai_n931_));
  AO210      m0903(.A0(mai_mai_n864_), .A1(mai_mai_n854_), .B0(mai_mai_n931_), .Y(mai_mai_n932_));
  NO3        m0904(.A(mai_mai_n932_), .B(mai_mai_n929_), .C(mai_mai_n927_), .Y(mai_mai_n933_));
  AO220      m0905(.A0(mai_mai_n455_), .A1(mai_mai_n759_), .B0(mai_mai_n177_), .B1(f), .Y(mai_mai_n934_));
  OAI210     m0906(.A0(mai_mai_n934_), .A1(mai_mai_n458_), .B0(mai_mai_n914_), .Y(mai_mai_n935_));
  NA2        m0907(.A(mai_mai_n857_), .B(mai_mai_n713_), .Y(mai_mai_n936_));
  AN4        m0908(.A(mai_mai_n936_), .B(mai_mai_n935_), .C(mai_mai_n933_), .D(mai_mai_n924_), .Y(mai_mai_n937_));
  NA4        m0909(.A(mai_mai_n937_), .B(mai_mai_n922_), .C(mai_mai_n904_), .D(mai_mai_n851_), .Y(mai12));
  NO2        m0910(.A(mai_mai_n453_), .B(c), .Y(mai_mai_n939_));
  NO4        m0911(.A(mai_mai_n442_), .B(mai_mai_n258_), .C(mai_mai_n588_), .D(mai_mai_n217_), .Y(mai_mai_n940_));
  NA2        m0912(.A(mai_mai_n940_), .B(mai_mai_n939_), .Y(mai_mai_n941_));
  NO2        m0913(.A(mai_mai_n453_), .B(mai_mai_n117_), .Y(mai_mai_n942_));
  NO2        m0914(.A(mai_mai_n860_), .B(mai_mai_n355_), .Y(mai_mai_n943_));
  NO2        m0915(.A(mai_mai_n668_), .B(mai_mai_n378_), .Y(mai_mai_n944_));
  AOI220     m0916(.A0(mai_mai_n944_), .A1(mai_mai_n548_), .B0(mai_mai_n943_), .B1(mai_mai_n942_), .Y(mai_mai_n945_));
  NA3        m0917(.A(mai_mai_n945_), .B(mai_mai_n941_), .C(mai_mai_n441_), .Y(mai_mai_n946_));
  AOI210     m0918(.A0(mai_mai_n237_), .A1(mai_mai_n339_), .B0(mai_mai_n204_), .Y(mai_mai_n947_));
  OR2        m0919(.A(mai_mai_n947_), .B(mai_mai_n940_), .Y(mai_mai_n948_));
  AOI210     m0920(.A0(mai_mai_n336_), .A1(mai_mai_n390_), .B0(mai_mai_n217_), .Y(mai_mai_n949_));
  OAI210     m0921(.A0(mai_mai_n949_), .A1(mai_mai_n948_), .B0(mai_mai_n403_), .Y(mai_mai_n950_));
  NO2        m0922(.A(mai_mai_n648_), .B(mai_mai_n269_), .Y(mai_mai_n951_));
  NO2        m0923(.A(mai_mai_n596_), .B(mai_mai_n853_), .Y(mai_mai_n952_));
  AOI220     m0924(.A0(mai_mai_n952_), .A1(mai_mai_n570_), .B0(mai_mai_n832_), .B1(mai_mai_n951_), .Y(mai_mai_n953_));
  NO2        m0925(.A(mai_mai_n151_), .B(mai_mai_n241_), .Y(mai_mai_n954_));
  NA2        m0926(.A(mai_mai_n953_), .B(mai_mai_n950_), .Y(mai_mai_n955_));
  OR2        m0927(.A(mai_mai_n324_), .B(mai_mai_n942_), .Y(mai_mai_n956_));
  NA2        m0928(.A(mai_mai_n956_), .B(mai_mai_n356_), .Y(mai_mai_n957_));
  NO3        m0929(.A(mai_mai_n131_), .B(mai_mai_n152_), .C(mai_mai_n217_), .Y(mai_mai_n958_));
  NA2        m0930(.A(mai_mai_n958_), .B(mai_mai_n536_), .Y(mai_mai_n959_));
  NA4        m0931(.A(mai_mai_n443_), .B(mai_mai_n435_), .C(mai_mai_n183_), .D(m), .Y(mai_mai_n960_));
  NA3        m0932(.A(mai_mai_n960_), .B(mai_mai_n959_), .C(mai_mai_n957_), .Y(mai_mai_n961_));
  NO3        m0933(.A(mai_mai_n671_), .B(mai_mai_n91_), .C(mai_mai_n45_), .Y(mai_mai_n962_));
  NO4        m0934(.A(mai_mai_n962_), .B(mai_mai_n961_), .C(mai_mai_n955_), .D(mai_mai_n946_), .Y(mai_mai_n963_));
  NO2        m0935(.A(mai_mai_n371_), .B(mai_mai_n370_), .Y(mai_mai_n964_));
  NA2        m0936(.A(mai_mai_n593_), .B(mai_mai_n70_), .Y(mai_mai_n965_));
  NA2        m0937(.A(mai_mai_n560_), .B(mai_mai_n144_), .Y(mai_mai_n966_));
  NOi21      m0938(.An(mai_mai_n34_), .B(mai_mai_n662_), .Y(mai_mai_n967_));
  AOI220     m0939(.A0(mai_mai_n967_), .A1(mai_mai_n966_), .B0(mai_mai_n965_), .B1(mai_mai_n964_), .Y(mai_mai_n968_));
  OAI210     m0940(.A0(mai_mai_n256_), .A1(mai_mai_n45_), .B0(mai_mai_n968_), .Y(mai_mai_n969_));
  NO3        m0941(.A(mai_mai_n834_), .B(mai_mai_n88_), .C(mai_mai_n408_), .Y(mai_mai_n970_));
  NAi21      m0942(.An(mai_mai_n970_), .B(mai_mai_n320_), .Y(mai_mai_n971_));
  NO2        m0943(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n972_));
  NO2        m0944(.A(mai_mai_n507_), .B(mai_mai_n301_), .Y(mai_mai_n973_));
  INV        m0945(.A(mai_mai_n973_), .Y(mai_mai_n974_));
  NO2        m0946(.A(mai_mai_n974_), .B(mai_mai_n144_), .Y(mai_mai_n975_));
  NA2        m0947(.A(mai_mai_n641_), .B(mai_mai_n365_), .Y(mai_mai_n976_));
  OAI210     m0948(.A0(mai_mai_n745_), .A1(mai_mai_n976_), .B0(mai_mai_n369_), .Y(mai_mai_n977_));
  NO4        m0949(.A(mai_mai_n977_), .B(mai_mai_n975_), .C(mai_mai_n971_), .D(mai_mai_n969_), .Y(mai_mai_n978_));
  NA2        m0950(.A(mai_mai_n349_), .B(m), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n162_), .B(i), .Y(mai_mai_n980_));
  NA2        m0952(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n981_));
  OAI220     m0953(.A0(mai_mai_n981_), .A1(mai_mai_n203_), .B0(mai_mai_n980_), .B1(mai_mai_n91_), .Y(mai_mai_n982_));
  AOI210     m0954(.A0(mai_mai_n419_), .A1(mai_mai_n37_), .B0(mai_mai_n982_), .Y(mai_mai_n983_));
  NO2        m0955(.A(mai_mai_n144_), .B(mai_mai_n83_), .Y(mai_mai_n984_));
  OR2        m0956(.A(mai_mai_n984_), .B(mai_mai_n559_), .Y(mai_mai_n985_));
  NA2        m0957(.A(mai_mai_n560_), .B(mai_mai_n382_), .Y(mai_mai_n986_));
  AOI210     m0958(.A0(mai_mai_n986_), .A1(n), .B0(mai_mai_n985_), .Y(mai_mai_n987_));
  OAI220     m0959(.A0(mai_mai_n987_), .A1(mai_mai_n979_), .B0(mai_mai_n983_), .B1(mai_mai_n333_), .Y(mai_mai_n988_));
  NO2        m0960(.A(mai_mai_n668_), .B(mai_mai_n500_), .Y(mai_mai_n989_));
  NA3        m0961(.A(mai_mai_n344_), .B(mai_mai_n636_), .C(i), .Y(mai_mai_n990_));
  OAI210     m0962(.A0(mai_mai_n437_), .A1(mai_mai_n310_), .B0(mai_mai_n990_), .Y(mai_mai_n991_));
  OAI220     m0963(.A0(mai_mai_n991_), .A1(mai_mai_n989_), .B0(mai_mai_n684_), .B1(mai_mai_n770_), .Y(mai_mai_n992_));
  NA2        m0964(.A(mai_mai_n616_), .B(mai_mai_n114_), .Y(mai_mai_n993_));
  OR3        m0965(.A(mai_mai_n310_), .B(mai_mai_n433_), .C(f), .Y(mai_mai_n994_));
  NA3        m0966(.A(mai_mai_n636_), .B(mai_mai_n79_), .C(i), .Y(mai_mai_n995_));
  OA220      m0967(.A0(mai_mai_n995_), .A1(mai_mai_n993_), .B0(mai_mai_n994_), .B1(mai_mai_n595_), .Y(mai_mai_n996_));
  NA3        m0968(.A(mai_mai_n325_), .B(mai_mai_n119_), .C(m), .Y(mai_mai_n997_));
  AOI210     m0969(.A0(mai_mai_n681_), .A1(mai_mai_n997_), .B0(m), .Y(mai_mai_n998_));
  OAI210     m0970(.A0(mai_mai_n998_), .A1(mai_mai_n943_), .B0(mai_mai_n324_), .Y(mai_mai_n999_));
  NA2        m0971(.A(mai_mai_n700_), .B(mai_mai_n891_), .Y(mai_mai_n1000_));
  INV        m0972(.A(mai_mai_n438_), .Y(mai_mai_n1001_));
  NA2        m0973(.A(mai_mai_n225_), .B(mai_mai_n76_), .Y(mai_mai_n1002_));
  NA3        m0974(.A(mai_mai_n1002_), .B(mai_mai_n995_), .C(mai_mai_n994_), .Y(mai_mai_n1003_));
  AOI220     m0975(.A0(mai_mai_n1003_), .A1(mai_mai_n264_), .B0(mai_mai_n1001_), .B1(mai_mai_n1000_), .Y(mai_mai_n1004_));
  NA4        m0976(.A(mai_mai_n1004_), .B(mai_mai_n999_), .C(mai_mai_n996_), .D(mai_mai_n992_), .Y(mai_mai_n1005_));
  NO2        m0977(.A(mai_mai_n378_), .B(mai_mai_n90_), .Y(mai_mai_n1006_));
  OAI210     m0978(.A0(mai_mai_n1006_), .A1(mai_mai_n951_), .B0(mai_mai_n242_), .Y(mai_mai_n1007_));
  NA2        m0979(.A(mai_mai_n670_), .B(mai_mai_n87_), .Y(mai_mai_n1008_));
  NO2        m0980(.A(mai_mai_n461_), .B(mai_mai_n217_), .Y(mai_mai_n1009_));
  AOI220     m0981(.A0(mai_mai_n1009_), .A1(mai_mai_n383_), .B0(mai_mai_n956_), .B1(mai_mai_n221_), .Y(mai_mai_n1010_));
  AOI220     m0982(.A0(mai_mai_n944_), .A1(mai_mai_n954_), .B0(mai_mai_n594_), .B1(mai_mai_n89_), .Y(mai_mai_n1011_));
  NA4        m0983(.A(mai_mai_n1011_), .B(mai_mai_n1010_), .C(mai_mai_n1008_), .D(mai_mai_n1007_), .Y(mai_mai_n1012_));
  OAI210     m0984(.A0(mai_mai_n1001_), .A1(mai_mai_n952_), .B0(mai_mai_n548_), .Y(mai_mai_n1013_));
  AOI210     m0985(.A0(mai_mai_n420_), .A1(mai_mai_n412_), .B0(mai_mai_n834_), .Y(mai_mai_n1014_));
  OAI210     m0986(.A0(mai_mai_n371_), .A1(mai_mai_n370_), .B0(mai_mai_n110_), .Y(mai_mai_n1015_));
  AOI210     m0987(.A0(mai_mai_n1015_), .A1(mai_mai_n540_), .B0(mai_mai_n1014_), .Y(mai_mai_n1016_));
  NA2        m0988(.A(mai_mai_n998_), .B(mai_mai_n942_), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n653_), .B(mai_mai_n536_), .Y(mai_mai_n1018_));
  NA4        m0990(.A(mai_mai_n1018_), .B(mai_mai_n1017_), .C(mai_mai_n1016_), .D(mai_mai_n1013_), .Y(mai_mai_n1019_));
  NO4        m0991(.A(mai_mai_n1019_), .B(mai_mai_n1012_), .C(mai_mai_n1005_), .D(mai_mai_n988_), .Y(mai_mai_n1020_));
  NAi31      m0992(.An(mai_mai_n140_), .B(mai_mai_n421_), .C(n), .Y(mai_mai_n1021_));
  NO3        m0993(.A(mai_mai_n127_), .B(mai_mai_n342_), .C(mai_mai_n861_), .Y(mai_mai_n1022_));
  NO2        m0994(.A(mai_mai_n1022_), .B(mai_mai_n1021_), .Y(mai_mai_n1023_));
  NO3        m0995(.A(mai_mai_n278_), .B(mai_mai_n140_), .C(mai_mai_n408_), .Y(mai_mai_n1024_));
  AOI210     m0996(.A0(mai_mai_n1024_), .A1(mai_mai_n501_), .B0(mai_mai_n1023_), .Y(mai_mai_n1025_));
  NA2        m0997(.A(mai_mai_n493_), .B(i), .Y(mai_mai_n1026_));
  NA2        m0998(.A(mai_mai_n1026_), .B(mai_mai_n1025_), .Y(mai_mai_n1027_));
  NA2        m0999(.A(mai_mai_n234_), .B(mai_mai_n173_), .Y(mai_mai_n1028_));
  NO3        m1000(.A(mai_mai_n308_), .B(mai_mai_n443_), .C(mai_mai_n177_), .Y(mai_mai_n1029_));
  NOi31      m1001(.An(mai_mai_n1028_), .B(mai_mai_n1029_), .C(mai_mai_n217_), .Y(mai_mai_n1030_));
  NAi21      m1002(.An(mai_mai_n560_), .B(mai_mai_n1009_), .Y(mai_mai_n1031_));
  NA2        m1003(.A(mai_mai_n436_), .B(mai_mai_n891_), .Y(mai_mai_n1032_));
  NO3        m1004(.A(mai_mai_n437_), .B(mai_mai_n310_), .C(mai_mai_n72_), .Y(mai_mai_n1033_));
  AOI220     m1005(.A0(mai_mai_n1033_), .A1(mai_mai_n1032_), .B0(mai_mai_n484_), .B1(m), .Y(mai_mai_n1034_));
  NA2        m1006(.A(mai_mai_n1034_), .B(mai_mai_n1031_), .Y(mai_mai_n1035_));
  OAI220     m1007(.A0(mai_mai_n1021_), .A1(mai_mai_n237_), .B0(mai_mai_n990_), .B1(mai_mai_n611_), .Y(mai_mai_n1036_));
  NA2        m1008(.A(mai_mai_n947_), .B(mai_mai_n939_), .Y(mai_mai_n1037_));
  NO3        m1009(.A(mai_mai_n549_), .B(mai_mai_n149_), .C(mai_mai_n216_), .Y(mai_mai_n1038_));
  OAI210     m1010(.A0(mai_mai_n1038_), .A1(mai_mai_n530_), .B0(mai_mai_n379_), .Y(mai_mai_n1039_));
  OAI220     m1011(.A0(mai_mai_n944_), .A1(mai_mai_n952_), .B0(mai_mai_n550_), .B1(mai_mai_n427_), .Y(mai_mai_n1040_));
  NA4        m1012(.A(mai_mai_n1040_), .B(mai_mai_n1039_), .C(mai_mai_n1037_), .D(mai_mai_n630_), .Y(mai_mai_n1041_));
  OAI210     m1013(.A0(mai_mai_n947_), .A1(mai_mai_n940_), .B0(mai_mai_n1028_), .Y(mai_mai_n1042_));
  NA3        m1014(.A(mai_mai_n986_), .B(mai_mai_n489_), .C(mai_mai_n46_), .Y(mai_mai_n1043_));
  AOI210     m1015(.A0(mai_mai_n381_), .A1(mai_mai_n379_), .B0(mai_mai_n332_), .Y(mai_mai_n1044_));
  NA3        m1016(.A(mai_mai_n1044_), .B(mai_mai_n1043_), .C(mai_mai_n1042_), .Y(mai_mai_n1045_));
  OR3        m1017(.A(mai_mai_n1045_), .B(mai_mai_n1041_), .C(mai_mai_n1036_), .Y(mai_mai_n1046_));
  NO4        m1018(.A(mai_mai_n1046_), .B(mai_mai_n1035_), .C(mai_mai_n1030_), .D(mai_mai_n1027_), .Y(mai_mai_n1047_));
  NA4        m1019(.A(mai_mai_n1047_), .B(mai_mai_n1020_), .C(mai_mai_n978_), .D(mai_mai_n963_), .Y(mai13));
  AN2        m1020(.A(c), .B(b), .Y(mai_mai_n1049_));
  NA3        m1021(.A(mai_mai_n255_), .B(mai_mai_n1049_), .C(m), .Y(mai_mai_n1050_));
  NA2        m1022(.A(mai_mai_n498_), .B(f), .Y(mai_mai_n1051_));
  NO4        m1023(.A(mai_mai_n1051_), .B(mai_mai_n1050_), .C(mai_mai_n1547_), .D(mai_mai_n589_), .Y(mai_mai_n1052_));
  NA2        m1024(.A(mai_mai_n271_), .B(mai_mai_n1049_), .Y(mai_mai_n1053_));
  NO4        m1025(.A(mai_mai_n1053_), .B(mai_mai_n1051_), .C(mai_mai_n980_), .D(a), .Y(mai_mai_n1054_));
  NAi32      m1026(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1055_));
  NA2        m1027(.A(mai_mai_n139_), .B(mai_mai_n45_), .Y(mai_mai_n1056_));
  NO4        m1028(.A(mai_mai_n1056_), .B(mai_mai_n1055_), .C(mai_mai_n596_), .D(mai_mai_n307_), .Y(mai_mai_n1057_));
  NA2        m1029(.A(mai_mai_n674_), .B(mai_mai_n228_), .Y(mai_mai_n1058_));
  NA2        m1030(.A(mai_mai_n411_), .B(mai_mai_n216_), .Y(mai_mai_n1059_));
  AN2        m1031(.A(d), .B(c), .Y(mai_mai_n1060_));
  NA2        m1032(.A(mai_mai_n1060_), .B(mai_mai_n117_), .Y(mai_mai_n1061_));
  NO4        m1033(.A(mai_mai_n1061_), .B(mai_mai_n1059_), .C(mai_mai_n178_), .D(mai_mai_n169_), .Y(mai_mai_n1062_));
  NA2        m1034(.A(mai_mai_n498_), .B(c), .Y(mai_mai_n1063_));
  NO4        m1035(.A(mai_mai_n1056_), .B(mai_mai_n592_), .C(mai_mai_n1063_), .D(mai_mai_n307_), .Y(mai_mai_n1064_));
  AO210      m1036(.A0(mai_mai_n1062_), .A1(mai_mai_n1058_), .B0(mai_mai_n1064_), .Y(mai_mai_n1065_));
  OR4        m1037(.A(mai_mai_n1065_), .B(mai_mai_n1057_), .C(mai_mai_n1054_), .D(mai_mai_n1052_), .Y(mai_mai_n1066_));
  NAi32      m1038(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1067_));
  NO2        m1039(.A(mai_mai_n1067_), .B(mai_mai_n146_), .Y(mai_mai_n1068_));
  NA2        m1040(.A(mai_mai_n1068_), .B(m), .Y(mai_mai_n1069_));
  OR3        m1041(.A(mai_mai_n228_), .B(mai_mai_n178_), .C(mai_mai_n169_), .Y(mai_mai_n1070_));
  NO2        m1042(.A(mai_mai_n1070_), .B(mai_mai_n1069_), .Y(mai_mai_n1071_));
  NO2        m1043(.A(mai_mai_n1063_), .B(mai_mai_n307_), .Y(mai_mai_n1072_));
  NO2        m1044(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1073_));
  NA2        m1045(.A(mai_mai_n638_), .B(mai_mai_n1073_), .Y(mai_mai_n1074_));
  NOi21      m1046(.An(mai_mai_n1072_), .B(mai_mai_n1074_), .Y(mai_mai_n1075_));
  NO2        m1047(.A(mai_mai_n774_), .B(mai_mai_n113_), .Y(mai_mai_n1076_));
  NOi41      m1048(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1077_));
  NA2        m1049(.A(mai_mai_n1077_), .B(mai_mai_n1076_), .Y(mai_mai_n1078_));
  NO2        m1050(.A(mai_mai_n1078_), .B(mai_mai_n1069_), .Y(mai_mai_n1079_));
  OR3        m1051(.A(e), .B(d), .C(c), .Y(mai_mai_n1080_));
  NA3        m1052(.A(k), .B(j), .C(i), .Y(mai_mai_n1081_));
  NO3        m1053(.A(mai_mai_n1081_), .B(mai_mai_n307_), .C(mai_mai_n90_), .Y(mai_mai_n1082_));
  NOi21      m1054(.An(mai_mai_n1082_), .B(mai_mai_n1080_), .Y(mai_mai_n1083_));
  OR4        m1055(.A(mai_mai_n1083_), .B(mai_mai_n1079_), .C(mai_mai_n1075_), .D(mai_mai_n1071_), .Y(mai_mai_n1084_));
  NO2        m1056(.A(f), .B(c), .Y(mai_mai_n1085_));
  NOi21      m1057(.An(mai_mai_n1085_), .B(mai_mai_n442_), .Y(mai_mai_n1086_));
  NA2        m1058(.A(mai_mai_n1086_), .B(mai_mai_n59_), .Y(mai_mai_n1087_));
  OR2        m1059(.A(k), .B(i), .Y(mai_mai_n1088_));
  NO3        m1060(.A(mai_mai_n1088_), .B(mai_mai_n248_), .C(l), .Y(mai_mai_n1089_));
  NOi31      m1061(.An(mai_mai_n1089_), .B(mai_mai_n1087_), .C(j), .Y(mai_mai_n1090_));
  OR3        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1084_), .C(mai_mai_n1066_), .Y(mai02));
  OR2        m1063(.A(l), .B(k), .Y(mai_mai_n1092_));
  OR3        m1064(.A(h), .B(m), .C(f), .Y(mai_mai_n1093_));
  OR3        m1065(.A(n), .B(m), .C(i), .Y(mai_mai_n1094_));
  NO4        m1066(.A(mai_mai_n1094_), .B(mai_mai_n1093_), .C(mai_mai_n1092_), .D(mai_mai_n1080_), .Y(mai_mai_n1095_));
  NOi31      m1067(.An(e), .B(d), .C(c), .Y(mai_mai_n1096_));
  AOI210     m1068(.A0(mai_mai_n1082_), .A1(mai_mai_n1096_), .B0(mai_mai_n1057_), .Y(mai_mai_n1097_));
  AN3        m1069(.A(m), .B(f), .C(c), .Y(mai_mai_n1098_));
  INV        m1070(.A(mai_mai_n1071_), .Y(mai_mai_n1099_));
  NA3        m1071(.A(l), .B(k), .C(j), .Y(mai_mai_n1100_));
  NA2        m1072(.A(i), .B(h), .Y(mai_mai_n1101_));
  NO3        m1073(.A(mai_mai_n1101_), .B(mai_mai_n1100_), .C(mai_mai_n131_), .Y(mai_mai_n1102_));
  NO3        m1074(.A(mai_mai_n141_), .B(mai_mai_n289_), .C(mai_mai_n217_), .Y(mai_mai_n1103_));
  INV        m1075(.A(mai_mai_n1075_), .Y(mai_mai_n1104_));
  NA3        m1076(.A(c), .B(b), .C(a), .Y(mai_mai_n1105_));
  NO3        m1077(.A(mai_mai_n1105_), .B(mai_mai_n913_), .C(mai_mai_n216_), .Y(mai_mai_n1106_));
  NO3        m1078(.A(mai_mai_n1081_), .B(mai_mai_n49_), .C(mai_mai_n113_), .Y(mai_mai_n1107_));
  NA2        m1079(.A(mai_mai_n1107_), .B(mai_mai_n1106_), .Y(mai_mai_n1108_));
  AN3        m1080(.A(mai_mai_n1108_), .B(mai_mai_n1104_), .C(mai_mai_n1099_), .Y(mai_mai_n1109_));
  NO2        m1081(.A(mai_mai_n1061_), .B(mai_mai_n1059_), .Y(mai_mai_n1110_));
  NA2        m1082(.A(mai_mai_n1078_), .B(mai_mai_n1070_), .Y(mai_mai_n1111_));
  AOI210     m1083(.A0(mai_mai_n1111_), .A1(mai_mai_n1110_), .B0(mai_mai_n1052_), .Y(mai_mai_n1112_));
  NAi41      m1084(.An(mai_mai_n1095_), .B(mai_mai_n1112_), .C(mai_mai_n1109_), .D(mai_mai_n1097_), .Y(mai03));
  NO2        m1085(.A(mai_mai_n532_), .B(mai_mai_n605_), .Y(mai_mai_n1114_));
  NA4        m1086(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(m), .D(mai_mai_n216_), .Y(mai_mai_n1115_));
  NA4        m1087(.A(mai_mai_n580_), .B(m), .C(mai_mai_n113_), .D(mai_mai_n216_), .Y(mai_mai_n1116_));
  NA3        m1088(.A(mai_mai_n1116_), .B(mai_mai_n372_), .C(mai_mai_n1115_), .Y(mai_mai_n1117_));
  NO3        m1089(.A(mai_mai_n1117_), .B(mai_mai_n1114_), .C(mai_mai_n1015_), .Y(mai_mai_n1118_));
  NOi41      m1090(.An(mai_mai_n819_), .B(mai_mai_n866_), .C(mai_mai_n855_), .D(mai_mai_n727_), .Y(mai_mai_n1119_));
  OAI220     m1091(.A0(mai_mai_n1119_), .A1(mai_mai_n700_), .B0(mai_mai_n1118_), .B1(mai_mai_n593_), .Y(mai_mai_n1120_));
  NOi31      m1092(.An(m), .B(n), .C(f), .Y(mai_mai_n1121_));
  NA2        m1093(.A(mai_mai_n1121_), .B(mai_mai_n51_), .Y(mai_mai_n1122_));
  AN2        m1094(.A(e), .B(c), .Y(mai_mai_n1123_));
  NA2        m1095(.A(mai_mai_n1123_), .B(a), .Y(mai_mai_n1124_));
  OAI220     m1096(.A0(mai_mai_n1124_), .A1(mai_mai_n1122_), .B0(mai_mai_n899_), .B1(mai_mai_n426_), .Y(mai_mai_n1125_));
  NA2        m1097(.A(mai_mai_n511_), .B(l), .Y(mai_mai_n1126_));
  NOi31      m1098(.An(mai_mai_n877_), .B(mai_mai_n1050_), .C(mai_mai_n1126_), .Y(mai_mai_n1127_));
  NO3        m1099(.A(mai_mai_n1127_), .B(mai_mai_n1125_), .C(mai_mai_n1014_), .Y(mai_mai_n1128_));
  NO2        m1100(.A(mai_mai_n289_), .B(a), .Y(mai_mai_n1129_));
  INV        m1101(.A(mai_mai_n1057_), .Y(mai_mai_n1130_));
  NO2        m1102(.A(mai_mai_n1101_), .B(mai_mai_n487_), .Y(mai_mai_n1131_));
  NO2        m1103(.A(mai_mai_n86_), .B(m), .Y(mai_mai_n1132_));
  AOI210     m1104(.A0(mai_mai_n1132_), .A1(mai_mai_n1131_), .B0(mai_mai_n1089_), .Y(mai_mai_n1133_));
  OR2        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1087_), .Y(mai_mai_n1134_));
  NA3        m1106(.A(mai_mai_n1134_), .B(mai_mai_n1130_), .C(mai_mai_n1128_), .Y(mai_mai_n1135_));
  NO4        m1107(.A(mai_mai_n1135_), .B(mai_mai_n1120_), .C(mai_mai_n835_), .D(mai_mai_n569_), .Y(mai_mai_n1136_));
  NA2        m1108(.A(c), .B(b), .Y(mai_mai_n1137_));
  NO2        m1109(.A(mai_mai_n712_), .B(mai_mai_n1137_), .Y(mai_mai_n1138_));
  OAI210     m1110(.A0(mai_mai_n875_), .A1(mai_mai_n847_), .B0(mai_mai_n415_), .Y(mai_mai_n1139_));
  OAI210     m1111(.A0(mai_mai_n1139_), .A1(mai_mai_n876_), .B0(mai_mai_n1138_), .Y(mai_mai_n1140_));
  NAi21      m1112(.An(mai_mai_n423_), .B(mai_mai_n1138_), .Y(mai_mai_n1141_));
  OAI210     m1113(.A0(mai_mai_n554_), .A1(mai_mai_n39_), .B0(mai_mai_n1129_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n1142_), .B(mai_mai_n1141_), .Y(mai_mai_n1143_));
  NA2        m1115(.A(mai_mai_n267_), .B(mai_mai_n120_), .Y(mai_mai_n1144_));
  NA2        m1116(.A(mai_mai_n1144_), .B(m), .Y(mai_mai_n1145_));
  NAi21      m1117(.An(f), .B(d), .Y(mai_mai_n1146_));
  NO2        m1118(.A(mai_mai_n1146_), .B(mai_mai_n1105_), .Y(mai_mai_n1147_));
  INV        m1119(.A(mai_mai_n1147_), .Y(mai_mai_n1148_));
  AOI210     m1120(.A0(mai_mai_n1145_), .A1(mai_mai_n293_), .B0(mai_mai_n1148_), .Y(mai_mai_n1149_));
  AOI210     m1121(.A0(mai_mai_n1149_), .A1(mai_mai_n114_), .B0(mai_mai_n1143_), .Y(mai_mai_n1150_));
  NO2        m1122(.A(mai_mai_n184_), .B(mai_mai_n241_), .Y(mai_mai_n1151_));
  NA2        m1123(.A(mai_mai_n1151_), .B(m), .Y(mai_mai_n1152_));
  NA3        m1124(.A(mai_mai_n930_), .B(mai_mai_n1126_), .C(mai_mai_n165_), .Y(mai_mai_n1153_));
  OAI210     m1125(.A0(mai_mai_n1153_), .A1(mai_mai_n311_), .B0(mai_mai_n473_), .Y(mai_mai_n1154_));
  NO2        m1126(.A(mai_mai_n1154_), .B(mai_mai_n1152_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n158_), .B(mai_mai_n33_), .Y(mai_mai_n1156_));
  AOI210     m1128(.A0(mai_mai_n976_), .A1(mai_mai_n1156_), .B0(mai_mai_n217_), .Y(mai_mai_n1157_));
  OAI210     m1129(.A0(mai_mai_n1157_), .A1(mai_mai_n446_), .B0(mai_mai_n1147_), .Y(mai_mai_n1158_));
  AOI210     m1130(.A0(mai_mai_n1151_), .A1(mai_mai_n429_), .B0(mai_mai_n970_), .Y(mai_mai_n1159_));
  NA2        m1131(.A(mai_mai_n1159_), .B(mai_mai_n1158_), .Y(mai_mai_n1160_));
  NO2        m1132(.A(mai_mai_n1160_), .B(mai_mai_n1155_), .Y(mai_mai_n1161_));
  NA4        m1133(.A(mai_mai_n1161_), .B(mai_mai_n1150_), .C(mai_mai_n1140_), .D(mai_mai_n1136_), .Y(mai00));
  AOI210     m1134(.A0(mai_mai_n300_), .A1(mai_mai_n217_), .B0(mai_mai_n281_), .Y(mai_mai_n1163_));
  NO2        m1135(.A(mai_mai_n1163_), .B(mai_mai_n583_), .Y(mai_mai_n1164_));
  NA2        m1136(.A(mai_mai_n911_), .B(mai_mai_n954_), .Y(mai_mai_n1165_));
  NO2        m1137(.A(mai_mai_n970_), .B(mai_mai_n724_), .Y(mai_mai_n1166_));
  NA3        m1138(.A(mai_mai_n1166_), .B(mai_mai_n1165_), .C(mai_mai_n1016_), .Y(mai_mai_n1167_));
  NA2        m1139(.A(mai_mai_n513_), .B(f), .Y(mai_mai_n1168_));
  OAI210     m1140(.A0(mai_mai_n1022_), .A1(mai_mai_n40_), .B0(mai_mai_n655_), .Y(mai_mai_n1169_));
  NA3        m1141(.A(mai_mai_n1169_), .B(mai_mai_n263_), .C(n), .Y(mai_mai_n1170_));
  AOI210     m1142(.A0(mai_mai_n1170_), .A1(mai_mai_n1168_), .B0(mai_mai_n1061_), .Y(mai_mai_n1171_));
  NO4        m1143(.A(mai_mai_n1171_), .B(mai_mai_n1167_), .C(mai_mai_n1164_), .D(mai_mai_n1084_), .Y(mai_mai_n1172_));
  NA3        m1144(.A(mai_mai_n168_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1173_));
  NA3        m1145(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1174_));
  NOi31      m1146(.An(n), .B(m), .C(i), .Y(mai_mai_n1175_));
  NA3        m1147(.A(mai_mai_n1175_), .B(mai_mai_n658_), .C(mai_mai_n51_), .Y(mai_mai_n1176_));
  OAI210     m1148(.A0(mai_mai_n1174_), .A1(mai_mai_n1173_), .B0(mai_mai_n1176_), .Y(mai_mai_n1177_));
  INV        m1149(.A(mai_mai_n582_), .Y(mai_mai_n1178_));
  NO2        m1150(.A(mai_mai_n1178_), .B(mai_mai_n1177_), .Y(mai_mai_n1179_));
  NO4        m1151(.A(mai_mai_n490_), .B(mai_mai_n358_), .C(mai_mai_n1137_), .D(mai_mai_n59_), .Y(mai_mai_n1180_));
  NA3        m1152(.A(mai_mai_n384_), .B(mai_mai_n224_), .C(m), .Y(mai_mai_n1181_));
  OR2        m1153(.A(mai_mai_n1181_), .B(mai_mai_n1174_), .Y(mai_mai_n1182_));
  NO2        m1154(.A(h), .B(m), .Y(mai_mai_n1183_));
  NA4        m1155(.A(mai_mai_n501_), .B(mai_mai_n469_), .C(mai_mai_n1183_), .D(mai_mai_n1049_), .Y(mai_mai_n1184_));
  OAI220     m1156(.A0(mai_mai_n532_), .A1(mai_mai_n605_), .B0(mai_mai_n91_), .B1(mai_mai_n90_), .Y(mai_mai_n1185_));
  AOI220     m1157(.A0(mai_mai_n1185_), .A1(mai_mai_n540_), .B0(mai_mai_n958_), .B1(mai_mai_n581_), .Y(mai_mai_n1186_));
  AOI220     m1158(.A0(mai_mai_n317_), .A1(mai_mai_n252_), .B0(mai_mai_n179_), .B1(mai_mai_n148_), .Y(mai_mai_n1187_));
  NA4        m1159(.A(mai_mai_n1187_), .B(mai_mai_n1186_), .C(mai_mai_n1184_), .D(mai_mai_n1182_), .Y(mai_mai_n1188_));
  NO3        m1160(.A(mai_mai_n1188_), .B(mai_mai_n1180_), .C(mai_mai_n273_), .Y(mai_mai_n1189_));
  INV        m1161(.A(mai_mai_n322_), .Y(mai_mai_n1190_));
  AOI210     m1162(.A0(mai_mai_n252_), .A1(mai_mai_n349_), .B0(mai_mai_n584_), .Y(mai_mai_n1191_));
  NA2        m1163(.A(mai_mai_n1191_), .B(mai_mai_n1190_), .Y(mai_mai_n1192_));
  NO2        m1164(.A(mai_mai_n243_), .B(mai_mai_n183_), .Y(mai_mai_n1193_));
  NA2        m1165(.A(mai_mai_n1193_), .B(mai_mai_n427_), .Y(mai_mai_n1194_));
  NAi31      m1166(.An(mai_mai_n188_), .B(mai_mai_n872_), .C(mai_mai_n469_), .Y(mai_mai_n1195_));
  NA2        m1167(.A(mai_mai_n1195_), .B(mai_mai_n1194_), .Y(mai_mai_n1196_));
  NO2        m1168(.A(mai_mai_n280_), .B(mai_mai_n72_), .Y(mai_mai_n1197_));
  NO3        m1169(.A(mai_mai_n426_), .B(mai_mai_n843_), .C(n), .Y(mai_mai_n1198_));
  AOI210     m1170(.A0(mai_mai_n1198_), .A1(mai_mai_n1197_), .B0(mai_mai_n1095_), .Y(mai_mai_n1199_));
  NAi31      m1171(.An(mai_mai_n1064_), .B(mai_mai_n1199_), .C(mai_mai_n71_), .Y(mai_mai_n1200_));
  NO4        m1172(.A(mai_mai_n1200_), .B(mai_mai_n1196_), .C(mai_mai_n1192_), .D(mai_mai_n523_), .Y(mai_mai_n1201_));
  AN3        m1173(.A(mai_mai_n1201_), .B(mai_mai_n1189_), .C(mai_mai_n1179_), .Y(mai_mai_n1202_));
  NA2        m1174(.A(mai_mai_n540_), .B(mai_mai_n101_), .Y(mai_mai_n1203_));
  NA3        m1175(.A(mai_mai_n1121_), .B(mai_mai_n616_), .C(mai_mai_n468_), .Y(mai_mai_n1204_));
  NA3        m1176(.A(mai_mai_n1204_), .B(mai_mai_n1203_), .C(mai_mai_n246_), .Y(mai_mai_n1205_));
  NA2        m1177(.A(mai_mai_n1117_), .B(mai_mai_n540_), .Y(mai_mai_n1206_));
  NA4        m1178(.A(mai_mai_n658_), .B(mai_mai_n209_), .C(mai_mai_n224_), .D(mai_mai_n162_), .Y(mai_mai_n1207_));
  NA3        m1179(.A(mai_mai_n1207_), .B(mai_mai_n1206_), .C(mai_mai_n297_), .Y(mai_mai_n1208_));
  OAI210     m1180(.A0(mai_mai_n467_), .A1(mai_mai_n121_), .B0(mai_mai_n878_), .Y(mai_mai_n1209_));
  NA2        m1181(.A(mai_mai_n1209_), .B(mai_mai_n1153_), .Y(mai_mai_n1210_));
  OR4        m1182(.A(mai_mai_n1061_), .B(mai_mai_n278_), .C(mai_mai_n226_), .D(e), .Y(mai_mai_n1211_));
  NO2        m1183(.A(mai_mai_n220_), .B(mai_mai_n217_), .Y(mai_mai_n1212_));
  NA2        m1184(.A(n), .B(e), .Y(mai_mai_n1213_));
  NO2        m1185(.A(mai_mai_n1213_), .B(mai_mai_n146_), .Y(mai_mai_n1214_));
  AOI220     m1186(.A0(mai_mai_n1214_), .A1(mai_mai_n279_), .B0(mai_mai_n859_), .B1(mai_mai_n1212_), .Y(mai_mai_n1215_));
  OAI210     m1187(.A0(mai_mai_n359_), .A1(mai_mai_n312_), .B0(mai_mai_n448_), .Y(mai_mai_n1216_));
  NA4        m1188(.A(mai_mai_n1216_), .B(mai_mai_n1215_), .C(mai_mai_n1211_), .D(mai_mai_n1210_), .Y(mai_mai_n1217_));
  NA2        m1189(.A(mai_mai_n1214_), .B(mai_mai_n863_), .Y(mai_mai_n1218_));
  AOI220     m1190(.A0(mai_mai_n967_), .A1(mai_mai_n581_), .B0(mai_mai_n658_), .B1(mai_mai_n249_), .Y(mai_mai_n1219_));
  NO2        m1191(.A(mai_mai_n65_), .B(h), .Y(mai_mai_n1220_));
  NO3        m1192(.A(mai_mai_n1061_), .B(mai_mai_n1059_), .C(mai_mai_n738_), .Y(mai_mai_n1221_));
  NO2        m1193(.A(mai_mai_n1092_), .B(mai_mai_n131_), .Y(mai_mai_n1222_));
  AN2        m1194(.A(mai_mai_n1222_), .B(mai_mai_n1103_), .Y(mai_mai_n1223_));
  OAI210     m1195(.A0(mai_mai_n1223_), .A1(mai_mai_n1221_), .B0(mai_mai_n1220_), .Y(mai_mai_n1224_));
  NA4        m1196(.A(mai_mai_n1224_), .B(mai_mai_n1219_), .C(mai_mai_n1218_), .D(mai_mai_n880_), .Y(mai_mai_n1225_));
  NO4        m1197(.A(mai_mai_n1225_), .B(mai_mai_n1217_), .C(mai_mai_n1208_), .D(mai_mai_n1205_), .Y(mai_mai_n1226_));
  NA2        m1198(.A(mai_mai_n848_), .B(mai_mai_n769_), .Y(mai_mai_n1227_));
  NA4        m1199(.A(mai_mai_n1227_), .B(mai_mai_n1226_), .C(mai_mai_n1202_), .D(mai_mai_n1172_), .Y(mai01));
  AN2        m1200(.A(mai_mai_n1039_), .B(mai_mai_n1037_), .Y(mai_mai_n1229_));
  NO2        m1201(.A(mai_mai_n481_), .B(mai_mai_n287_), .Y(mai_mai_n1230_));
  NA2        m1202(.A(mai_mai_n395_), .B(i), .Y(mai_mai_n1231_));
  NA3        m1203(.A(mai_mai_n1231_), .B(mai_mai_n1230_), .C(mai_mai_n1229_), .Y(mai_mai_n1232_));
  NA2        m1204(.A(mai_mai_n594_), .B(mai_mai_n89_), .Y(mai_mai_n1233_));
  NA2        m1205(.A(mai_mai_n560_), .B(mai_mai_n277_), .Y(mai_mai_n1234_));
  NA2        m1206(.A(mai_mai_n973_), .B(mai_mai_n1234_), .Y(mai_mai_n1235_));
  NA4        m1207(.A(mai_mai_n1235_), .B(mai_mai_n1233_), .C(mai_mai_n926_), .D(mai_mai_n334_), .Y(mai_mai_n1236_));
  NA2        m1208(.A(mai_mai_n45_), .B(f), .Y(mai_mai_n1237_));
  NA2        m1209(.A(mai_mai_n719_), .B(mai_mai_n96_), .Y(mai_mai_n1238_));
  NO2        m1210(.A(mai_mai_n1238_), .B(mai_mai_n1237_), .Y(mai_mai_n1239_));
  OAI210     m1211(.A0(mai_mai_n796_), .A1(mai_mai_n611_), .B0(mai_mai_n1207_), .Y(mai_mai_n1240_));
  INV        m1212(.A(mai_mai_n1240_), .Y(mai_mai_n1241_));
  INV        m1213(.A(mai_mai_n119_), .Y(mai_mai_n1242_));
  OA220      m1214(.A0(mai_mai_n1242_), .A1(mai_mai_n591_), .B0(mai_mai_n669_), .B1(mai_mai_n372_), .Y(mai_mai_n1243_));
  NAi41      m1215(.An(mai_mai_n161_), .B(mai_mai_n1243_), .C(mai_mai_n1241_), .D(mai_mai_n910_), .Y(mai_mai_n1244_));
  NO3        m1216(.A(mai_mai_n797_), .B(mai_mai_n683_), .C(mai_mai_n516_), .Y(mai_mai_n1245_));
  NA4        m1217(.A(mai_mai_n719_), .B(mai_mai_n96_), .C(mai_mai_n45_), .D(mai_mai_n216_), .Y(mai_mai_n1246_));
  OA220      m1218(.A0(mai_mai_n1246_), .A1(mai_mai_n677_), .B0(mai_mai_n198_), .B1(mai_mai_n196_), .Y(mai_mai_n1247_));
  NA3        m1219(.A(mai_mai_n1247_), .B(mai_mai_n1245_), .C(mai_mai_n136_), .Y(mai_mai_n1248_));
  NO4        m1220(.A(mai_mai_n1248_), .B(mai_mai_n1244_), .C(mai_mai_n1236_), .D(mai_mai_n1232_), .Y(mai_mai_n1249_));
  INV        m1221(.A(mai_mai_n1181_), .Y(mai_mai_n1250_));
  NA2        m1222(.A(mai_mai_n1250_), .B(mai_mai_n536_), .Y(mai_mai_n1251_));
  NA2        m1223(.A(mai_mai_n543_), .B(mai_mai_n397_), .Y(mai_mai_n1252_));
  NOi21      m1224(.An(mai_mai_n566_), .B(mai_mai_n588_), .Y(mai_mai_n1253_));
  NA2        m1225(.A(mai_mai_n1253_), .B(mai_mai_n1252_), .Y(mai_mai_n1254_));
  AOI210     m1226(.A0(mai_mai_n207_), .A1(mai_mai_n88_), .B0(mai_mai_n216_), .Y(mai_mai_n1255_));
  OAI210     m1227(.A0(mai_mai_n822_), .A1(mai_mai_n427_), .B0(mai_mai_n1255_), .Y(mai_mai_n1256_));
  AN3        m1228(.A(m), .B(l), .C(k), .Y(mai_mai_n1257_));
  OAI210     m1229(.A0(mai_mai_n361_), .A1(mai_mai_n34_), .B0(mai_mai_n1257_), .Y(mai_mai_n1258_));
  NA2        m1230(.A(mai_mai_n206_), .B(mai_mai_n34_), .Y(mai_mai_n1259_));
  AO210      m1231(.A0(mai_mai_n1259_), .A1(mai_mai_n1258_), .B0(mai_mai_n333_), .Y(mai_mai_n1260_));
  NA4        m1232(.A(mai_mai_n1260_), .B(mai_mai_n1256_), .C(mai_mai_n1254_), .D(mai_mai_n1251_), .Y(mai_mai_n1261_));
  AOI210     m1233(.A0(mai_mai_n603_), .A1(mai_mai_n119_), .B0(mai_mai_n609_), .Y(mai_mai_n1262_));
  OAI210     m1234(.A0(mai_mai_n1242_), .A1(mai_mai_n600_), .B0(mai_mai_n1262_), .Y(mai_mai_n1263_));
  NA2        m1235(.A(mai_mai_n286_), .B(mai_mai_n198_), .Y(mai_mai_n1264_));
  NA2        m1236(.A(mai_mai_n1264_), .B(mai_mai_n673_), .Y(mai_mai_n1265_));
  INV        m1237(.A(mai_mai_n970_), .Y(mai_mai_n1266_));
  OAI210     m1238(.A0(mai_mai_n1239_), .A1(mai_mai_n327_), .B0(mai_mai_n684_), .Y(mai_mai_n1267_));
  NA4        m1239(.A(mai_mai_n1267_), .B(mai_mai_n1266_), .C(mai_mai_n1265_), .D(mai_mai_n800_), .Y(mai_mai_n1268_));
  NO3        m1240(.A(mai_mai_n1268_), .B(mai_mai_n1263_), .C(mai_mai_n1261_), .Y(mai_mai_n1269_));
  NA3        m1241(.A(mai_mai_n612_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1270_));
  NO2        m1242(.A(mai_mai_n1270_), .B(mai_mai_n207_), .Y(mai_mai_n1271_));
  AOI210     m1243(.A0(mai_mai_n508_), .A1(mai_mai_n58_), .B0(mai_mai_n1271_), .Y(mai_mai_n1272_));
  OR3        m1244(.A(mai_mai_n1238_), .B(mai_mai_n613_), .C(mai_mai_n1237_), .Y(mai_mai_n1273_));
  NO2        m1245(.A(mai_mai_n1246_), .B(mai_mai_n993_), .Y(mai_mai_n1274_));
  NO2        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1177_), .Y(mai_mai_n1275_));
  NA4        m1247(.A(mai_mai_n1275_), .B(mai_mai_n1273_), .C(mai_mai_n1272_), .D(mai_mai_n768_), .Y(mai_mai_n1276_));
  NO2        m1248(.A(mai_mai_n980_), .B(mai_mai_n236_), .Y(mai_mai_n1277_));
  NO2        m1249(.A(mai_mai_n981_), .B(mai_mai_n562_), .Y(mai_mai_n1278_));
  OAI210     m1250(.A0(mai_mai_n1278_), .A1(mai_mai_n1277_), .B0(mai_mai_n342_), .Y(mai_mai_n1279_));
  NA2        m1251(.A(mai_mai_n576_), .B(mai_mai_n574_), .Y(mai_mai_n1280_));
  NO3        m1252(.A(mai_mai_n78_), .B(mai_mai_n301_), .C(mai_mai_n45_), .Y(mai_mai_n1281_));
  NA2        m1253(.A(mai_mai_n1281_), .B(mai_mai_n559_), .Y(mai_mai_n1282_));
  NA3        m1254(.A(mai_mai_n1282_), .B(mai_mai_n1280_), .C(mai_mai_n679_), .Y(mai_mai_n1283_));
  OR2        m1255(.A(mai_mai_n1181_), .B(mai_mai_n1174_), .Y(mai_mai_n1284_));
  NO2        m1256(.A(mai_mai_n372_), .B(mai_mai_n70_), .Y(mai_mai_n1285_));
  INV        m1257(.A(mai_mai_n1285_), .Y(mai_mai_n1286_));
  NA2        m1258(.A(mai_mai_n1281_), .B(mai_mai_n825_), .Y(mai_mai_n1287_));
  NA4        m1259(.A(mai_mai_n1287_), .B(mai_mai_n1286_), .C(mai_mai_n1284_), .D(mai_mai_n387_), .Y(mai_mai_n1288_));
  NOi41      m1260(.An(mai_mai_n1279_), .B(mai_mai_n1288_), .C(mai_mai_n1283_), .D(mai_mai_n1276_), .Y(mai_mai_n1289_));
  NO2        m1261(.A(mai_mai_n130_), .B(mai_mai_n45_), .Y(mai_mai_n1290_));
  NO2        m1262(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1291_));
  AO220      m1263(.A0(mai_mai_n1291_), .A1(mai_mai_n633_), .B0(mai_mai_n1290_), .B1(mai_mai_n717_), .Y(mai_mai_n1292_));
  NA2        m1264(.A(mai_mai_n1292_), .B(mai_mai_n342_), .Y(mai_mai_n1293_));
  INV        m1265(.A(mai_mai_n134_), .Y(mai_mai_n1294_));
  NO3        m1266(.A(mai_mai_n1101_), .B(mai_mai_n178_), .C(mai_mai_n86_), .Y(mai_mai_n1295_));
  AOI220     m1267(.A0(mai_mai_n1295_), .A1(mai_mai_n1294_), .B0(mai_mai_n1281_), .B1(mai_mai_n984_), .Y(mai_mai_n1296_));
  NA2        m1268(.A(mai_mai_n1296_), .B(mai_mai_n1293_), .Y(mai_mai_n1297_));
  NO2        m1269(.A(mai_mai_n624_), .B(mai_mai_n623_), .Y(mai_mai_n1298_));
  NO4        m1270(.A(mai_mai_n1101_), .B(mai_mai_n1298_), .C(mai_mai_n176_), .D(mai_mai_n86_), .Y(mai_mai_n1299_));
  NO3        m1271(.A(mai_mai_n1299_), .B(mai_mai_n1297_), .C(mai_mai_n647_), .Y(mai_mai_n1300_));
  NA4        m1272(.A(mai_mai_n1300_), .B(mai_mai_n1289_), .C(mai_mai_n1269_), .D(mai_mai_n1249_), .Y(mai06));
  NO2        m1273(.A(mai_mai_n228_), .B(mai_mai_n103_), .Y(mai_mai_n1302_));
  OAI210     m1274(.A0(mai_mai_n1302_), .A1(mai_mai_n1295_), .B0(mai_mai_n383_), .Y(mai_mai_n1303_));
  NO3        m1275(.A(mai_mai_n607_), .B(mai_mai_n820_), .C(mai_mai_n610_), .Y(mai_mai_n1304_));
  OR2        m1276(.A(mai_mai_n1304_), .B(mai_mai_n899_), .Y(mai_mai_n1305_));
  NA3        m1277(.A(mai_mai_n1305_), .B(mai_mai_n1303_), .C(mai_mai_n1279_), .Y(mai_mai_n1306_));
  NO3        m1278(.A(mai_mai_n1306_), .B(mai_mai_n1283_), .C(mai_mai_n262_), .Y(mai_mai_n1307_));
  NO2        m1279(.A(mai_mai_n301_), .B(mai_mai_n45_), .Y(mai_mai_n1308_));
  AOI210     m1280(.A0(mai_mai_n1308_), .A1(mai_mai_n985_), .B0(mai_mai_n1277_), .Y(mai_mai_n1309_));
  AOI210     m1281(.A0(mai_mai_n1308_), .A1(mai_mai_n563_), .B0(mai_mai_n1292_), .Y(mai_mai_n1310_));
  AOI210     m1282(.A0(mai_mai_n1310_), .A1(mai_mai_n1309_), .B0(mai_mai_n339_), .Y(mai_mai_n1311_));
  INV        m1283(.A(mai_mai_n682_), .Y(mai_mai_n1312_));
  NA2        m1284(.A(mai_mai_n1312_), .B(mai_mai_n651_), .Y(mai_mai_n1313_));
  NO2        m1285(.A(mai_mai_n519_), .B(mai_mai_n173_), .Y(mai_mai_n1314_));
  NO2        m1286(.A(mai_mai_n617_), .B(mai_mai_n1122_), .Y(mai_mai_n1315_));
  OAI210     m1287(.A0(mai_mai_n462_), .A1(mai_mai_n253_), .B0(mai_mai_n920_), .Y(mai_mai_n1316_));
  NO3        m1288(.A(mai_mai_n1316_), .B(mai_mai_n1315_), .C(mai_mai_n1314_), .Y(mai_mai_n1317_));
  OR2        m1289(.A(mai_mai_n608_), .B(mai_mai_n606_), .Y(mai_mai_n1318_));
  NO2        m1290(.A(mai_mai_n371_), .B(mai_mai_n135_), .Y(mai_mai_n1319_));
  AOI210     m1291(.A0(mai_mai_n1319_), .A1(mai_mai_n594_), .B0(mai_mai_n1318_), .Y(mai_mai_n1320_));
  NA3        m1292(.A(mai_mai_n1320_), .B(mai_mai_n1317_), .C(mai_mai_n1313_), .Y(mai_mai_n1321_));
  NO2        m1293(.A(mai_mai_n760_), .B(mai_mai_n370_), .Y(mai_mai_n1322_));
  NO3        m1294(.A(mai_mai_n684_), .B(mai_mai_n770_), .C(mai_mai_n643_), .Y(mai_mai_n1323_));
  NOi21      m1295(.An(mai_mai_n1322_), .B(mai_mai_n1323_), .Y(mai_mai_n1324_));
  AN2        m1296(.A(mai_mai_n967_), .B(mai_mai_n654_), .Y(mai_mai_n1325_));
  NO4        m1297(.A(mai_mai_n1325_), .B(mai_mai_n1324_), .C(mai_mai_n1321_), .D(mai_mai_n1311_), .Y(mai_mai_n1326_));
  OAI220     m1298(.A0(mai_mai_n744_), .A1(mai_mai_n47_), .B0(mai_mai_n228_), .B1(mai_mai_n626_), .Y(mai_mai_n1327_));
  NA2        m1299(.A(mai_mai_n364_), .B(mai_mai_n1327_), .Y(mai_mai_n1328_));
  NO3        m1300(.A(mai_mai_n248_), .B(mai_mai_n103_), .C(mai_mai_n289_), .Y(mai_mai_n1329_));
  OAI220     m1301(.A0(mai_mai_n709_), .A1(mai_mai_n253_), .B0(mai_mai_n515_), .B1(mai_mai_n519_), .Y(mai_mai_n1330_));
  OAI210     m1302(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1331_));
  NO3        m1303(.A(mai_mai_n1331_), .B(mai_mai_n605_), .C(j), .Y(mai_mai_n1332_));
  NOi21      m1304(.An(mai_mai_n1332_), .B(mai_mai_n677_), .Y(mai_mai_n1333_));
  NO4        m1305(.A(mai_mai_n1333_), .B(mai_mai_n1330_), .C(mai_mai_n1329_), .D(mai_mai_n1125_), .Y(mai_mai_n1334_));
  NA4        m1306(.A(mai_mai_n808_), .B(mai_mai_n807_), .C(mai_mai_n436_), .D(mai_mai_n891_), .Y(mai_mai_n1335_));
  NAi31      m1307(.An(mai_mai_n760_), .B(mai_mai_n1335_), .C(mai_mai_n206_), .Y(mai_mai_n1336_));
  NA4        m1308(.A(mai_mai_n1336_), .B(mai_mai_n1334_), .C(mai_mai_n1328_), .D(mai_mai_n1219_), .Y(mai_mai_n1337_));
  NOi21      m1309(.An(mai_mai_n1304_), .B(mai_mai_n466_), .Y(mai_mai_n1338_));
  OR3        m1310(.A(mai_mai_n1338_), .B(mai_mai_n796_), .C(mai_mai_n546_), .Y(mai_mai_n1339_));
  NA2        m1311(.A(mai_mai_n576_), .B(mai_mai_n448_), .Y(mai_mai_n1340_));
  NA2        m1312(.A(mai_mai_n1332_), .B(mai_mai_n804_), .Y(mai_mai_n1341_));
  NA3        m1313(.A(mai_mai_n1341_), .B(mai_mai_n1340_), .C(mai_mai_n1339_), .Y(mai_mai_n1342_));
  AOI220     m1314(.A0(mai_mai_n1322_), .A1(mai_mai_n769_), .B0(mai_mai_n1319_), .B1(mai_mai_n242_), .Y(mai_mai_n1343_));
  AN2        m1315(.A(mai_mai_n940_), .B(mai_mai_n939_), .Y(mai_mai_n1344_));
  NO4        m1316(.A(mai_mai_n1344_), .B(mai_mai_n889_), .C(mai_mai_n504_), .D(mai_mai_n484_), .Y(mai_mai_n1345_));
  NA3        m1317(.A(mai_mai_n1345_), .B(mai_mai_n1343_), .C(mai_mai_n1287_), .Y(mai_mai_n1346_));
  NAi21      m1318(.An(j), .B(i), .Y(mai_mai_n1347_));
  NO4        m1319(.A(mai_mai_n1298_), .B(mai_mai_n1347_), .C(mai_mai_n442_), .D(mai_mai_n239_), .Y(mai_mai_n1348_));
  NO4        m1320(.A(mai_mai_n1348_), .B(mai_mai_n1346_), .C(mai_mai_n1342_), .D(mai_mai_n1337_), .Y(mai_mai_n1349_));
  NA4        m1321(.A(mai_mai_n1349_), .B(mai_mai_n1326_), .C(mai_mai_n1307_), .D(mai_mai_n1300_), .Y(mai07));
  NAi32      m1322(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1351_));
  NO3        m1323(.A(mai_mai_n1351_), .B(m), .C(f), .Y(mai_mai_n1352_));
  OAI210     m1324(.A0(mai_mai_n321_), .A1(mai_mai_n486_), .B0(mai_mai_n1352_), .Y(mai_mai_n1353_));
  NAi21      m1325(.An(f), .B(c), .Y(mai_mai_n1354_));
  OR2        m1326(.A(e), .B(d), .Y(mai_mai_n1355_));
  OAI220     m1327(.A0(mai_mai_n1355_), .A1(mai_mai_n1354_), .B0(mai_mai_n637_), .B1(mai_mai_n323_), .Y(mai_mai_n1356_));
  NA3        m1328(.A(mai_mai_n1356_), .B(mai_mai_n1073_), .C(mai_mai_n181_), .Y(mai_mai_n1357_));
  NOi31      m1329(.An(n), .B(m), .C(b), .Y(mai_mai_n1358_));
  NO3        m1330(.A(mai_mai_n131_), .B(mai_mai_n450_), .C(h), .Y(mai_mai_n1359_));
  NA2        m1331(.A(mai_mai_n1357_), .B(mai_mai_n1353_), .Y(mai_mai_n1360_));
  NOi41      m1332(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1361_));
  INV        m1333(.A(k), .Y(mai_mai_n1362_));
  NA2        m1334(.A(mai_mai_n1103_), .B(mai_mai_n224_), .Y(mai_mai_n1363_));
  NO2        m1335(.A(mai_mai_n1363_), .B(mai_mai_n60_), .Y(mai_mai_n1364_));
  NO2        m1336(.A(k), .B(i), .Y(mai_mai_n1365_));
  NA3        m1337(.A(mai_mai_n1365_), .B(mai_mai_n909_), .C(mai_mai_n181_), .Y(mai_mai_n1366_));
  NA2        m1338(.A(mai_mai_n86_), .B(mai_mai_n45_), .Y(mai_mai_n1367_));
  NO2        m1339(.A(mai_mai_n1067_), .B(mai_mai_n442_), .Y(mai_mai_n1368_));
  NA3        m1340(.A(mai_mai_n1368_), .B(mai_mai_n1367_), .C(mai_mai_n217_), .Y(mai_mai_n1369_));
  NO2        m1341(.A(mai_mai_n1081_), .B(mai_mai_n307_), .Y(mai_mai_n1370_));
  NA2        m1342(.A(mai_mai_n547_), .B(mai_mai_n79_), .Y(mai_mai_n1371_));
  NA2        m1343(.A(mai_mai_n1220_), .B(mai_mai_n291_), .Y(mai_mai_n1372_));
  NA4        m1344(.A(mai_mai_n1372_), .B(mai_mai_n1371_), .C(mai_mai_n1369_), .D(mai_mai_n1366_), .Y(mai_mai_n1373_));
  NO3        m1345(.A(mai_mai_n1373_), .B(mai_mai_n1364_), .C(mai_mai_n1360_), .Y(mai_mai_n1374_));
  NO3        m1346(.A(e), .B(d), .C(c), .Y(mai_mai_n1375_));
  OAI210     m1347(.A0(mai_mai_n131_), .A1(mai_mai_n217_), .B0(mai_mai_n614_), .Y(mai_mai_n1376_));
  NA2        m1348(.A(mai_mai_n1376_), .B(mai_mai_n1375_), .Y(mai_mai_n1377_));
  NO2        m1349(.A(mai_mai_n1377_), .B(c), .Y(mai_mai_n1378_));
  OR2        m1350(.A(h), .B(f), .Y(mai_mai_n1379_));
  NO3        m1351(.A(n), .B(m), .C(i), .Y(mai_mai_n1380_));
  OAI210     m1352(.A0(mai_mai_n1123_), .A1(mai_mai_n156_), .B0(mai_mai_n1380_), .Y(mai_mai_n1381_));
  NO2        m1353(.A(mai_mai_n1381_), .B(mai_mai_n1379_), .Y(mai_mai_n1382_));
  NA3        m1354(.A(mai_mai_n706_), .B(mai_mai_n692_), .C(mai_mai_n113_), .Y(mai_mai_n1383_));
  NO2        m1355(.A(mai_mai_n1383_), .B(mai_mai_n45_), .Y(mai_mai_n1384_));
  NO2        m1356(.A(l), .B(k), .Y(mai_mai_n1385_));
  NOi31      m1357(.An(mai_mai_n552_), .B(mai_mai_n479_), .C(mai_mai_n442_), .Y(mai_mai_n1386_));
  NO3        m1358(.A(mai_mai_n442_), .B(d), .C(c), .Y(mai_mai_n1387_));
  NO4        m1359(.A(mai_mai_n1386_), .B(mai_mai_n1384_), .C(mai_mai_n1382_), .D(mai_mai_n1378_), .Y(mai_mai_n1388_));
  NO2        m1360(.A(mai_mai_n147_), .B(h), .Y(mai_mai_n1389_));
  NO2        m1361(.A(mai_mai_n1088_), .B(l), .Y(mai_mai_n1390_));
  NO2        m1362(.A(m), .B(c), .Y(mai_mai_n1391_));
  NA3        m1363(.A(mai_mai_n1391_), .B(mai_mai_n141_), .C(mai_mai_n189_), .Y(mai_mai_n1392_));
  NO2        m1364(.A(mai_mai_n1392_), .B(mai_mai_n1390_), .Y(mai_mai_n1393_));
  NA2        m1365(.A(mai_mai_n1393_), .B(mai_mai_n181_), .Y(mai_mai_n1394_));
  NA2        m1366(.A(mai_mai_n1362_), .B(mai_mai_n1088_), .Y(mai_mai_n1395_));
  NO2        m1367(.A(mai_mai_n453_), .B(a), .Y(mai_mai_n1396_));
  NA3        m1368(.A(mai_mai_n1396_), .B(mai_mai_n1395_), .C(mai_mai_n114_), .Y(mai_mai_n1397_));
  NO2        m1369(.A(i), .B(h), .Y(mai_mai_n1398_));
  NA2        m1370(.A(mai_mai_n1146_), .B(h), .Y(mai_mai_n1399_));
  NA2        m1371(.A(mai_mai_n137_), .B(mai_mai_n224_), .Y(mai_mai_n1400_));
  NO2        m1372(.A(mai_mai_n1400_), .B(mai_mai_n1399_), .Y(mai_mai_n1401_));
  NO2        m1373(.A(mai_mai_n767_), .B(mai_mai_n190_), .Y(mai_mai_n1402_));
  NOi31      m1374(.An(m), .B(n), .C(b), .Y(mai_mai_n1403_));
  NOi31      m1375(.An(f), .B(d), .C(c), .Y(mai_mai_n1404_));
  NA2        m1376(.A(mai_mai_n1404_), .B(mai_mai_n1403_), .Y(mai_mai_n1405_));
  INV        m1377(.A(mai_mai_n1405_), .Y(mai_mai_n1406_));
  NO3        m1378(.A(mai_mai_n1406_), .B(mai_mai_n1402_), .C(mai_mai_n1401_), .Y(mai_mai_n1407_));
  NA2        m1379(.A(mai_mai_n1098_), .B(mai_mai_n469_), .Y(mai_mai_n1408_));
  NO3        m1380(.A(mai_mai_n1408_), .B(mai_mai_n442_), .C(mai_mai_n45_), .Y(mai_mai_n1409_));
  OAI210     m1381(.A0(mai_mai_n184_), .A1(mai_mai_n531_), .B0(mai_mai_n1077_), .Y(mai_mai_n1410_));
  NO3        m1382(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1411_));
  INV        m1383(.A(mai_mai_n1410_), .Y(mai_mai_n1412_));
  NO2        m1384(.A(mai_mai_n1412_), .B(mai_mai_n1409_), .Y(mai_mai_n1413_));
  AN4        m1385(.A(mai_mai_n1413_), .B(mai_mai_n1407_), .C(mai_mai_n1397_), .D(mai_mai_n1394_), .Y(mai_mai_n1414_));
  NA2        m1386(.A(mai_mai_n1358_), .B(mai_mai_n380_), .Y(mai_mai_n1415_));
  NO2        m1387(.A(mai_mai_n1415_), .B(mai_mai_n1058_), .Y(mai_mai_n1416_));
  NA2        m1388(.A(mai_mai_n1387_), .B(mai_mai_n218_), .Y(mai_mai_n1417_));
  NO2        m1389(.A(mai_mai_n190_), .B(b), .Y(mai_mai_n1418_));
  AOI210     m1390(.A0(mai_mai_n1175_), .A1(mai_mai_n1418_), .B0(mai_mai_n1102_), .Y(mai_mai_n1419_));
  NAi31      m1391(.An(mai_mai_n1416_), .B(mai_mai_n1419_), .C(mai_mai_n1417_), .Y(mai_mai_n1420_));
  NO4        m1392(.A(mai_mai_n131_), .B(m), .C(f), .D(e), .Y(mai_mai_n1421_));
  NA3        m1393(.A(mai_mai_n1365_), .B(mai_mai_n292_), .C(h), .Y(mai_mai_n1422_));
  OR2        m1394(.A(e), .B(a), .Y(mai_mai_n1423_));
  NO2        m1395(.A(mai_mai_n1355_), .B(mai_mai_n1354_), .Y(mai_mai_n1424_));
  AOI210     m1396(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1424_), .Y(mai_mai_n1425_));
  NO2        m1397(.A(mai_mai_n1425_), .B(mai_mai_n1094_), .Y(mai_mai_n1426_));
  NA2        m1398(.A(mai_mai_n1361_), .B(mai_mai_n1385_), .Y(mai_mai_n1427_));
  INV        m1399(.A(mai_mai_n1427_), .Y(mai_mai_n1428_));
  OR3        m1400(.A(mai_mai_n546_), .B(mai_mai_n545_), .C(mai_mai_n113_), .Y(mai_mai_n1429_));
  NA2        m1401(.A(mai_mai_n1121_), .B(mai_mai_n408_), .Y(mai_mai_n1430_));
  OAI220     m1402(.A0(mai_mai_n1430_), .A1(mai_mai_n435_), .B0(mai_mai_n1429_), .B1(mai_mai_n301_), .Y(mai_mai_n1431_));
  AO210      m1403(.A0(mai_mai_n1431_), .A1(mai_mai_n117_), .B0(mai_mai_n1428_), .Y(mai_mai_n1432_));
  NO3        m1404(.A(mai_mai_n1432_), .B(mai_mai_n1426_), .C(mai_mai_n1420_), .Y(mai_mai_n1433_));
  NA4        m1405(.A(mai_mai_n1433_), .B(mai_mai_n1414_), .C(mai_mai_n1388_), .D(mai_mai_n1374_), .Y(mai_mai_n1434_));
  NO2        m1406(.A(mai_mai_n1137_), .B(mai_mai_n111_), .Y(mai_mai_n1435_));
  NO2        m1407(.A(mai_mai_n392_), .B(j), .Y(mai_mai_n1436_));
  NA3        m1408(.A(mai_mai_n1411_), .B(mai_mai_n1355_), .C(mai_mai_n1121_), .Y(mai_mai_n1437_));
  NAi41      m1409(.An(mai_mai_n1398_), .B(mai_mai_n1086_), .C(mai_mai_n169_), .D(mai_mai_n150_), .Y(mai_mai_n1438_));
  NA2        m1410(.A(mai_mai_n1438_), .B(mai_mai_n1437_), .Y(mai_mai_n1439_));
  NA3        m1411(.A(m), .B(mai_mai_n1436_), .C(mai_mai_n158_), .Y(mai_mai_n1440_));
  INV        m1412(.A(mai_mai_n1440_), .Y(mai_mai_n1441_));
  NO2        m1413(.A(mai_mai_n760_), .B(mai_mai_n176_), .Y(mai_mai_n1442_));
  NO3        m1414(.A(mai_mai_n1442_), .B(mai_mai_n1441_), .C(mai_mai_n1439_), .Y(mai_mai_n1443_));
  OR2        m1415(.A(n), .B(i), .Y(mai_mai_n1444_));
  OAI210     m1416(.A0(mai_mai_n1444_), .A1(mai_mai_n1085_), .B0(mai_mai_n49_), .Y(mai_mai_n1445_));
  AOI220     m1417(.A0(mai_mai_n1445_), .A1(mai_mai_n1183_), .B0(mai_mai_n837_), .B1(mai_mai_n197_), .Y(mai_mai_n1446_));
  INV        m1418(.A(mai_mai_n1446_), .Y(mai_mai_n1447_));
  NO2        m1419(.A(mai_mai_n131_), .B(l), .Y(mai_mai_n1448_));
  NO2        m1420(.A(mai_mai_n228_), .B(k), .Y(mai_mai_n1449_));
  OAI210     m1421(.A0(mai_mai_n1449_), .A1(mai_mai_n1398_), .B0(mai_mai_n1448_), .Y(mai_mai_n1450_));
  NO2        m1422(.A(mai_mai_n1450_), .B(mai_mai_n31_), .Y(mai_mai_n1451_));
  NO3        m1423(.A(mai_mai_n1429_), .B(mai_mai_n469_), .C(mai_mai_n355_), .Y(mai_mai_n1452_));
  NO3        m1424(.A(mai_mai_n1452_), .B(mai_mai_n1451_), .C(mai_mai_n1447_), .Y(mai_mai_n1453_));
  INV        m1425(.A(mai_mai_n49_), .Y(mai_mai_n1454_));
  NO3        m1426(.A(mai_mai_n1105_), .B(mai_mai_n1355_), .C(mai_mai_n49_), .Y(mai_mai_n1455_));
  NA2        m1427(.A(mai_mai_n1106_), .B(mai_mai_n1454_), .Y(mai_mai_n1456_));
  NO2        m1428(.A(mai_mai_n1094_), .B(h), .Y(mai_mai_n1457_));
  NA2        m1429(.A(mai_mai_n1457_), .B(d), .Y(mai_mai_n1458_));
  OAI220     m1430(.A0(mai_mai_n1458_), .A1(c), .B0(mai_mai_n1456_), .B1(j), .Y(mai_mai_n1459_));
  NA3        m1431(.A(mai_mai_n1435_), .B(mai_mai_n469_), .C(f), .Y(mai_mai_n1460_));
  NA2        m1432(.A(mai_mai_n181_), .B(mai_mai_n113_), .Y(mai_mai_n1461_));
  NO2        m1433(.A(mai_mai_n1347_), .B(mai_mai_n176_), .Y(mai_mai_n1462_));
  NOi21      m1434(.An(d), .B(f), .Y(mai_mai_n1463_));
  NO2        m1435(.A(mai_mai_n1355_), .B(f), .Y(mai_mai_n1464_));
  INV        m1436(.A(mai_mai_n1459_), .Y(mai_mai_n1465_));
  NA3        m1437(.A(mai_mai_n1465_), .B(mai_mai_n1453_), .C(mai_mai_n1443_), .Y(mai_mai_n1466_));
  NO2        m1438(.A(mai_mai_n1085_), .B(mai_mai_n40_), .Y(mai_mai_n1467_));
  NO2        m1439(.A(mai_mai_n469_), .B(mai_mai_n301_), .Y(mai_mai_n1468_));
  OAI210     m1440(.A0(mai_mai_n1468_), .A1(mai_mai_n1467_), .B0(mai_mai_n1370_), .Y(mai_mai_n1469_));
  OAI210     m1441(.A0(mai_mai_n1421_), .A1(mai_mai_n1358_), .B0(mai_mai_n896_), .Y(mai_mai_n1470_));
  NO2        m1442(.A(mai_mai_n1055_), .B(mai_mai_n131_), .Y(mai_mai_n1471_));
  NA2        m1443(.A(mai_mai_n1471_), .B(mai_mai_n632_), .Y(mai_mai_n1472_));
  NA3        m1444(.A(mai_mai_n1472_), .B(mai_mai_n1470_), .C(mai_mai_n1469_), .Y(mai_mai_n1473_));
  NA2        m1445(.A(mai_mai_n1391_), .B(mai_mai_n1463_), .Y(mai_mai_n1474_));
  NO2        m1446(.A(mai_mai_n1474_), .B(m), .Y(mai_mai_n1475_));
  NO2        m1447(.A(mai_mai_n151_), .B(mai_mai_n183_), .Y(mai_mai_n1476_));
  OAI210     m1448(.A0(mai_mai_n1476_), .A1(mai_mai_n111_), .B0(mai_mai_n1403_), .Y(mai_mai_n1477_));
  INV        m1449(.A(mai_mai_n1477_), .Y(mai_mai_n1478_));
  NO3        m1450(.A(mai_mai_n1478_), .B(mai_mai_n1475_), .C(mai_mai_n1473_), .Y(mai_mai_n1479_));
  NO2        m1451(.A(mai_mai_n1354_), .B(e), .Y(mai_mai_n1480_));
  NA2        m1452(.A(mai_mai_n1480_), .B(mai_mai_n406_), .Y(mai_mai_n1481_));
  NA2        m1453(.A(mai_mai_n1132_), .B(mai_mai_n641_), .Y(mai_mai_n1482_));
  OR3        m1454(.A(mai_mai_n1449_), .B(mai_mai_n1220_), .C(mai_mai_n131_), .Y(mai_mai_n1483_));
  OAI220     m1455(.A0(mai_mai_n1483_), .A1(mai_mai_n1481_), .B0(mai_mai_n1482_), .B1(mai_mai_n444_), .Y(mai_mai_n1484_));
  NO3        m1456(.A(mai_mai_n1429_), .B(mai_mai_n355_), .C(a), .Y(mai_mai_n1485_));
  NO2        m1457(.A(mai_mai_n1485_), .B(mai_mai_n1484_), .Y(mai_mai_n1486_));
  NO2        m1458(.A(mai_mai_n183_), .B(c), .Y(mai_mai_n1487_));
  OAI210     m1459(.A0(mai_mai_n1487_), .A1(mai_mai_n1480_), .B0(mai_mai_n181_), .Y(mai_mai_n1488_));
  AOI220     m1460(.A0(mai_mai_n1488_), .A1(mai_mai_n1087_), .B0(mai_mai_n538_), .B1(mai_mai_n370_), .Y(mai_mai_n1489_));
  AOI210     m1461(.A0(i), .A1(mai_mai_n1387_), .B0(mai_mai_n1455_), .Y(mai_mai_n1490_));
  NO2        m1462(.A(mai_mai_n1423_), .B(f), .Y(mai_mai_n1491_));
  AOI210     m1463(.A0(mai_mai_n1132_), .A1(a), .B0(mai_mai_n1491_), .Y(mai_mai_n1492_));
  OAI220     m1464(.A0(mai_mai_n1492_), .A1(mai_mai_n66_), .B0(mai_mai_n1490_), .B1(mai_mai_n216_), .Y(mai_mai_n1493_));
  OR2        m1465(.A(h), .B(mai_mai_n545_), .Y(mai_mai_n1494_));
  NA2        m1466(.A(mai_mai_n1491_), .B(mai_mai_n1367_), .Y(mai_mai_n1495_));
  OAI220     m1467(.A0(mai_mai_n1495_), .A1(mai_mai_n49_), .B0(mai_mai_n1494_), .B1(mai_mai_n176_), .Y(mai_mai_n1496_));
  NA3        m1468(.A(mai_mai_n1103_), .B(mai_mai_n224_), .C(mai_mai_n65_), .Y(mai_mai_n1497_));
  NA2        m1469(.A(mai_mai_n1359_), .B(mai_mai_n184_), .Y(mai_mai_n1498_));
  NO2        m1470(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1499_));
  OAI210     m1471(.A0(mai_mai_n1423_), .A1(mai_mai_n874_), .B0(mai_mai_n486_), .Y(mai_mai_n1500_));
  OAI210     m1472(.A0(mai_mai_n1500_), .A1(mai_mai_n1106_), .B0(mai_mai_n1499_), .Y(mai_mai_n1501_));
  NO2        m1473(.A(mai_mai_n258_), .B(m), .Y(mai_mai_n1502_));
  NO2        m1474(.A(m), .B(i), .Y(mai_mai_n1503_));
  BUFFER     m1475(.A(mai_mai_n1503_), .Y(mai_mai_n1504_));
  AOI220     m1476(.A0(mai_mai_n1504_), .A1(mai_mai_n1389_), .B0(mai_mai_n1086_), .B1(mai_mai_n1502_), .Y(mai_mai_n1505_));
  NA4        m1477(.A(mai_mai_n1505_), .B(mai_mai_n1501_), .C(mai_mai_n1498_), .D(mai_mai_n1497_), .Y(mai_mai_n1506_));
  NO4        m1478(.A(mai_mai_n1506_), .B(mai_mai_n1496_), .C(mai_mai_n1493_), .D(mai_mai_n1489_), .Y(mai_mai_n1507_));
  NA3        m1479(.A(mai_mai_n1507_), .B(mai_mai_n1486_), .C(mai_mai_n1479_), .Y(mai_mai_n1508_));
  NA3        m1480(.A(mai_mai_n972_), .B(mai_mai_n137_), .C(mai_mai_n46_), .Y(mai_mai_n1509_));
  AOI210     m1481(.A0(mai_mai_n148_), .A1(c), .B0(mai_mai_n1509_), .Y(mai_mai_n1510_));
  INV        m1482(.A(mai_mai_n187_), .Y(mai_mai_n1511_));
  NA2        m1483(.A(mai_mai_n1511_), .B(mai_mai_n1457_), .Y(mai_mai_n1512_));
  OR2        m1484(.A(mai_mai_n132_), .B(mai_mai_n1415_), .Y(mai_mai_n1513_));
  NO2        m1485(.A(mai_mai_n69_), .B(c), .Y(mai_mai_n1514_));
  NO4        m1486(.A(mai_mai_n1379_), .B(mai_mai_n188_), .C(mai_mai_n450_), .D(mai_mai_n45_), .Y(mai_mai_n1515_));
  AOI210     m1487(.A0(mai_mai_n1462_), .A1(mai_mai_n1514_), .B0(mai_mai_n1515_), .Y(mai_mai_n1516_));
  NA3        m1488(.A(mai_mai_n1516_), .B(mai_mai_n1513_), .C(mai_mai_n1512_), .Y(mai_mai_n1517_));
  NO2        m1489(.A(mai_mai_n1517_), .B(mai_mai_n1510_), .Y(mai_mai_n1518_));
  NO4        m1490(.A(mai_mai_n228_), .B(mai_mai_n188_), .C(mai_mai_n263_), .D(k), .Y(mai_mai_n1519_));
  AOI210     m1491(.A0(mai_mai_n156_), .A1(mai_mai_n56_), .B0(mai_mai_n1480_), .Y(mai_mai_n1520_));
  NO2        m1492(.A(mai_mai_n1520_), .B(mai_mai_n1461_), .Y(mai_mai_n1521_));
  NO2        m1493(.A(mai_mai_n1509_), .B(mai_mai_n111_), .Y(mai_mai_n1522_));
  NOi21      m1494(.An(mai_mai_n1359_), .B(e), .Y(mai_mai_n1523_));
  NO4        m1495(.A(mai_mai_n1523_), .B(mai_mai_n1522_), .C(mai_mai_n1521_), .D(mai_mai_n1519_), .Y(mai_mai_n1524_));
  AN2        m1496(.A(mai_mai_n1103_), .B(mai_mai_n1092_), .Y(mai_mai_n1525_));
  AOI220     m1497(.A0(mai_mai_n1503_), .A1(mai_mai_n649_), .B0(mai_mai_n1073_), .B1(mai_mai_n159_), .Y(mai_mai_n1526_));
  NOi31      m1498(.An(mai_mai_n30_), .B(mai_mai_n1526_), .C(n), .Y(mai_mai_n1527_));
  AOI210     m1499(.A0(mai_mai_n1525_), .A1(mai_mai_n1175_), .B0(mai_mai_n1527_), .Y(mai_mai_n1528_));
  NO2        m1500(.A(mai_mai_n1460_), .B(mai_mai_n66_), .Y(mai_mai_n1529_));
  NA2        m1501(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1530_));
  NO2        m1502(.A(mai_mai_n1365_), .B(mai_mai_n119_), .Y(mai_mai_n1531_));
  OAI220     m1503(.A0(mai_mai_n1531_), .A1(mai_mai_n1415_), .B0(mai_mai_n1430_), .B1(mai_mai_n1530_), .Y(mai_mai_n1532_));
  NO2        m1504(.A(mai_mai_n1532_), .B(mai_mai_n1529_), .Y(mai_mai_n1533_));
  NA4        m1505(.A(mai_mai_n1533_), .B(mai_mai_n1528_), .C(mai_mai_n1524_), .D(mai_mai_n1518_), .Y(mai_mai_n1534_));
  OR4        m1506(.A(mai_mai_n1534_), .B(mai_mai_n1508_), .C(mai_mai_n1466_), .D(mai_mai_n1434_), .Y(mai04));
  NOi31      m1507(.An(mai_mai_n1421_), .B(mai_mai_n1422_), .C(mai_mai_n1061_), .Y(mai_mai_n1536_));
  NA2        m1508(.A(mai_mai_n1464_), .B(mai_mai_n837_), .Y(mai_mai_n1537_));
  NO4        m1509(.A(mai_mai_n1537_), .B(mai_mai_n1050_), .C(mai_mai_n487_), .D(j), .Y(mai_mai_n1538_));
  OR3        m1510(.A(mai_mai_n1538_), .B(mai_mai_n1536_), .C(mai_mai_n1079_), .Y(mai_mai_n1539_));
  NO3        m1511(.A(mai_mai_n1367_), .B(mai_mai_n90_), .C(k), .Y(mai_mai_n1540_));
  NA2        m1512(.A(mai_mai_n1540_), .B(mai_mai_n1072_), .Y(mai_mai_n1541_));
  NA2        m1513(.A(mai_mai_n1541_), .B(mai_mai_n1224_), .Y(mai_mai_n1542_));
  NO3        m1514(.A(mai_mai_n1542_), .B(mai_mai_n1539_), .C(mai_mai_n1066_), .Y(mai_mai_n1543_));
  NA3        m1515(.A(mai_mai_n1543_), .B(mai_mai_n1134_), .C(mai_mai_n1109_), .Y(mai05));
  INV        m1516(.A(m), .Y(mai_mai_n1547_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(u), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(u), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(u), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(u), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(u), .Y(men_men_n51_));
  INV        u0023(.A(men_men_n51_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO2        u0025(.A(men_men_n53_), .B(men_men_n43_), .Y(men_men_n54_));
  NO2        u0026(.A(men_men_n54_), .B(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(u), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  NO2        u0034(.A(men_men_n61_), .B(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(u), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(u), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(u), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(u), .Y(men_men_n91_));
  NAi32      u0063(.An(u), .Bn(f), .C(h), .Y(men_men_n92_));
  NAi31      u0064(.An(j), .B(m), .C(l), .Y(men_men_n93_));
  NA2        u0065(.A(m), .B(l), .Y(men_men_n94_));
  NAi31      u0066(.An(k), .B(j), .C(u), .Y(men_men_n95_));
  NO3        u0067(.A(men_men_n95_), .B(men_men_n94_), .C(f), .Y(men_men_n96_));
  AN2        u0068(.A(j), .B(u), .Y(men_men_n97_));
  NOi32      u0069(.An(m), .Bn(l), .C(i), .Y(men_men_n98_));
  NOi21      u0070(.An(u), .B(i), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(j), .C(k), .Y(men_men_n100_));
  AOI220     u0072(.A0(men_men_n100_), .A1(men_men_n99_), .B0(men_men_n98_), .B1(men_men_n97_), .Y(men_men_n101_));
  NO2        u0073(.A(men_men_n101_), .B(f), .Y(men_men_n102_));
  NAi41      u0074(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n103_));
  AN2        u0075(.A(e), .B(b), .Y(men_men_n104_));
  NOi31      u0076(.An(c), .B(h), .C(f), .Y(men_men_n105_));
  NA2        u0077(.A(men_men_n105_), .B(men_men_n104_), .Y(men_men_n106_));
  NO2        u0078(.A(men_men_n106_), .B(men_men_n103_), .Y(men_men_n107_));
  NOi21      u0079(.An(u), .B(f), .Y(men_men_n108_));
  NOi21      u0080(.An(i), .B(h), .Y(men_men_n109_));
  NA3        u0081(.A(men_men_n109_), .B(men_men_n108_), .C(men_men_n36_), .Y(men_men_n110_));
  INV        u0082(.A(a), .Y(men_men_n111_));
  NA2        u0083(.A(men_men_n104_), .B(men_men_n111_), .Y(men_men_n112_));
  INV        u0084(.A(l), .Y(men_men_n113_));
  NOi21      u0085(.An(m), .B(n), .Y(men_men_n114_));
  AN2        u0086(.A(k), .B(h), .Y(men_men_n115_));
  NO2        u0087(.A(men_men_n110_), .B(men_men_n88_), .Y(men_men_n116_));
  INV        u0088(.A(b), .Y(men_men_n117_));
  NA2        u0089(.A(l), .B(j), .Y(men_men_n118_));
  AN2        u0090(.A(k), .B(i), .Y(men_men_n119_));
  NA2        u0091(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NA2        u0092(.A(u), .B(e), .Y(men_men_n121_));
  NOi32      u0093(.An(c), .Bn(a), .C(d), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n114_), .Y(men_men_n123_));
  NO4        u0095(.A(men_men_n123_), .B(men_men_n121_), .C(men_men_n120_), .D(men_men_n117_), .Y(men_men_n124_));
  NO3        u0096(.A(men_men_n124_), .B(men_men_n116_), .C(men_men_n107_), .Y(men_men_n125_));
  OAI210     u0097(.A0(men_men_n101_), .A1(men_men_n88_), .B0(men_men_n125_), .Y(men_men_n126_));
  NOi31      u0098(.An(k), .B(m), .C(j), .Y(men_men_n127_));
  NA3        u0099(.A(men_men_n127_), .B(men_men_n79_), .C(men_men_n78_), .Y(men_men_n128_));
  NOi31      u0100(.An(k), .B(m), .C(i), .Y(men_men_n129_));
  NA3        u0101(.A(men_men_n129_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n130_));
  NA2        u0102(.A(men_men_n130_), .B(men_men_n128_), .Y(men_men_n131_));
  NOi32      u0103(.An(f), .Bn(b), .C(e), .Y(men_men_n132_));
  NAi21      u0104(.An(u), .B(h), .Y(men_men_n133_));
  NAi21      u0105(.An(m), .B(n), .Y(men_men_n134_));
  NAi21      u0106(.An(j), .B(k), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n133_), .Y(men_men_n136_));
  NAi41      u0108(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n137_));
  NAi31      u0109(.An(j), .B(k), .C(h), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n134_), .Y(men_men_n139_));
  AOI210     u0111(.A0(men_men_n136_), .A1(men_men_n132_), .B0(men_men_n139_), .Y(men_men_n140_));
  NO2        u0112(.A(k), .B(j), .Y(men_men_n141_));
  AN2        u0113(.A(k), .B(j), .Y(men_men_n142_));
  NAi21      u0114(.An(c), .B(b), .Y(men_men_n143_));
  NA2        u0115(.A(f), .B(d), .Y(men_men_n144_));
  NA2        u0116(.A(h), .B(c), .Y(men_men_n145_));
  NAi31      u0117(.An(f), .B(e), .C(b), .Y(men_men_n146_));
  NA2        u0118(.A(d), .B(b), .Y(men_men_n147_));
  NAi21      u0119(.An(e), .B(f), .Y(men_men_n148_));
  NO2        u0120(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n149_));
  NA2        u0121(.A(b), .B(a), .Y(men_men_n150_));
  NAi21      u0122(.An(e), .B(u), .Y(men_men_n151_));
  NAi21      u0123(.An(c), .B(d), .Y(men_men_n152_));
  NAi31      u0124(.An(l), .B(k), .C(h), .Y(men_men_n153_));
  NO2        u0125(.A(men_men_n134_), .B(men_men_n153_), .Y(men_men_n154_));
  NA2        u0126(.A(men_men_n154_), .B(men_men_n149_), .Y(men_men_n155_));
  NAi31      u0127(.An(men_men_n131_), .B(men_men_n155_), .C(men_men_n140_), .Y(men_men_n156_));
  NAi31      u0128(.An(e), .B(f), .C(b), .Y(men_men_n157_));
  NOi21      u0129(.An(u), .B(d), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n158_), .B(men_men_n157_), .Y(men_men_n159_));
  NOi21      u0131(.An(h), .B(i), .Y(men_men_n160_));
  NOi21      u0132(.An(k), .B(m), .Y(men_men_n161_));
  NA3        u0133(.A(men_men_n161_), .B(men_men_n160_), .C(n), .Y(men_men_n162_));
  NOi21      u0134(.An(men_men_n159_), .B(men_men_n162_), .Y(men_men_n163_));
  NOi21      u0135(.An(h), .B(u), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n144_), .B(men_men_n143_), .Y(men_men_n165_));
  NA2        u0137(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  NAi31      u0138(.An(l), .B(j), .C(h), .Y(men_men_n167_));
  NOi32      u0139(.An(n), .Bn(k), .C(m), .Y(men_men_n168_));
  NA2        u0140(.A(l), .B(i), .Y(men_men_n169_));
  NA2        u0141(.A(men_men_n169_), .B(men_men_n168_), .Y(men_men_n170_));
  NO2        u0142(.A(men_men_n170_), .B(men_men_n166_), .Y(men_men_n171_));
  NAi31      u0143(.An(d), .B(f), .C(c), .Y(men_men_n172_));
  NAi31      u0144(.An(e), .B(f), .C(c), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  NA2        u0146(.A(j), .B(h), .Y(men_men_n175_));
  OR3        u0147(.A(n), .B(m), .C(k), .Y(men_men_n176_));
  NO2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  NAi32      u0149(.An(m), .Bn(k), .C(n), .Y(men_men_n178_));
  NO2        u0150(.A(men_men_n178_), .B(men_men_n175_), .Y(men_men_n179_));
  AOI220     u0151(.A0(men_men_n179_), .A1(men_men_n159_), .B0(men_men_n177_), .B1(men_men_n174_), .Y(men_men_n180_));
  NO2        u0152(.A(n), .B(m), .Y(men_men_n181_));
  NA2        u0153(.A(men_men_n181_), .B(men_men_n50_), .Y(men_men_n182_));
  NAi21      u0154(.An(f), .B(e), .Y(men_men_n183_));
  NA2        u0155(.A(d), .B(c), .Y(men_men_n184_));
  NO2        u0156(.A(men_men_n184_), .B(men_men_n183_), .Y(men_men_n185_));
  NOi21      u0157(.An(men_men_n185_), .B(men_men_n182_), .Y(men_men_n186_));
  NAi21      u0158(.An(d), .B(c), .Y(men_men_n187_));
  NAi31      u0159(.An(m), .B(n), .C(b), .Y(men_men_n188_));
  NA2        u0160(.A(k), .B(i), .Y(men_men_n189_));
  NAi21      u0161(.An(h), .B(f), .Y(men_men_n190_));
  NO2        u0162(.A(men_men_n190_), .B(men_men_n189_), .Y(men_men_n191_));
  NO2        u0163(.A(men_men_n188_), .B(men_men_n152_), .Y(men_men_n192_));
  NA2        u0164(.A(men_men_n192_), .B(men_men_n191_), .Y(men_men_n193_));
  NOi32      u0165(.An(f), .Bn(c), .C(d), .Y(men_men_n194_));
  NOi32      u0166(.An(f), .Bn(c), .C(e), .Y(men_men_n195_));
  NO2        u0167(.A(men_men_n195_), .B(men_men_n194_), .Y(men_men_n196_));
  NO3        u0168(.A(n), .B(m), .C(j), .Y(men_men_n197_));
  NA2        u0169(.A(men_men_n197_), .B(men_men_n115_), .Y(men_men_n198_));
  AO210      u0170(.A0(men_men_n198_), .A1(men_men_n182_), .B0(men_men_n196_), .Y(men_men_n199_));
  NAi41      u0171(.An(men_men_n186_), .B(men_men_n199_), .C(men_men_n193_), .D(men_men_n180_), .Y(men_men_n200_));
  OR4        u0172(.A(men_men_n200_), .B(men_men_n171_), .C(men_men_n163_), .D(men_men_n156_), .Y(men_men_n201_));
  NO4        u0173(.A(men_men_n201_), .B(men_men_n126_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n202_));
  NA3        u0174(.A(m), .B(men_men_n113_), .C(j), .Y(men_men_n203_));
  NAi31      u0175(.An(n), .B(h), .C(u), .Y(men_men_n204_));
  NO2        u0176(.A(men_men_n204_), .B(men_men_n203_), .Y(men_men_n205_));
  NOi32      u0177(.An(m), .Bn(k), .C(l), .Y(men_men_n206_));
  NA3        u0178(.A(men_men_n206_), .B(men_men_n89_), .C(u), .Y(men_men_n207_));
  NO2        u0179(.A(men_men_n207_), .B(n), .Y(men_men_n208_));
  NOi21      u0180(.An(k), .B(j), .Y(men_men_n209_));
  NA4        u0181(.A(men_men_n209_), .B(men_men_n114_), .C(i), .D(u), .Y(men_men_n210_));
  AN2        u0182(.A(i), .B(u), .Y(men_men_n211_));
  NA3        u0183(.A(men_men_n76_), .B(men_men_n211_), .C(men_men_n114_), .Y(men_men_n212_));
  NA2        u0184(.A(men_men_n212_), .B(men_men_n210_), .Y(men_men_n213_));
  INV        u0185(.A(men_men_n213_), .Y(men_men_n214_));
  NAi41      u0186(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n215_));
  INV        u0187(.A(men_men_n215_), .Y(men_men_n216_));
  INV        u0188(.A(f), .Y(men_men_n217_));
  INV        u0189(.A(u), .Y(men_men_n218_));
  NOi31      u0190(.An(i), .B(j), .C(h), .Y(men_men_n219_));
  NOi21      u0191(.An(l), .B(m), .Y(men_men_n220_));
  NA2        u0192(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n221_));
  NO3        u0193(.A(men_men_n221_), .B(men_men_n218_), .C(men_men_n217_), .Y(men_men_n222_));
  NA2        u0194(.A(men_men_n222_), .B(men_men_n216_), .Y(men_men_n223_));
  OAI210     u0195(.A0(men_men_n214_), .A1(men_men_n32_), .B0(men_men_n223_), .Y(men_men_n224_));
  NOi21      u0196(.An(n), .B(m), .Y(men_men_n225_));
  NOi32      u0197(.An(l), .Bn(i), .C(j), .Y(men_men_n226_));
  NA2        u0198(.A(men_men_n226_), .B(men_men_n225_), .Y(men_men_n227_));
  OA220      u0199(.A0(men_men_n227_), .A1(men_men_n106_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n228_));
  NAi21      u0200(.An(j), .B(h), .Y(men_men_n229_));
  XN2        u0201(.A(i), .B(h), .Y(men_men_n230_));
  NA2        u0202(.A(men_men_n230_), .B(men_men_n229_), .Y(men_men_n231_));
  NOi31      u0203(.An(k), .B(n), .C(m), .Y(men_men_n232_));
  NOi31      u0204(.An(men_men_n232_), .B(men_men_n184_), .C(men_men_n183_), .Y(men_men_n233_));
  NA2        u0205(.A(men_men_n233_), .B(men_men_n231_), .Y(men_men_n234_));
  NAi31      u0206(.An(f), .B(e), .C(c), .Y(men_men_n235_));
  NO4        u0207(.A(men_men_n235_), .B(men_men_n176_), .C(men_men_n175_), .D(men_men_n59_), .Y(men_men_n236_));
  NA3        u0208(.A(e), .B(c), .C(b), .Y(men_men_n237_));
  NAi32      u0209(.An(m), .Bn(i), .C(k), .Y(men_men_n238_));
  INV        u0210(.A(k), .Y(men_men_n239_));
  INV        u0211(.A(men_men_n236_), .Y(men_men_n240_));
  NAi21      u0212(.An(n), .B(a), .Y(men_men_n241_));
  NO2        u0213(.A(men_men_n241_), .B(men_men_n147_), .Y(men_men_n242_));
  NAi41      u0214(.An(u), .B(m), .C(k), .D(h), .Y(men_men_n243_));
  NO2        u0215(.A(men_men_n243_), .B(e), .Y(men_men_n244_));
  NO3        u0216(.A(men_men_n148_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n245_));
  OAI210     u0217(.A0(men_men_n245_), .A1(men_men_n244_), .B0(men_men_n242_), .Y(men_men_n246_));
  AN4        u0218(.A(men_men_n246_), .B(men_men_n240_), .C(men_men_n234_), .D(men_men_n228_), .Y(men_men_n247_));
  OR2        u0219(.A(h), .B(u), .Y(men_men_n248_));
  NO2        u0220(.A(men_men_n248_), .B(men_men_n103_), .Y(men_men_n249_));
  NA2        u0221(.A(men_men_n249_), .B(men_men_n132_), .Y(men_men_n250_));
  NA2        u0222(.A(men_men_n161_), .B(men_men_n109_), .Y(men_men_n251_));
  NO2        u0223(.A(n), .B(a), .Y(men_men_n252_));
  NAi31      u0224(.An(men_men_n243_), .B(men_men_n252_), .C(men_men_n104_), .Y(men_men_n253_));
  NAi21      u0225(.An(h), .B(i), .Y(men_men_n254_));
  NA2        u0226(.A(men_men_n181_), .B(k), .Y(men_men_n255_));
  NO2        u0227(.A(men_men_n255_), .B(men_men_n254_), .Y(men_men_n256_));
  NA2        u0228(.A(men_men_n256_), .B(men_men_n194_), .Y(men_men_n257_));
  NA3        u0229(.A(men_men_n257_), .B(men_men_n253_), .C(men_men_n250_), .Y(men_men_n258_));
  NOi21      u0230(.An(u), .B(e), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n260_));
  NA2        u0232(.A(men_men_n260_), .B(men_men_n259_), .Y(men_men_n261_));
  NOi32      u0233(.An(l), .Bn(j), .C(i), .Y(men_men_n262_));
  AOI210     u0234(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n262_), .Y(men_men_n263_));
  NO2        u0235(.A(men_men_n254_), .B(men_men_n44_), .Y(men_men_n264_));
  NAi21      u0236(.An(f), .B(u), .Y(men_men_n265_));
  NO2        u0237(.A(men_men_n265_), .B(men_men_n65_), .Y(men_men_n266_));
  NO2        u0238(.A(men_men_n69_), .B(men_men_n118_), .Y(men_men_n267_));
  AOI220     u0239(.A0(men_men_n267_), .A1(men_men_n266_), .B0(men_men_n264_), .B1(men_men_n67_), .Y(men_men_n268_));
  OAI210     u0240(.A0(men_men_n263_), .A1(men_men_n261_), .B0(men_men_n268_), .Y(men_men_n269_));
  NO3        u0241(.A(men_men_n135_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n270_));
  NOi41      u0242(.An(men_men_n247_), .B(men_men_n269_), .C(men_men_n258_), .D(men_men_n224_), .Y(men_men_n271_));
  NO4        u0243(.A(men_men_n205_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n272_), .B(men_men_n112_), .Y(men_men_n273_));
  NA3        u0245(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n274_));
  NAi21      u0246(.An(h), .B(u), .Y(men_men_n275_));
  OR4        u0247(.A(men_men_n275_), .B(men_men_n274_), .C(men_men_n227_), .D(e), .Y(men_men_n276_));
  NO2        u0248(.A(men_men_n251_), .B(men_men_n265_), .Y(men_men_n277_));
  NAi31      u0249(.An(u), .B(k), .C(h), .Y(men_men_n278_));
  NO3        u0250(.A(men_men_n134_), .B(men_men_n278_), .C(l), .Y(men_men_n279_));
  NAi31      u0251(.An(e), .B(d), .C(a), .Y(men_men_n280_));
  NA2        u0252(.A(men_men_n279_), .B(men_men_n132_), .Y(men_men_n281_));
  NA2        u0253(.A(men_men_n281_), .B(men_men_n276_), .Y(men_men_n282_));
  NA4        u0254(.A(men_men_n161_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n118_), .Y(men_men_n283_));
  NA3        u0255(.A(men_men_n161_), .B(men_men_n160_), .C(men_men_n86_), .Y(men_men_n284_));
  NO2        u0256(.A(men_men_n284_), .B(men_men_n196_), .Y(men_men_n285_));
  NOi21      u0257(.An(men_men_n283_), .B(men_men_n285_), .Y(men_men_n286_));
  NA3        u0258(.A(e), .B(c), .C(b), .Y(men_men_n287_));
  NO2        u0259(.A(men_men_n60_), .B(men_men_n287_), .Y(men_men_n288_));
  NAi32      u0260(.An(k), .Bn(i), .C(j), .Y(men_men_n289_));
  NAi31      u0261(.An(h), .B(l), .C(i), .Y(men_men_n290_));
  NA3        u0262(.A(men_men_n290_), .B(men_men_n289_), .C(men_men_n167_), .Y(men_men_n291_));
  NOi21      u0263(.An(men_men_n291_), .B(men_men_n49_), .Y(men_men_n292_));
  OAI210     u0264(.A0(men_men_n266_), .A1(men_men_n288_), .B0(men_men_n292_), .Y(men_men_n293_));
  NAi21      u0265(.An(l), .B(k), .Y(men_men_n294_));
  NO2        u0266(.A(men_men_n294_), .B(men_men_n49_), .Y(men_men_n295_));
  NOi21      u0267(.An(l), .B(j), .Y(men_men_n296_));
  NA2        u0268(.A(men_men_n164_), .B(men_men_n296_), .Y(men_men_n297_));
  NAi32      u0269(.An(j), .Bn(h), .C(i), .Y(men_men_n298_));
  NAi21      u0270(.An(m), .B(l), .Y(men_men_n299_));
  NO3        u0271(.A(men_men_n299_), .B(men_men_n298_), .C(men_men_n86_), .Y(men_men_n300_));
  NA2        u0272(.A(h), .B(u), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n168_), .B(men_men_n45_), .Y(men_men_n302_));
  NO2        u0274(.A(men_men_n302_), .B(men_men_n301_), .Y(men_men_n303_));
  OAI210     u0275(.A0(men_men_n303_), .A1(men_men_n300_), .B0(men_men_n165_), .Y(men_men_n304_));
  NA3        u0276(.A(men_men_n304_), .B(men_men_n293_), .C(men_men_n286_), .Y(men_men_n305_));
  NO2        u0277(.A(men_men_n146_), .B(d), .Y(men_men_n306_));
  NA2        u0278(.A(men_men_n306_), .B(men_men_n53_), .Y(men_men_n307_));
  NO2        u0279(.A(men_men_n106_), .B(men_men_n103_), .Y(men_men_n308_));
  NAi32      u0280(.An(n), .Bn(m), .C(l), .Y(men_men_n309_));
  NO2        u0281(.A(men_men_n309_), .B(men_men_n298_), .Y(men_men_n310_));
  NA2        u0282(.A(men_men_n310_), .B(men_men_n185_), .Y(men_men_n311_));
  NO2        u0283(.A(men_men_n123_), .B(men_men_n117_), .Y(men_men_n312_));
  NAi31      u0284(.An(k), .B(l), .C(j), .Y(men_men_n313_));
  OAI210     u0285(.A0(men_men_n294_), .A1(j), .B0(men_men_n313_), .Y(men_men_n314_));
  NOi21      u0286(.An(men_men_n314_), .B(men_men_n121_), .Y(men_men_n315_));
  NA2        u0287(.A(men_men_n315_), .B(men_men_n312_), .Y(men_men_n316_));
  NA3        u0288(.A(men_men_n316_), .B(men_men_n311_), .C(men_men_n307_), .Y(men_men_n317_));
  NO4        u0289(.A(men_men_n317_), .B(men_men_n305_), .C(men_men_n282_), .D(men_men_n273_), .Y(men_men_n318_));
  NA2        u0290(.A(men_men_n256_), .B(men_men_n195_), .Y(men_men_n319_));
  NAi21      u0291(.An(m), .B(k), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n230_), .B(men_men_n320_), .Y(men_men_n321_));
  NAi41      u0293(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n322_));
  NO2        u0294(.A(men_men_n322_), .B(men_men_n151_), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n323_), .B(men_men_n321_), .Y(men_men_n324_));
  NAi31      u0296(.An(i), .B(l), .C(h), .Y(men_men_n325_));
  NA2        u0297(.A(e), .B(c), .Y(men_men_n326_));
  NO3        u0298(.A(men_men_n326_), .B(n), .C(d), .Y(men_men_n327_));
  NOi21      u0299(.An(f), .B(h), .Y(men_men_n328_));
  NA2        u0300(.A(men_men_n328_), .B(men_men_n119_), .Y(men_men_n329_));
  NO2        u0301(.A(men_men_n329_), .B(men_men_n218_), .Y(men_men_n330_));
  NAi31      u0302(.An(d), .B(e), .C(b), .Y(men_men_n331_));
  NO2        u0303(.A(men_men_n134_), .B(men_men_n331_), .Y(men_men_n332_));
  NA2        u0304(.A(men_men_n332_), .B(men_men_n330_), .Y(men_men_n333_));
  NA3        u0305(.A(men_men_n333_), .B(men_men_n324_), .C(men_men_n319_), .Y(men_men_n334_));
  NO4        u0306(.A(men_men_n322_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n218_), .Y(men_men_n335_));
  NA2        u0307(.A(men_men_n252_), .B(men_men_n104_), .Y(men_men_n336_));
  OR2        u0308(.A(men_men_n336_), .B(men_men_n207_), .Y(men_men_n337_));
  NOi31      u0309(.An(l), .B(n), .C(m), .Y(men_men_n338_));
  NA2        u0310(.A(men_men_n338_), .B(men_men_n219_), .Y(men_men_n339_));
  NO2        u0311(.A(men_men_n339_), .B(men_men_n196_), .Y(men_men_n340_));
  NAi32      u0312(.An(men_men_n340_), .Bn(men_men_n335_), .C(men_men_n337_), .Y(men_men_n341_));
  NAi32      u0313(.An(m), .Bn(j), .C(k), .Y(men_men_n342_));
  NAi41      u0314(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n343_));
  OAI210     u0315(.A0(men_men_n215_), .A1(men_men_n342_), .B0(men_men_n343_), .Y(men_men_n344_));
  NOi31      u0316(.An(j), .B(m), .C(k), .Y(men_men_n345_));
  NO2        u0317(.A(men_men_n127_), .B(men_men_n345_), .Y(men_men_n346_));
  AN3        u0318(.A(h), .B(u), .C(f), .Y(men_men_n347_));
  NAi31      u0319(.An(men_men_n346_), .B(men_men_n347_), .C(men_men_n344_), .Y(men_men_n348_));
  NOi32      u0320(.An(m), .Bn(j), .C(l), .Y(men_men_n349_));
  NO2        u0321(.A(men_men_n349_), .B(men_men_n98_), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n299_), .B(men_men_n298_), .Y(men_men_n351_));
  NO2        u0323(.A(men_men_n221_), .B(u), .Y(men_men_n352_));
  NO2        u0324(.A(men_men_n157_), .B(men_men_n86_), .Y(men_men_n353_));
  NA2        u0325(.A(men_men_n353_), .B(men_men_n352_), .Y(men_men_n354_));
  NA2        u0326(.A(men_men_n238_), .B(men_men_n81_), .Y(men_men_n355_));
  NA3        u0327(.A(men_men_n355_), .B(men_men_n347_), .C(men_men_n216_), .Y(men_men_n356_));
  NA3        u0328(.A(men_men_n356_), .B(men_men_n354_), .C(men_men_n348_), .Y(men_men_n357_));
  NA3        u0329(.A(h), .B(u), .C(f), .Y(men_men_n358_));
  NO2        u0330(.A(men_men_n358_), .B(men_men_n77_), .Y(men_men_n359_));
  NA2        u0331(.A(men_men_n343_), .B(men_men_n215_), .Y(men_men_n360_));
  NA2        u0332(.A(men_men_n164_), .B(e), .Y(men_men_n361_));
  NO2        u0333(.A(men_men_n361_), .B(men_men_n41_), .Y(men_men_n362_));
  AOI220     u0334(.A0(men_men_n362_), .A1(men_men_n312_), .B0(men_men_n360_), .B1(men_men_n359_), .Y(men_men_n363_));
  NOi32      u0335(.An(j), .Bn(u), .C(i), .Y(men_men_n364_));
  NA3        u0336(.A(men_men_n364_), .B(men_men_n294_), .C(men_men_n114_), .Y(men_men_n365_));
  AO210      u0337(.A0(men_men_n112_), .A1(men_men_n32_), .B0(men_men_n365_), .Y(men_men_n366_));
  NOi32      u0338(.An(e), .Bn(b), .C(a), .Y(men_men_n367_));
  AN2        u0339(.A(l), .B(j), .Y(men_men_n368_));
  NO2        u0340(.A(men_men_n320_), .B(men_men_n368_), .Y(men_men_n369_));
  NO3        u0341(.A(men_men_n322_), .B(men_men_n72_), .C(men_men_n218_), .Y(men_men_n370_));
  NA3        u0342(.A(men_men_n212_), .B(men_men_n210_), .C(men_men_n35_), .Y(men_men_n371_));
  AOI220     u0343(.A0(men_men_n371_), .A1(men_men_n367_), .B0(men_men_n370_), .B1(men_men_n369_), .Y(men_men_n372_));
  NO2        u0344(.A(men_men_n331_), .B(n), .Y(men_men_n373_));
  NA2        u0345(.A(men_men_n211_), .B(k), .Y(men_men_n374_));
  NA3        u0346(.A(m), .B(men_men_n113_), .C(men_men_n217_), .Y(men_men_n375_));
  NA4        u0347(.A(men_men_n206_), .B(men_men_n89_), .C(u), .D(men_men_n217_), .Y(men_men_n376_));
  OAI210     u0348(.A0(men_men_n375_), .A1(men_men_n374_), .B0(men_men_n376_), .Y(men_men_n377_));
  NAi41      u0349(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n378_));
  NA2        u0350(.A(men_men_n51_), .B(men_men_n114_), .Y(men_men_n379_));
  NO2        u0351(.A(men_men_n379_), .B(men_men_n378_), .Y(men_men_n380_));
  AOI220     u0352(.A0(men_men_n380_), .A1(b), .B0(men_men_n377_), .B1(men_men_n373_), .Y(men_men_n381_));
  NA4        u0353(.A(men_men_n381_), .B(men_men_n372_), .C(men_men_n366_), .D(men_men_n363_), .Y(men_men_n382_));
  NO4        u0354(.A(men_men_n382_), .B(men_men_n357_), .C(men_men_n341_), .D(men_men_n334_), .Y(men_men_n383_));
  NA4        u0355(.A(men_men_n383_), .B(men_men_n318_), .C(men_men_n271_), .D(men_men_n202_), .Y(men10));
  NA3        u0356(.A(m), .B(k), .C(i), .Y(men_men_n385_));
  NO3        u0357(.A(men_men_n385_), .B(j), .C(men_men_n218_), .Y(men_men_n386_));
  NOi21      u0358(.An(e), .B(f), .Y(men_men_n387_));
  NO4        u0359(.A(men_men_n152_), .B(men_men_n387_), .C(n), .D(men_men_n111_), .Y(men_men_n388_));
  NAi31      u0360(.An(b), .B(f), .C(c), .Y(men_men_n389_));
  INV        u0361(.A(men_men_n389_), .Y(men_men_n390_));
  NOi32      u0362(.An(k), .Bn(h), .C(j), .Y(men_men_n391_));
  NA2        u0363(.A(men_men_n391_), .B(men_men_n225_), .Y(men_men_n392_));
  NA2        u0364(.A(men_men_n162_), .B(men_men_n392_), .Y(men_men_n393_));
  NA2        u0365(.A(men_men_n393_), .B(men_men_n390_), .Y(men_men_n394_));
  AN2        u0366(.A(j), .B(h), .Y(men_men_n395_));
  NO3        u0367(.A(n), .B(m), .C(k), .Y(men_men_n396_));
  NA2        u0368(.A(men_men_n396_), .B(men_men_n395_), .Y(men_men_n397_));
  NO3        u0369(.A(men_men_n397_), .B(men_men_n152_), .C(men_men_n217_), .Y(men_men_n398_));
  OR2        u0370(.A(m), .B(k), .Y(men_men_n399_));
  NO2        u0371(.A(men_men_n175_), .B(men_men_n399_), .Y(men_men_n400_));
  NA4        u0372(.A(n), .B(f), .C(c), .D(men_men_n117_), .Y(men_men_n401_));
  NOi21      u0373(.An(men_men_n400_), .B(men_men_n401_), .Y(men_men_n402_));
  NOi32      u0374(.An(d), .Bn(a), .C(c), .Y(men_men_n403_));
  NA2        u0375(.A(men_men_n403_), .B(men_men_n183_), .Y(men_men_n404_));
  NAi21      u0376(.An(i), .B(u), .Y(men_men_n405_));
  NAi31      u0377(.An(k), .B(m), .C(j), .Y(men_men_n406_));
  NO3        u0378(.A(men_men_n406_), .B(men_men_n405_), .C(n), .Y(men_men_n407_));
  NOi21      u0379(.An(men_men_n407_), .B(men_men_n404_), .Y(men_men_n408_));
  NO3        u0380(.A(men_men_n408_), .B(men_men_n402_), .C(men_men_n398_), .Y(men_men_n409_));
  NO2        u0381(.A(men_men_n401_), .B(men_men_n299_), .Y(men_men_n410_));
  NOi32      u0382(.An(f), .Bn(d), .C(c), .Y(men_men_n411_));
  AOI220     u0383(.A0(men_men_n411_), .A1(men_men_n310_), .B0(men_men_n410_), .B1(men_men_n219_), .Y(men_men_n412_));
  NA3        u0384(.A(men_men_n412_), .B(men_men_n409_), .C(men_men_n394_), .Y(men_men_n413_));
  NO2        u0385(.A(men_men_n59_), .B(men_men_n117_), .Y(men_men_n414_));
  NA2        u0386(.A(men_men_n252_), .B(men_men_n414_), .Y(men_men_n415_));
  INV        u0387(.A(e), .Y(men_men_n416_));
  NA2        u0388(.A(men_men_n46_), .B(e), .Y(men_men_n417_));
  OAI220     u0389(.A0(men_men_n417_), .A1(men_men_n203_), .B0(men_men_n207_), .B1(men_men_n416_), .Y(men_men_n418_));
  AN2        u0390(.A(u), .B(e), .Y(men_men_n419_));
  NA3        u0391(.A(men_men_n419_), .B(men_men_n206_), .C(i), .Y(men_men_n420_));
  OAI210     u0392(.A0(men_men_n91_), .A1(men_men_n416_), .B0(men_men_n420_), .Y(men_men_n421_));
  NO2        u0393(.A(men_men_n101_), .B(men_men_n416_), .Y(men_men_n422_));
  NO3        u0394(.A(men_men_n422_), .B(men_men_n421_), .C(men_men_n418_), .Y(men_men_n423_));
  NOi32      u0395(.An(h), .Bn(e), .C(u), .Y(men_men_n424_));
  NA3        u0396(.A(men_men_n424_), .B(men_men_n296_), .C(m), .Y(men_men_n425_));
  NOi21      u0397(.An(u), .B(h), .Y(men_men_n426_));
  AN3        u0398(.A(m), .B(l), .C(i), .Y(men_men_n427_));
  NA3        u0399(.A(men_men_n427_), .B(men_men_n426_), .C(e), .Y(men_men_n428_));
  AN3        u0400(.A(h), .B(u), .C(e), .Y(men_men_n429_));
  NA2        u0401(.A(men_men_n429_), .B(men_men_n98_), .Y(men_men_n430_));
  AN3        u0402(.A(men_men_n430_), .B(men_men_n428_), .C(men_men_n425_), .Y(men_men_n431_));
  AOI210     u0403(.A0(men_men_n431_), .A1(men_men_n423_), .B0(men_men_n415_), .Y(men_men_n432_));
  NA3        u0404(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n433_));
  NO2        u0405(.A(men_men_n433_), .B(men_men_n415_), .Y(men_men_n434_));
  NA3        u0406(.A(men_men_n403_), .B(men_men_n183_), .C(men_men_n86_), .Y(men_men_n435_));
  NAi31      u0407(.An(b), .B(c), .C(a), .Y(men_men_n436_));
  NO2        u0408(.A(men_men_n436_), .B(n), .Y(men_men_n437_));
  NA2        u0409(.A(men_men_n51_), .B(m), .Y(men_men_n438_));
  NO2        u0410(.A(men_men_n438_), .B(men_men_n148_), .Y(men_men_n439_));
  NA2        u0411(.A(men_men_n439_), .B(men_men_n437_), .Y(men_men_n440_));
  INV        u0412(.A(men_men_n440_), .Y(men_men_n441_));
  NO4        u0413(.A(men_men_n441_), .B(men_men_n434_), .C(men_men_n432_), .D(men_men_n413_), .Y(men_men_n442_));
  NA2        u0414(.A(i), .B(u), .Y(men_men_n443_));
  NO3        u0415(.A(men_men_n280_), .B(men_men_n443_), .C(c), .Y(men_men_n444_));
  NOi21      u0416(.An(a), .B(n), .Y(men_men_n445_));
  NOi21      u0417(.An(d), .B(c), .Y(men_men_n446_));
  NA2        u0418(.A(men_men_n446_), .B(men_men_n445_), .Y(men_men_n447_));
  NA3        u0419(.A(i), .B(u), .C(f), .Y(men_men_n448_));
  OR2        u0420(.A(men_men_n448_), .B(men_men_n71_), .Y(men_men_n449_));
  NA3        u0421(.A(men_men_n427_), .B(men_men_n426_), .C(men_men_n183_), .Y(men_men_n450_));
  AOI210     u0422(.A0(men_men_n450_), .A1(men_men_n449_), .B0(men_men_n447_), .Y(men_men_n451_));
  AOI210     u0423(.A0(men_men_n444_), .A1(men_men_n295_), .B0(men_men_n451_), .Y(men_men_n452_));
  OR2        u0424(.A(n), .B(m), .Y(men_men_n453_));
  NO2        u0425(.A(men_men_n453_), .B(men_men_n153_), .Y(men_men_n454_));
  NO2        u0426(.A(men_men_n184_), .B(men_men_n148_), .Y(men_men_n455_));
  OAI210     u0427(.A0(men_men_n454_), .A1(men_men_n177_), .B0(men_men_n455_), .Y(men_men_n456_));
  INV        u0428(.A(men_men_n379_), .Y(men_men_n457_));
  NA3        u0429(.A(men_men_n457_), .B(men_men_n367_), .C(d), .Y(men_men_n458_));
  NO2        u0430(.A(men_men_n436_), .B(men_men_n49_), .Y(men_men_n459_));
  NO3        u0431(.A(men_men_n66_), .B(men_men_n113_), .C(e), .Y(men_men_n460_));
  NAi21      u0432(.An(k), .B(j), .Y(men_men_n461_));
  NA3        u0433(.A(i), .B(men_men_n460_), .C(men_men_n459_), .Y(men_men_n462_));
  NAi21      u0434(.An(e), .B(d), .Y(men_men_n463_));
  INV        u0435(.A(men_men_n463_), .Y(men_men_n464_));
  NO2        u0436(.A(men_men_n255_), .B(men_men_n217_), .Y(men_men_n465_));
  NA3        u0437(.A(men_men_n465_), .B(men_men_n464_), .C(men_men_n231_), .Y(men_men_n466_));
  NA4        u0438(.A(men_men_n466_), .B(men_men_n462_), .C(men_men_n458_), .D(men_men_n456_), .Y(men_men_n467_));
  NO2        u0439(.A(men_men_n339_), .B(men_men_n217_), .Y(men_men_n468_));
  NA2        u0440(.A(men_men_n468_), .B(men_men_n464_), .Y(men_men_n469_));
  NOi31      u0441(.An(n), .B(m), .C(k), .Y(men_men_n470_));
  AOI220     u0442(.A0(men_men_n470_), .A1(men_men_n395_), .B0(men_men_n225_), .B1(men_men_n50_), .Y(men_men_n471_));
  NAi31      u0443(.An(u), .B(f), .C(c), .Y(men_men_n472_));
  OR3        u0444(.A(men_men_n472_), .B(men_men_n471_), .C(e), .Y(men_men_n473_));
  NA3        u0445(.A(men_men_n473_), .B(men_men_n469_), .C(men_men_n311_), .Y(men_men_n474_));
  NOi41      u0446(.An(men_men_n452_), .B(men_men_n474_), .C(men_men_n467_), .D(men_men_n269_), .Y(men_men_n475_));
  NOi32      u0447(.An(c), .Bn(a), .C(b), .Y(men_men_n476_));
  NA2        u0448(.A(men_men_n476_), .B(men_men_n114_), .Y(men_men_n477_));
  INV        u0449(.A(men_men_n278_), .Y(men_men_n478_));
  AN2        u0450(.A(e), .B(d), .Y(men_men_n479_));
  NA2        u0451(.A(men_men_n479_), .B(men_men_n478_), .Y(men_men_n480_));
  INV        u0452(.A(men_men_n148_), .Y(men_men_n481_));
  NO2        u0453(.A(men_men_n133_), .B(men_men_n41_), .Y(men_men_n482_));
  NO2        u0454(.A(men_men_n66_), .B(e), .Y(men_men_n483_));
  NOi31      u0455(.An(j), .B(k), .C(i), .Y(men_men_n484_));
  NOi21      u0456(.An(men_men_n167_), .B(men_men_n484_), .Y(men_men_n485_));
  NA4        u0457(.A(men_men_n325_), .B(men_men_n485_), .C(men_men_n263_), .D(men_men_n120_), .Y(men_men_n486_));
  AOI220     u0458(.A0(men_men_n486_), .A1(men_men_n483_), .B0(men_men_n482_), .B1(men_men_n481_), .Y(men_men_n487_));
  AOI210     u0459(.A0(men_men_n487_), .A1(men_men_n480_), .B0(men_men_n477_), .Y(men_men_n488_));
  NO2        u0460(.A(men_men_n213_), .B(men_men_n208_), .Y(men_men_n489_));
  NOi21      u0461(.An(a), .B(b), .Y(men_men_n490_));
  NA3        u0462(.A(e), .B(d), .C(c), .Y(men_men_n491_));
  NAi21      u0463(.An(men_men_n491_), .B(men_men_n490_), .Y(men_men_n492_));
  NO2        u0464(.A(men_men_n435_), .B(men_men_n207_), .Y(men_men_n493_));
  NOi21      u0465(.An(men_men_n492_), .B(men_men_n493_), .Y(men_men_n494_));
  AOI210     u0466(.A0(men_men_n272_), .A1(men_men_n489_), .B0(men_men_n494_), .Y(men_men_n495_));
  NO4        u0467(.A(men_men_n190_), .B(men_men_n103_), .C(men_men_n56_), .D(b), .Y(men_men_n496_));
  NA2        u0468(.A(men_men_n390_), .B(men_men_n154_), .Y(men_men_n497_));
  OR2        u0469(.A(k), .B(j), .Y(men_men_n498_));
  NA2        u0470(.A(l), .B(k), .Y(men_men_n499_));
  NA3        u0471(.A(men_men_n499_), .B(men_men_n498_), .C(men_men_n225_), .Y(men_men_n500_));
  AOI210     u0472(.A0(men_men_n238_), .A1(men_men_n342_), .B0(men_men_n86_), .Y(men_men_n501_));
  NOi21      u0473(.An(men_men_n500_), .B(men_men_n501_), .Y(men_men_n502_));
  OR3        u0474(.A(men_men_n502_), .B(men_men_n145_), .C(men_men_n137_), .Y(men_men_n503_));
  NA3        u0475(.A(men_men_n283_), .B(men_men_n130_), .C(men_men_n128_), .Y(men_men_n504_));
  NA2        u0476(.A(men_men_n403_), .B(men_men_n114_), .Y(men_men_n505_));
  NO4        u0477(.A(men_men_n505_), .B(men_men_n95_), .C(men_men_n113_), .D(e), .Y(men_men_n506_));
  NO3        u0478(.A(men_men_n435_), .B(men_men_n93_), .C(men_men_n133_), .Y(men_men_n507_));
  NO3        u0479(.A(men_men_n507_), .B(men_men_n506_), .C(men_men_n504_), .Y(men_men_n508_));
  NA3        u0480(.A(men_men_n508_), .B(men_men_n503_), .C(men_men_n497_), .Y(men_men_n509_));
  NO4        u0481(.A(men_men_n509_), .B(men_men_n496_), .C(men_men_n495_), .D(men_men_n488_), .Y(men_men_n510_));
  NA2        u0482(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n511_));
  NAi31      u0483(.An(j), .B(l), .C(i), .Y(men_men_n512_));
  OAI210     u0484(.A0(men_men_n512_), .A1(men_men_n134_), .B0(men_men_n103_), .Y(men_men_n513_));
  NO3        u0485(.A(men_men_n404_), .B(men_men_n350_), .C(men_men_n204_), .Y(men_men_n514_));
  NO2        u0486(.A(men_men_n404_), .B(men_men_n379_), .Y(men_men_n515_));
  NO4        u0487(.A(men_men_n515_), .B(men_men_n514_), .C(men_men_n186_), .D(men_men_n308_), .Y(men_men_n516_));
  NA3        u0488(.A(men_men_n516_), .B(men_men_n511_), .C(men_men_n247_), .Y(men_men_n517_));
  OAI210     u0489(.A0(men_men_n129_), .A1(men_men_n127_), .B0(n), .Y(men_men_n518_));
  NO2        u0490(.A(men_men_n518_), .B(men_men_n133_), .Y(men_men_n519_));
  OR2        u0491(.A(men_men_n300_), .B(men_men_n249_), .Y(men_men_n520_));
  OA210      u0492(.A0(men_men_n520_), .A1(men_men_n519_), .B0(men_men_n195_), .Y(men_men_n521_));
  XO2        u0493(.A(i), .B(h), .Y(men_men_n522_));
  NA3        u0494(.A(men_men_n522_), .B(men_men_n161_), .C(n), .Y(men_men_n523_));
  NAi41      u0495(.An(men_men_n300_), .B(men_men_n523_), .C(men_men_n471_), .D(men_men_n392_), .Y(men_men_n524_));
  NOi32      u0496(.An(men_men_n524_), .Bn(men_men_n483_), .C(men_men_n274_), .Y(men_men_n525_));
  NAi31      u0497(.An(c), .B(f), .C(d), .Y(men_men_n526_));
  AOI210     u0498(.A0(men_men_n284_), .A1(men_men_n198_), .B0(men_men_n526_), .Y(men_men_n527_));
  NOi21      u0499(.An(men_men_n84_), .B(men_men_n527_), .Y(men_men_n528_));
  NA3        u0500(.A(men_men_n388_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n529_));
  NA2        u0501(.A(men_men_n232_), .B(men_men_n109_), .Y(men_men_n530_));
  AOI210     u0502(.A0(men_men_n530_), .A1(men_men_n182_), .B0(men_men_n526_), .Y(men_men_n531_));
  AOI210     u0503(.A0(men_men_n365_), .A1(men_men_n35_), .B0(men_men_n492_), .Y(men_men_n532_));
  NOi31      u0504(.An(men_men_n529_), .B(men_men_n532_), .C(men_men_n531_), .Y(men_men_n533_));
  AN2        u0505(.A(men_men_n292_), .B(men_men_n266_), .Y(men_men_n534_));
  NA3        u0506(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n535_));
  NO2        u0507(.A(men_men_n535_), .B(men_men_n447_), .Y(men_men_n536_));
  INV        u0508(.A(men_men_n536_), .Y(men_men_n537_));
  NAi41      u0509(.An(men_men_n534_), .B(men_men_n537_), .C(men_men_n533_), .D(men_men_n528_), .Y(men_men_n538_));
  NO4        u0510(.A(men_men_n538_), .B(men_men_n525_), .C(men_men_n521_), .D(men_men_n517_), .Y(men_men_n539_));
  NA4        u0511(.A(men_men_n539_), .B(men_men_n510_), .C(men_men_n475_), .D(men_men_n442_), .Y(men11));
  NO2        u0512(.A(men_men_n73_), .B(f), .Y(men_men_n541_));
  NA2        u0513(.A(j), .B(u), .Y(men_men_n542_));
  NAi31      u0514(.An(i), .B(m), .C(l), .Y(men_men_n543_));
  NA3        u0515(.A(m), .B(k), .C(j), .Y(men_men_n544_));
  OAI220     u0516(.A0(men_men_n544_), .A1(men_men_n133_), .B0(men_men_n543_), .B1(men_men_n542_), .Y(men_men_n545_));
  NA2        u0517(.A(men_men_n545_), .B(men_men_n541_), .Y(men_men_n546_));
  NOi32      u0518(.An(e), .Bn(b), .C(f), .Y(men_men_n547_));
  NA2        u0519(.A(men_men_n262_), .B(men_men_n114_), .Y(men_men_n548_));
  NA2        u0520(.A(men_men_n46_), .B(j), .Y(men_men_n549_));
  NO2        u0521(.A(men_men_n549_), .B(men_men_n302_), .Y(men_men_n550_));
  NAi31      u0522(.An(d), .B(e), .C(a), .Y(men_men_n551_));
  NO2        u0523(.A(men_men_n551_), .B(n), .Y(men_men_n552_));
  AOI220     u0524(.A0(men_men_n552_), .A1(men_men_n102_), .B0(men_men_n550_), .B1(men_men_n547_), .Y(men_men_n553_));
  NAi41      u0525(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n554_));
  AN2        u0526(.A(men_men_n554_), .B(men_men_n378_), .Y(men_men_n555_));
  AOI210     u0527(.A0(men_men_n555_), .A1(men_men_n404_), .B0(men_men_n275_), .Y(men_men_n556_));
  NA2        u0528(.A(j), .B(i), .Y(men_men_n557_));
  NAi31      u0529(.An(n), .B(m), .C(k), .Y(men_men_n558_));
  NO3        u0530(.A(men_men_n558_), .B(men_men_n557_), .C(men_men_n113_), .Y(men_men_n559_));
  NO4        u0531(.A(n), .B(d), .C(men_men_n117_), .D(a), .Y(men_men_n560_));
  OR2        u0532(.A(n), .B(c), .Y(men_men_n561_));
  NO2        u0533(.A(men_men_n561_), .B(men_men_n150_), .Y(men_men_n562_));
  NO2        u0534(.A(men_men_n562_), .B(men_men_n560_), .Y(men_men_n563_));
  NOi32      u0535(.An(u), .Bn(f), .C(i), .Y(men_men_n564_));
  AOI220     u0536(.A0(men_men_n564_), .A1(men_men_n100_), .B0(men_men_n545_), .B1(f), .Y(men_men_n565_));
  NO2        u0537(.A(men_men_n278_), .B(men_men_n49_), .Y(men_men_n566_));
  NO2        u0538(.A(men_men_n565_), .B(men_men_n563_), .Y(men_men_n567_));
  AOI210     u0539(.A0(men_men_n559_), .A1(men_men_n556_), .B0(men_men_n567_), .Y(men_men_n568_));
  NA2        u0540(.A(men_men_n142_), .B(men_men_n34_), .Y(men_men_n569_));
  OAI220     u0541(.A0(men_men_n569_), .A1(m), .B0(men_men_n549_), .B1(men_men_n238_), .Y(men_men_n570_));
  NOi41      u0542(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n571_));
  NAi32      u0543(.An(e), .Bn(b), .C(c), .Y(men_men_n572_));
  OR2        u0544(.A(men_men_n572_), .B(men_men_n86_), .Y(men_men_n573_));
  AN2        u0545(.A(men_men_n343_), .B(men_men_n322_), .Y(men_men_n574_));
  NA2        u0546(.A(men_men_n574_), .B(men_men_n573_), .Y(men_men_n575_));
  OA210      u0547(.A0(men_men_n575_), .A1(men_men_n571_), .B0(men_men_n570_), .Y(men_men_n576_));
  OAI220     u0548(.A0(men_men_n406_), .A1(men_men_n405_), .B0(men_men_n543_), .B1(men_men_n542_), .Y(men_men_n577_));
  NAi31      u0549(.An(d), .B(c), .C(a), .Y(men_men_n578_));
  NO2        u0550(.A(men_men_n578_), .B(n), .Y(men_men_n579_));
  NA3        u0551(.A(men_men_n579_), .B(men_men_n577_), .C(e), .Y(men_men_n580_));
  NO3        u0552(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n218_), .Y(men_men_n581_));
  NO2        u0553(.A(men_men_n235_), .B(men_men_n111_), .Y(men_men_n582_));
  OAI210     u0554(.A0(men_men_n581_), .A1(men_men_n407_), .B0(men_men_n582_), .Y(men_men_n583_));
  NA2        u0555(.A(men_men_n583_), .B(men_men_n580_), .Y(men_men_n584_));
  NO2        u0556(.A(men_men_n280_), .B(n), .Y(men_men_n585_));
  NO2        u0557(.A(men_men_n437_), .B(men_men_n585_), .Y(men_men_n586_));
  NA2        u0558(.A(men_men_n577_), .B(f), .Y(men_men_n587_));
  NAi32      u0559(.An(d), .Bn(a), .C(b), .Y(men_men_n588_));
  NO2        u0560(.A(men_men_n588_), .B(men_men_n49_), .Y(men_men_n589_));
  NA2        u0561(.A(h), .B(f), .Y(men_men_n590_));
  NO2        u0562(.A(men_men_n590_), .B(men_men_n95_), .Y(men_men_n591_));
  NO3        u0563(.A(men_men_n178_), .B(men_men_n175_), .C(u), .Y(men_men_n592_));
  AOI220     u0564(.A0(men_men_n592_), .A1(men_men_n58_), .B0(men_men_n591_), .B1(men_men_n589_), .Y(men_men_n593_));
  OAI210     u0565(.A0(men_men_n587_), .A1(men_men_n586_), .B0(men_men_n593_), .Y(men_men_n594_));
  AN3        u0566(.A(j), .B(h), .C(u), .Y(men_men_n595_));
  NO2        u0567(.A(men_men_n147_), .B(c), .Y(men_men_n596_));
  NA3        u0568(.A(men_men_n596_), .B(men_men_n595_), .C(men_men_n470_), .Y(men_men_n597_));
  NA3        u0569(.A(f), .B(d), .C(b), .Y(men_men_n598_));
  NO4        u0570(.A(men_men_n598_), .B(men_men_n178_), .C(men_men_n175_), .D(u), .Y(men_men_n599_));
  INV        u0571(.A(men_men_n597_), .Y(men_men_n600_));
  NO4        u0572(.A(men_men_n600_), .B(men_men_n594_), .C(men_men_n584_), .D(men_men_n576_), .Y(men_men_n601_));
  AN4        u0573(.A(men_men_n601_), .B(men_men_n568_), .C(men_men_n553_), .D(men_men_n546_), .Y(men_men_n602_));
  INV        u0574(.A(k), .Y(men_men_n603_));
  NA3        u0575(.A(l), .B(men_men_n603_), .C(i), .Y(men_men_n604_));
  INV        u0576(.A(men_men_n604_), .Y(men_men_n605_));
  NA4        u0577(.A(men_men_n403_), .B(men_men_n426_), .C(men_men_n183_), .D(men_men_n114_), .Y(men_men_n606_));
  NAi32      u0578(.An(h), .Bn(f), .C(u), .Y(men_men_n607_));
  NAi41      u0579(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n608_));
  OAI210     u0580(.A0(men_men_n551_), .A1(n), .B0(men_men_n608_), .Y(men_men_n609_));
  NA2        u0581(.A(men_men_n609_), .B(m), .Y(men_men_n610_));
  NAi31      u0582(.An(h), .B(u), .C(f), .Y(men_men_n611_));
  OR3        u0583(.A(men_men_n611_), .B(men_men_n280_), .C(men_men_n49_), .Y(men_men_n612_));
  NA4        u0584(.A(men_men_n426_), .B(men_men_n122_), .C(men_men_n114_), .D(e), .Y(men_men_n613_));
  AN2        u0585(.A(men_men_n613_), .B(men_men_n612_), .Y(men_men_n614_));
  OA210      u0586(.A0(men_men_n610_), .A1(men_men_n607_), .B0(men_men_n614_), .Y(men_men_n615_));
  NA2        u0587(.A(men_men_n615_), .B(men_men_n606_), .Y(men_men_n616_));
  NAi31      u0588(.An(f), .B(h), .C(u), .Y(men_men_n617_));
  NO4        u0589(.A(men_men_n313_), .B(men_men_n617_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n618_));
  NOi32      u0590(.An(b), .Bn(a), .C(c), .Y(men_men_n619_));
  NOi32      u0591(.An(d), .Bn(a), .C(e), .Y(men_men_n620_));
  NO2        u0592(.A(n), .B(c), .Y(men_men_n621_));
  NA3        u0593(.A(men_men_n621_), .B(men_men_n29_), .C(m), .Y(men_men_n622_));
  NOi32      u0594(.An(e), .Bn(a), .C(d), .Y(men_men_n623_));
  AOI210     u0595(.A0(men_men_n29_), .A1(d), .B0(men_men_n623_), .Y(men_men_n624_));
  AOI210     u0596(.A0(men_men_n616_), .A1(men_men_n605_), .B0(men_men_n618_), .Y(men_men_n625_));
  NO3        u0597(.A(men_men_n320_), .B(men_men_n61_), .C(n), .Y(men_men_n626_));
  NA3        u0598(.A(men_men_n526_), .B(men_men_n173_), .C(men_men_n172_), .Y(men_men_n627_));
  NA2        u0599(.A(men_men_n472_), .B(men_men_n235_), .Y(men_men_n628_));
  OR2        u0600(.A(men_men_n628_), .B(men_men_n627_), .Y(men_men_n629_));
  NA2        u0601(.A(men_men_n76_), .B(men_men_n114_), .Y(men_men_n630_));
  NO2        u0602(.A(men_men_n630_), .B(men_men_n45_), .Y(men_men_n631_));
  AOI220     u0603(.A0(men_men_n631_), .A1(men_men_n556_), .B0(men_men_n629_), .B1(men_men_n626_), .Y(men_men_n632_));
  NO2        u0604(.A(men_men_n632_), .B(men_men_n89_), .Y(men_men_n633_));
  NA3        u0605(.A(men_men_n571_), .B(men_men_n345_), .C(men_men_n46_), .Y(men_men_n634_));
  NOi32      u0606(.An(e), .Bn(c), .C(f), .Y(men_men_n635_));
  NOi21      u0607(.An(f), .B(u), .Y(men_men_n636_));
  NO2        u0608(.A(men_men_n636_), .B(men_men_n215_), .Y(men_men_n637_));
  AOI220     u0609(.A0(men_men_n637_), .A1(men_men_n400_), .B0(men_men_n635_), .B1(men_men_n177_), .Y(men_men_n638_));
  NA3        u0610(.A(men_men_n638_), .B(men_men_n634_), .C(men_men_n180_), .Y(men_men_n639_));
  AOI210     u0611(.A0(men_men_n555_), .A1(men_men_n404_), .B0(men_men_n301_), .Y(men_men_n640_));
  NA2        u0612(.A(men_men_n640_), .B(men_men_n267_), .Y(men_men_n641_));
  NOi21      u0613(.An(j), .B(l), .Y(men_men_n642_));
  NAi21      u0614(.An(k), .B(h), .Y(men_men_n643_));
  NO2        u0615(.A(men_men_n643_), .B(men_men_n265_), .Y(men_men_n644_));
  NOi31      u0616(.An(m), .B(n), .C(k), .Y(men_men_n645_));
  NA2        u0617(.A(men_men_n642_), .B(men_men_n645_), .Y(men_men_n646_));
  AOI210     u0618(.A0(men_men_n404_), .A1(men_men_n378_), .B0(men_men_n301_), .Y(men_men_n647_));
  NAi21      u0619(.An(men_men_n646_), .B(men_men_n647_), .Y(men_men_n648_));
  NO2        u0620(.A(men_men_n280_), .B(men_men_n49_), .Y(men_men_n649_));
  NO2        u0621(.A(men_men_n551_), .B(men_men_n49_), .Y(men_men_n650_));
  NA2        u0622(.A(men_men_n649_), .B(men_men_n591_), .Y(men_men_n651_));
  NA3        u0623(.A(men_men_n651_), .B(men_men_n648_), .C(men_men_n641_), .Y(men_men_n652_));
  NA2        u0624(.A(men_men_n109_), .B(men_men_n36_), .Y(men_men_n653_));
  NO2        u0625(.A(k), .B(men_men_n218_), .Y(men_men_n654_));
  INV        u0626(.A(men_men_n367_), .Y(men_men_n655_));
  NO2        u0627(.A(men_men_n655_), .B(n), .Y(men_men_n656_));
  NAi31      u0628(.An(men_men_n653_), .B(men_men_n656_), .C(men_men_n654_), .Y(men_men_n657_));
  NO2        u0629(.A(men_men_n549_), .B(men_men_n178_), .Y(men_men_n658_));
  NA3        u0630(.A(men_men_n572_), .B(men_men_n274_), .C(men_men_n146_), .Y(men_men_n659_));
  NA2        u0631(.A(men_men_n522_), .B(men_men_n161_), .Y(men_men_n660_));
  NO3        u0632(.A(men_men_n401_), .B(men_men_n660_), .C(men_men_n89_), .Y(men_men_n661_));
  AOI210     u0633(.A0(men_men_n659_), .A1(men_men_n658_), .B0(men_men_n661_), .Y(men_men_n662_));
  AN3        u0634(.A(f), .B(d), .C(b), .Y(men_men_n663_));
  OAI210     u0635(.A0(men_men_n663_), .A1(men_men_n132_), .B0(n), .Y(men_men_n664_));
  NA3        u0636(.A(men_men_n522_), .B(men_men_n161_), .C(men_men_n218_), .Y(men_men_n665_));
  AOI210     u0637(.A0(men_men_n664_), .A1(men_men_n237_), .B0(men_men_n665_), .Y(men_men_n666_));
  NAi31      u0638(.An(m), .B(n), .C(k), .Y(men_men_n667_));
  OR2        u0639(.A(men_men_n137_), .B(men_men_n61_), .Y(men_men_n668_));
  OAI210     u0640(.A0(men_men_n668_), .A1(men_men_n667_), .B0(men_men_n253_), .Y(men_men_n669_));
  OAI210     u0641(.A0(men_men_n669_), .A1(men_men_n666_), .B0(j), .Y(men_men_n670_));
  NA3        u0642(.A(men_men_n670_), .B(men_men_n662_), .C(men_men_n657_), .Y(men_men_n671_));
  NO4        u0643(.A(men_men_n671_), .B(men_men_n652_), .C(men_men_n639_), .D(men_men_n633_), .Y(men_men_n672_));
  NA2        u0644(.A(men_men_n388_), .B(men_men_n164_), .Y(men_men_n673_));
  NAi31      u0645(.An(u), .B(h), .C(f), .Y(men_men_n674_));
  OR3        u0646(.A(men_men_n674_), .B(men_men_n280_), .C(n), .Y(men_men_n675_));
  OA210      u0647(.A0(men_men_n551_), .A1(n), .B0(men_men_n608_), .Y(men_men_n676_));
  NA3        u0648(.A(men_men_n424_), .B(men_men_n122_), .C(men_men_n86_), .Y(men_men_n677_));
  OAI210     u0649(.A0(men_men_n676_), .A1(men_men_n92_), .B0(men_men_n677_), .Y(men_men_n678_));
  NOi21      u0650(.An(men_men_n675_), .B(men_men_n678_), .Y(men_men_n679_));
  AOI210     u0651(.A0(men_men_n679_), .A1(men_men_n673_), .B0(men_men_n544_), .Y(men_men_n680_));
  NO3        u0652(.A(u), .B(men_men_n217_), .C(men_men_n56_), .Y(men_men_n681_));
  NAi21      u0653(.An(h), .B(j), .Y(men_men_n682_));
  NO2        u0654(.A(men_men_n530_), .B(men_men_n89_), .Y(men_men_n683_));
  OAI210     u0655(.A0(men_men_n683_), .A1(men_men_n400_), .B0(men_men_n681_), .Y(men_men_n684_));
  OR2        u0656(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n685_));
  NA3        u0657(.A(men_men_n541_), .B(men_men_n100_), .C(men_men_n99_), .Y(men_men_n686_));
  AN2        u0658(.A(h), .B(f), .Y(men_men_n687_));
  NA2        u0659(.A(men_men_n687_), .B(men_men_n37_), .Y(men_men_n688_));
  NA2        u0660(.A(men_men_n100_), .B(men_men_n46_), .Y(men_men_n689_));
  OAI220     u0661(.A0(men_men_n689_), .A1(men_men_n336_), .B0(men_men_n688_), .B1(men_men_n477_), .Y(men_men_n690_));
  AOI210     u0662(.A0(men_men_n588_), .A1(men_men_n436_), .B0(men_men_n49_), .Y(men_men_n691_));
  OAI220     u0663(.A0(men_men_n611_), .A1(men_men_n604_), .B0(men_men_n329_), .B1(men_men_n542_), .Y(men_men_n692_));
  AOI210     u0664(.A0(men_men_n692_), .A1(men_men_n691_), .B0(men_men_n690_), .Y(men_men_n693_));
  NA3        u0665(.A(men_men_n693_), .B(men_men_n686_), .C(men_men_n684_), .Y(men_men_n694_));
  NO2        u0666(.A(men_men_n254_), .B(f), .Y(men_men_n695_));
  NO2        u0667(.A(men_men_n636_), .B(men_men_n61_), .Y(men_men_n696_));
  NO3        u0668(.A(men_men_n696_), .B(men_men_n695_), .C(men_men_n34_), .Y(men_men_n697_));
  NA2        u0669(.A(men_men_n332_), .B(men_men_n142_), .Y(men_men_n698_));
  NA2        u0670(.A(men_men_n134_), .B(men_men_n49_), .Y(men_men_n699_));
  AOI220     u0671(.A0(men_men_n699_), .A1(men_men_n547_), .B0(men_men_n367_), .B1(men_men_n114_), .Y(men_men_n700_));
  OA220      u0672(.A0(men_men_n700_), .A1(men_men_n569_), .B0(men_men_n365_), .B1(men_men_n112_), .Y(men_men_n701_));
  OAI210     u0673(.A0(men_men_n698_), .A1(men_men_n697_), .B0(men_men_n701_), .Y(men_men_n702_));
  NO3        u0674(.A(men_men_n411_), .B(men_men_n195_), .C(men_men_n194_), .Y(men_men_n703_));
  NA2        u0675(.A(men_men_n703_), .B(men_men_n235_), .Y(men_men_n704_));
  NA3        u0676(.A(men_men_n704_), .B(men_men_n256_), .C(j), .Y(men_men_n705_));
  NO3        u0677(.A(men_men_n472_), .B(men_men_n175_), .C(i), .Y(men_men_n706_));
  NA2        u0678(.A(men_men_n476_), .B(men_men_n86_), .Y(men_men_n707_));
  NO4        u0679(.A(men_men_n544_), .B(men_men_n707_), .C(men_men_n133_), .D(men_men_n217_), .Y(men_men_n708_));
  INV        u0680(.A(men_men_n708_), .Y(men_men_n709_));
  NA4        u0681(.A(men_men_n709_), .B(men_men_n705_), .C(men_men_n529_), .D(men_men_n409_), .Y(men_men_n710_));
  NO4        u0682(.A(men_men_n710_), .B(men_men_n702_), .C(men_men_n694_), .D(men_men_n680_), .Y(men_men_n711_));
  NA4        u0683(.A(men_men_n711_), .B(men_men_n672_), .C(men_men_n625_), .D(men_men_n602_), .Y(men08));
  NO2        u0684(.A(k), .B(h), .Y(men_men_n713_));
  AO210      u0685(.A0(men_men_n254_), .A1(men_men_n461_), .B0(men_men_n713_), .Y(men_men_n714_));
  NO2        u0686(.A(men_men_n714_), .B(men_men_n299_), .Y(men_men_n715_));
  NA2        u0687(.A(men_men_n635_), .B(men_men_n86_), .Y(men_men_n716_));
  NA2        u0688(.A(men_men_n716_), .B(men_men_n472_), .Y(men_men_n717_));
  AOI210     u0689(.A0(men_men_n717_), .A1(men_men_n715_), .B0(men_men_n507_), .Y(men_men_n718_));
  NA2        u0690(.A(men_men_n86_), .B(men_men_n111_), .Y(men_men_n719_));
  NO2        u0691(.A(men_men_n719_), .B(men_men_n57_), .Y(men_men_n720_));
  NO4        u0692(.A(men_men_n385_), .B(men_men_n113_), .C(j), .D(men_men_n218_), .Y(men_men_n721_));
  NA2        u0693(.A(men_men_n598_), .B(men_men_n237_), .Y(men_men_n722_));
  AOI220     u0694(.A0(men_men_n722_), .A1(men_men_n352_), .B0(men_men_n721_), .B1(men_men_n720_), .Y(men_men_n723_));
  AOI210     u0695(.A0(men_men_n598_), .A1(men_men_n157_), .B0(men_men_n86_), .Y(men_men_n724_));
  NA4        u0696(.A(men_men_n220_), .B(men_men_n142_), .C(men_men_n45_), .D(h), .Y(men_men_n725_));
  AN2        u0697(.A(l), .B(k), .Y(men_men_n726_));
  NA4        u0698(.A(men_men_n726_), .B(men_men_n109_), .C(men_men_n75_), .D(men_men_n218_), .Y(men_men_n727_));
  OAI210     u0699(.A0(men_men_n725_), .A1(u), .B0(men_men_n727_), .Y(men_men_n728_));
  NA2        u0700(.A(men_men_n728_), .B(men_men_n724_), .Y(men_men_n729_));
  NA4        u0701(.A(men_men_n729_), .B(men_men_n723_), .C(men_men_n718_), .D(men_men_n354_), .Y(men_men_n730_));
  NO4        u0702(.A(men_men_n175_), .B(men_men_n399_), .C(men_men_n113_), .D(u), .Y(men_men_n731_));
  AOI210     u0703(.A0(men_men_n731_), .A1(men_men_n722_), .B0(men_men_n536_), .Y(men_men_n732_));
  NO2        u0704(.A(men_men_n38_), .B(men_men_n217_), .Y(men_men_n733_));
  AOI220     u0705(.A0(men_men_n637_), .A1(men_men_n351_), .B0(men_men_n733_), .B1(men_men_n585_), .Y(men_men_n734_));
  NA2        u0706(.A(men_men_n734_), .B(men_men_n732_), .Y(men_men_n735_));
  OAI210     u0707(.A0(men_men_n572_), .A1(men_men_n47_), .B0(men_men_n668_), .Y(men_men_n736_));
  NO2        u0708(.A(men_men_n499_), .B(men_men_n134_), .Y(men_men_n737_));
  NA2        u0709(.A(men_men_n737_), .B(men_men_n736_), .Y(men_men_n738_));
  NO3        u0710(.A(men_men_n320_), .B(men_men_n133_), .C(men_men_n41_), .Y(men_men_n739_));
  NAi21      u0711(.An(men_men_n739_), .B(men_men_n727_), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n714_), .B(men_men_n138_), .Y(men_men_n741_));
  AOI220     u0713(.A0(men_men_n741_), .A1(men_men_n410_), .B0(men_men_n740_), .B1(men_men_n78_), .Y(men_men_n742_));
  NA2        u0714(.A(men_men_n738_), .B(men_men_n742_), .Y(men_men_n743_));
  NA2        u0715(.A(men_men_n367_), .B(men_men_n43_), .Y(men_men_n744_));
  NA3        u0716(.A(men_men_n704_), .B(men_men_n338_), .C(men_men_n391_), .Y(men_men_n745_));
  NA2        u0717(.A(men_men_n726_), .B(men_men_n225_), .Y(men_men_n746_));
  NO2        u0718(.A(men_men_n746_), .B(men_men_n331_), .Y(men_men_n747_));
  AOI210     u0719(.A0(men_men_n747_), .A1(men_men_n695_), .B0(men_men_n506_), .Y(men_men_n748_));
  NA3        u0720(.A(m), .B(l), .C(k), .Y(men_men_n749_));
  AOI210     u0721(.A0(men_men_n677_), .A1(men_men_n675_), .B0(men_men_n749_), .Y(men_men_n750_));
  NO2        u0722(.A(men_men_n554_), .B(men_men_n275_), .Y(men_men_n751_));
  NOi21      u0723(.An(men_men_n751_), .B(men_men_n548_), .Y(men_men_n752_));
  NA4        u0724(.A(men_men_n114_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n753_));
  NA3        u0725(.A(men_men_n122_), .B(men_men_n419_), .C(i), .Y(men_men_n754_));
  NO2        u0726(.A(men_men_n754_), .B(men_men_n753_), .Y(men_men_n755_));
  NO3        u0727(.A(men_men_n755_), .B(men_men_n752_), .C(men_men_n750_), .Y(men_men_n756_));
  NA4        u0728(.A(men_men_n756_), .B(men_men_n748_), .C(men_men_n745_), .D(men_men_n744_), .Y(men_men_n757_));
  NO4        u0729(.A(men_men_n757_), .B(men_men_n743_), .C(men_men_n735_), .D(men_men_n730_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n637_), .B(men_men_n400_), .Y(men_men_n759_));
  NOi31      u0731(.An(u), .B(h), .C(f), .Y(men_men_n760_));
  NA2        u0732(.A(men_men_n650_), .B(men_men_n760_), .Y(men_men_n761_));
  AO210      u0733(.A0(men_men_n761_), .A1(men_men_n612_), .B0(men_men_n557_), .Y(men_men_n762_));
  NO3        u0734(.A(men_men_n404_), .B(men_men_n542_), .C(h), .Y(men_men_n763_));
  AOI210     u0735(.A0(men_men_n763_), .A1(men_men_n114_), .B0(men_men_n515_), .Y(men_men_n764_));
  NA4        u0736(.A(men_men_n764_), .B(men_men_n762_), .C(men_men_n759_), .D(men_men_n253_), .Y(men_men_n765_));
  NA2        u0737(.A(men_men_n726_), .B(men_men_n75_), .Y(men_men_n766_));
  NO4        u0738(.A(men_men_n703_), .B(men_men_n175_), .C(n), .D(i), .Y(men_men_n767_));
  NOi21      u0739(.An(h), .B(j), .Y(men_men_n768_));
  NA2        u0740(.A(men_men_n768_), .B(f), .Y(men_men_n769_));
  NO2        u0741(.A(men_men_n767_), .B(men_men_n706_), .Y(men_men_n770_));
  OAI220     u0742(.A0(men_men_n770_), .A1(men_men_n766_), .B0(men_men_n614_), .B1(men_men_n62_), .Y(men_men_n771_));
  AOI210     u0743(.A0(men_men_n765_), .A1(l), .B0(men_men_n771_), .Y(men_men_n772_));
  NO2        u0744(.A(j), .B(i), .Y(men_men_n773_));
  NA3        u0745(.A(men_men_n773_), .B(men_men_n82_), .C(l), .Y(men_men_n774_));
  NA2        u0746(.A(men_men_n773_), .B(men_men_n33_), .Y(men_men_n775_));
  NA2        u0747(.A(men_men_n429_), .B(men_men_n122_), .Y(men_men_n776_));
  OR2        u0748(.A(men_men_n776_), .B(men_men_n775_), .Y(men_men_n777_));
  NO3        u0749(.A(men_men_n152_), .B(men_men_n49_), .C(men_men_n111_), .Y(men_men_n778_));
  NO3        u0750(.A(men_men_n561_), .B(men_men_n150_), .C(men_men_n75_), .Y(men_men_n779_));
  NO3        u0751(.A(men_men_n499_), .B(men_men_n448_), .C(j), .Y(men_men_n780_));
  OAI210     u0752(.A0(men_men_n779_), .A1(men_men_n778_), .B0(men_men_n780_), .Y(men_men_n781_));
  OAI210     u0753(.A0(men_men_n761_), .A1(men_men_n62_), .B0(men_men_n781_), .Y(men_men_n782_));
  NA2        u0754(.A(k), .B(j), .Y(men_men_n783_));
  NO3        u0755(.A(men_men_n299_), .B(men_men_n783_), .C(men_men_n40_), .Y(men_men_n784_));
  AOI210     u0756(.A0(men_men_n547_), .A1(n), .B0(men_men_n571_), .Y(men_men_n785_));
  NA2        u0757(.A(men_men_n785_), .B(men_men_n574_), .Y(men_men_n786_));
  AN3        u0758(.A(men_men_n786_), .B(men_men_n784_), .C(men_men_n99_), .Y(men_men_n787_));
  NA2        u0759(.A(men_men_n628_), .B(men_men_n310_), .Y(men_men_n788_));
  INV        u0760(.A(men_men_n788_), .Y(men_men_n789_));
  NO2        u0761(.A(men_men_n299_), .B(men_men_n138_), .Y(men_men_n790_));
  AOI220     u0762(.A0(men_men_n790_), .A1(men_men_n637_), .B0(men_men_n739_), .B1(men_men_n724_), .Y(men_men_n791_));
  NO2        u0763(.A(men_men_n749_), .B(men_men_n92_), .Y(men_men_n792_));
  NA2        u0764(.A(men_men_n792_), .B(men_men_n609_), .Y(men_men_n793_));
  NO2        u0765(.A(men_men_n611_), .B(men_men_n118_), .Y(men_men_n794_));
  OAI210     u0766(.A0(men_men_n794_), .A1(men_men_n780_), .B0(men_men_n691_), .Y(men_men_n795_));
  NA3        u0767(.A(men_men_n795_), .B(men_men_n793_), .C(men_men_n791_), .Y(men_men_n796_));
  OR4        u0768(.A(men_men_n796_), .B(men_men_n789_), .C(men_men_n787_), .D(men_men_n782_), .Y(men_men_n797_));
  NA3        u0769(.A(men_men_n785_), .B(men_men_n574_), .C(men_men_n573_), .Y(men_men_n798_));
  NA4        u0770(.A(men_men_n798_), .B(men_men_n220_), .C(men_men_n461_), .D(men_men_n34_), .Y(men_men_n799_));
  NO4        u0771(.A(men_men_n499_), .B(men_men_n443_), .C(j), .D(f), .Y(men_men_n800_));
  OAI220     u0772(.A0(men_men_n725_), .A1(men_men_n716_), .B0(men_men_n336_), .B1(men_men_n38_), .Y(men_men_n801_));
  AOI210     u0773(.A0(men_men_n800_), .A1(men_men_n260_), .B0(men_men_n801_), .Y(men_men_n802_));
  NA3        u0774(.A(men_men_n564_), .B(men_men_n296_), .C(h), .Y(men_men_n803_));
  NOi21      u0775(.An(men_men_n691_), .B(men_men_n803_), .Y(men_men_n804_));
  NO2        u0776(.A(men_men_n93_), .B(men_men_n47_), .Y(men_men_n805_));
  OAI220     u0777(.A0(men_men_n803_), .A1(men_men_n622_), .B0(men_men_n774_), .B1(men_men_n685_), .Y(men_men_n806_));
  AOI210     u0778(.A0(men_men_n805_), .A1(men_men_n656_), .B0(men_men_n806_), .Y(men_men_n807_));
  NAi41      u0779(.An(men_men_n804_), .B(men_men_n807_), .C(men_men_n802_), .D(men_men_n799_), .Y(men_men_n808_));
  OR2        u0780(.A(men_men_n792_), .B(men_men_n96_), .Y(men_men_n809_));
  AOI220     u0781(.A0(men_men_n809_), .A1(men_men_n242_), .B0(men_men_n780_), .B1(men_men_n649_), .Y(men_men_n810_));
  INV        u0782(.A(men_men_n340_), .Y(men_men_n811_));
  OAI210     u0783(.A0(men_men_n749_), .A1(men_men_n674_), .B0(men_men_n535_), .Y(men_men_n812_));
  NA3        u0784(.A(men_men_n252_), .B(men_men_n59_), .C(b), .Y(men_men_n813_));
  AOI220     u0785(.A0(men_men_n621_), .A1(men_men_n29_), .B0(men_men_n476_), .B1(men_men_n86_), .Y(men_men_n814_));
  NA2        u0786(.A(men_men_n814_), .B(men_men_n813_), .Y(men_men_n815_));
  NO2        u0787(.A(men_men_n803_), .B(men_men_n505_), .Y(men_men_n816_));
  AOI210     u0788(.A0(men_men_n815_), .A1(men_men_n812_), .B0(men_men_n816_), .Y(men_men_n817_));
  NA3        u0789(.A(men_men_n817_), .B(men_men_n811_), .C(men_men_n810_), .Y(men_men_n818_));
  NOi41      u0790(.An(men_men_n777_), .B(men_men_n818_), .C(men_men_n808_), .D(men_men_n797_), .Y(men_men_n819_));
  NO3        u0791(.A(men_men_n346_), .B(men_men_n301_), .C(men_men_n113_), .Y(men_men_n820_));
  NA2        u0792(.A(men_men_n820_), .B(men_men_n786_), .Y(men_men_n821_));
  NA2        u0793(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n822_));
  NO3        u0794(.A(men_men_n822_), .B(men_men_n775_), .C(men_men_n280_), .Y(men_men_n823_));
  NO3        u0795(.A(men_men_n542_), .B(men_men_n94_), .C(h), .Y(men_men_n824_));
  AOI210     u0796(.A0(men_men_n824_), .A1(men_men_n720_), .B0(men_men_n823_), .Y(men_men_n825_));
  NA3        u0797(.A(men_men_n825_), .B(men_men_n821_), .C(men_men_n412_), .Y(men_men_n826_));
  OR2        u0798(.A(men_men_n674_), .B(men_men_n93_), .Y(men_men_n827_));
  NOi31      u0799(.An(b), .B(d), .C(a), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n828_), .B(men_men_n620_), .Y(men_men_n829_));
  NO2        u0801(.A(men_men_n829_), .B(n), .Y(men_men_n830_));
  NOi21      u0802(.An(men_men_n814_), .B(men_men_n830_), .Y(men_men_n831_));
  NO2        u0803(.A(men_men_n831_), .B(men_men_n827_), .Y(men_men_n832_));
  NO2        u0804(.A(men_men_n572_), .B(men_men_n86_), .Y(men_men_n833_));
  NA2        u0805(.A(men_men_n820_), .B(men_men_n833_), .Y(men_men_n834_));
  OAI210     u0806(.A0(men_men_n725_), .A1(men_men_n401_), .B0(men_men_n834_), .Y(men_men_n835_));
  NO2        u0807(.A(men_men_n703_), .B(n), .Y(men_men_n836_));
  AOI220     u0808(.A0(men_men_n790_), .A1(men_men_n681_), .B0(men_men_n836_), .B1(men_men_n715_), .Y(men_men_n837_));
  NO2        u0809(.A(men_men_n326_), .B(men_men_n241_), .Y(men_men_n838_));
  NA2        u0810(.A(men_men_n122_), .B(men_men_n86_), .Y(men_men_n839_));
  AOI210     u0811(.A0(men_men_n433_), .A1(men_men_n425_), .B0(men_men_n839_), .Y(men_men_n840_));
  NA2        u0812(.A(men_men_n747_), .B(men_men_n34_), .Y(men_men_n841_));
  NAi21      u0813(.An(men_men_n753_), .B(men_men_n444_), .Y(men_men_n842_));
  NO2        u0814(.A(men_men_n275_), .B(i), .Y(men_men_n843_));
  NA2        u0815(.A(men_men_n731_), .B(men_men_n353_), .Y(men_men_n844_));
  AN2        u0816(.A(men_men_n844_), .B(men_men_n842_), .Y(men_men_n845_));
  NAi41      u0817(.An(men_men_n840_), .B(men_men_n845_), .C(men_men_n841_), .D(men_men_n837_), .Y(men_men_n846_));
  NO4        u0818(.A(men_men_n846_), .B(men_men_n835_), .C(men_men_n832_), .D(men_men_n826_), .Y(men_men_n847_));
  NA4        u0819(.A(men_men_n847_), .B(men_men_n819_), .C(men_men_n772_), .D(men_men_n758_), .Y(men09));
  INV        u0820(.A(men_men_n123_), .Y(men_men_n849_));
  NA2        u0821(.A(f), .B(e), .Y(men_men_n850_));
  NO2        u0822(.A(men_men_n230_), .B(men_men_n113_), .Y(men_men_n851_));
  NA2        u0823(.A(men_men_n851_), .B(u), .Y(men_men_n852_));
  NA4        u0824(.A(men_men_n313_), .B(men_men_n485_), .C(men_men_n263_), .D(men_men_n120_), .Y(men_men_n853_));
  AOI210     u0825(.A0(men_men_n853_), .A1(u), .B0(men_men_n482_), .Y(men_men_n854_));
  AOI210     u0826(.A0(men_men_n854_), .A1(men_men_n852_), .B0(men_men_n850_), .Y(men_men_n855_));
  NA2        u0827(.A(men_men_n454_), .B(e), .Y(men_men_n856_));
  NO2        u0828(.A(men_men_n856_), .B(men_men_n526_), .Y(men_men_n857_));
  AOI210     u0829(.A0(men_men_n855_), .A1(men_men_n849_), .B0(men_men_n857_), .Y(men_men_n858_));
  NO2        u0830(.A(men_men_n207_), .B(men_men_n217_), .Y(men_men_n859_));
  NA3        u0831(.A(m), .B(l), .C(i), .Y(men_men_n860_));
  OAI220     u0832(.A0(men_men_n611_), .A1(men_men_n860_), .B0(men_men_n358_), .B1(men_men_n543_), .Y(men_men_n861_));
  NA4        u0833(.A(men_men_n90_), .B(men_men_n89_), .C(u), .D(f), .Y(men_men_n862_));
  NAi31      u0834(.An(men_men_n861_), .B(men_men_n862_), .C(men_men_n449_), .Y(men_men_n863_));
  OR2        u0835(.A(men_men_n863_), .B(men_men_n859_), .Y(men_men_n864_));
  NA3        u0836(.A(men_men_n827_), .B(men_men_n587_), .C(men_men_n535_), .Y(men_men_n865_));
  OA210      u0837(.A0(men_men_n865_), .A1(men_men_n864_), .B0(men_men_n830_), .Y(men_men_n866_));
  INV        u0838(.A(men_men_n343_), .Y(men_men_n867_));
  NO2        u0839(.A(men_men_n129_), .B(men_men_n127_), .Y(men_men_n868_));
  NOi31      u0840(.An(k), .B(m), .C(l), .Y(men_men_n869_));
  NO2        u0841(.A(men_men_n345_), .B(men_men_n869_), .Y(men_men_n870_));
  AOI210     u0842(.A0(men_men_n870_), .A1(men_men_n868_), .B0(men_men_n617_), .Y(men_men_n871_));
  NA2        u0843(.A(men_men_n813_), .B(men_men_n336_), .Y(men_men_n872_));
  NA2        u0844(.A(men_men_n347_), .B(men_men_n349_), .Y(men_men_n873_));
  OAI210     u0845(.A0(men_men_n207_), .A1(men_men_n217_), .B0(men_men_n873_), .Y(men_men_n874_));
  AOI220     u0846(.A0(men_men_n874_), .A1(men_men_n872_), .B0(men_men_n871_), .B1(men_men_n867_), .Y(men_men_n875_));
  NA2        u0847(.A(men_men_n169_), .B(men_men_n115_), .Y(men_men_n876_));
  NA3        u0848(.A(men_men_n876_), .B(men_men_n714_), .C(men_men_n138_), .Y(men_men_n877_));
  NA3        u0849(.A(men_men_n877_), .B(men_men_n192_), .C(men_men_n31_), .Y(men_men_n878_));
  NA4        u0850(.A(men_men_n878_), .B(men_men_n875_), .C(men_men_n638_), .D(men_men_n84_), .Y(men_men_n879_));
  NO2        u0851(.A(men_men_n607_), .B(men_men_n512_), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n880_), .B(men_men_n192_), .Y(men_men_n881_));
  NOi21      u0853(.An(f), .B(d), .Y(men_men_n882_));
  NA2        u0854(.A(men_men_n882_), .B(m), .Y(men_men_n883_));
  NO2        u0855(.A(men_men_n883_), .B(men_men_n52_), .Y(men_men_n884_));
  NOi32      u0856(.An(u), .Bn(f), .C(d), .Y(men_men_n885_));
  NA4        u0857(.A(men_men_n885_), .B(men_men_n621_), .C(men_men_n29_), .D(m), .Y(men_men_n886_));
  NA2        u0858(.A(men_men_n884_), .B(men_men_n562_), .Y(men_men_n887_));
  NA3        u0859(.A(men_men_n313_), .B(men_men_n263_), .C(men_men_n120_), .Y(men_men_n888_));
  AN2        u0860(.A(f), .B(d), .Y(men_men_n889_));
  NA3        u0861(.A(men_men_n490_), .B(men_men_n889_), .C(men_men_n86_), .Y(men_men_n890_));
  NO3        u0862(.A(men_men_n890_), .B(men_men_n75_), .C(men_men_n218_), .Y(men_men_n891_));
  NO2        u0863(.A(men_men_n289_), .B(men_men_n56_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n888_), .B(men_men_n891_), .Y(men_men_n893_));
  NAi41      u0865(.An(men_men_n504_), .B(men_men_n893_), .C(men_men_n887_), .D(men_men_n881_), .Y(men_men_n894_));
  NO4        u0866(.A(men_men_n636_), .B(men_men_n134_), .C(men_men_n331_), .D(men_men_n153_), .Y(men_men_n895_));
  NO2        u0867(.A(men_men_n667_), .B(men_men_n331_), .Y(men_men_n896_));
  AN2        u0868(.A(men_men_n896_), .B(men_men_n695_), .Y(men_men_n897_));
  NO2        u0869(.A(men_men_n897_), .B(men_men_n895_), .Y(men_men_n898_));
  NA2        u0870(.A(men_men_n620_), .B(men_men_n86_), .Y(men_men_n899_));
  NA3        u0871(.A(men_men_n161_), .B(men_men_n109_), .C(men_men_n108_), .Y(men_men_n900_));
  OAI220     u0872(.A0(men_men_n890_), .A1(men_men_n438_), .B0(men_men_n343_), .B1(men_men_n900_), .Y(men_men_n901_));
  NOi31      u0873(.An(men_men_n228_), .B(men_men_n901_), .C(men_men_n308_), .Y(men_men_n902_));
  NA2        u0874(.A(c), .B(men_men_n117_), .Y(men_men_n903_));
  NO2        u0875(.A(men_men_n903_), .B(men_men_n416_), .Y(men_men_n904_));
  NA3        u0876(.A(men_men_n904_), .B(men_men_n524_), .C(f), .Y(men_men_n905_));
  OR2        u0877(.A(men_men_n674_), .B(men_men_n558_), .Y(men_men_n906_));
  INV        u0878(.A(men_men_n906_), .Y(men_men_n907_));
  NA2        u0879(.A(men_men_n829_), .B(men_men_n112_), .Y(men_men_n908_));
  NA2        u0880(.A(men_men_n908_), .B(men_men_n907_), .Y(men_men_n909_));
  NA4        u0881(.A(men_men_n909_), .B(men_men_n905_), .C(men_men_n902_), .D(men_men_n898_), .Y(men_men_n910_));
  NO4        u0882(.A(men_men_n910_), .B(men_men_n894_), .C(men_men_n879_), .D(men_men_n866_), .Y(men_men_n911_));
  OR2        u0883(.A(men_men_n890_), .B(men_men_n75_), .Y(men_men_n912_));
  NA2        u0884(.A(men_men_n113_), .B(j), .Y(men_men_n913_));
  NA2        u0885(.A(men_men_n851_), .B(u), .Y(men_men_n914_));
  AOI210     u0886(.A0(men_men_n914_), .A1(men_men_n297_), .B0(men_men_n912_), .Y(men_men_n915_));
  NO2        u0887(.A(men_men_n336_), .B(men_men_n862_), .Y(men_men_n916_));
  NO2        u0888(.A(men_men_n138_), .B(men_men_n134_), .Y(men_men_n917_));
  NO2        u0889(.A(men_men_n235_), .B(men_men_n229_), .Y(men_men_n918_));
  AOI220     u0890(.A0(men_men_n918_), .A1(men_men_n232_), .B0(men_men_n306_), .B1(men_men_n917_), .Y(men_men_n919_));
  NO2        u0891(.A(men_men_n438_), .B(men_men_n850_), .Y(men_men_n920_));
  NA2        u0892(.A(men_men_n920_), .B(men_men_n579_), .Y(men_men_n921_));
  NA2        u0893(.A(men_men_n921_), .B(men_men_n919_), .Y(men_men_n922_));
  NA2        u0894(.A(e), .B(d), .Y(men_men_n923_));
  OAI220     u0895(.A0(men_men_n923_), .A1(c), .B0(men_men_n326_), .B1(d), .Y(men_men_n924_));
  NA3        u0896(.A(men_men_n924_), .B(men_men_n465_), .C(men_men_n522_), .Y(men_men_n925_));
  AOI210     u0897(.A0(men_men_n530_), .A1(men_men_n182_), .B0(men_men_n235_), .Y(men_men_n926_));
  AOI210     u0898(.A0(men_men_n637_), .A1(men_men_n351_), .B0(men_men_n926_), .Y(men_men_n927_));
  NA2        u0899(.A(men_men_n289_), .B(men_men_n167_), .Y(men_men_n928_));
  NA2        u0900(.A(men_men_n891_), .B(men_men_n928_), .Y(men_men_n929_));
  NA3        u0901(.A(men_men_n168_), .B(men_men_n87_), .C(men_men_n34_), .Y(men_men_n930_));
  NA4        u0902(.A(men_men_n930_), .B(men_men_n929_), .C(men_men_n927_), .D(men_men_n925_), .Y(men_men_n931_));
  NO4        u0903(.A(men_men_n931_), .B(men_men_n922_), .C(men_men_n916_), .D(men_men_n915_), .Y(men_men_n932_));
  NA2        u0904(.A(men_men_n867_), .B(men_men_n31_), .Y(men_men_n933_));
  AO210      u0905(.A0(men_men_n933_), .A1(men_men_n716_), .B0(men_men_n221_), .Y(men_men_n934_));
  OAI220     u0906(.A0(men_men_n636_), .A1(men_men_n61_), .B0(men_men_n301_), .B1(j), .Y(men_men_n935_));
  AOI220     u0907(.A0(men_men_n935_), .A1(men_men_n896_), .B0(men_men_n626_), .B1(men_men_n635_), .Y(men_men_n936_));
  OAI210     u0908(.A0(men_men_n856_), .A1(men_men_n172_), .B0(men_men_n936_), .Y(men_men_n937_));
  OAI210     u0909(.A0(men_men_n851_), .A1(men_men_n928_), .B0(men_men_n885_), .Y(men_men_n938_));
  NO2        u0910(.A(men_men_n938_), .B(men_men_n622_), .Y(men_men_n939_));
  AOI210     u0911(.A0(men_men_n119_), .A1(men_men_n118_), .B0(men_men_n262_), .Y(men_men_n940_));
  NO2        u0912(.A(men_men_n940_), .B(men_men_n886_), .Y(men_men_n941_));
  AO210      u0913(.A0(men_men_n872_), .A1(men_men_n861_), .B0(men_men_n941_), .Y(men_men_n942_));
  NOi31      u0914(.An(men_men_n562_), .B(men_men_n883_), .C(men_men_n297_), .Y(men_men_n943_));
  NO4        u0915(.A(men_men_n943_), .B(men_men_n942_), .C(men_men_n939_), .D(men_men_n937_), .Y(men_men_n944_));
  AO220      u0916(.A0(men_men_n465_), .A1(men_men_n768_), .B0(men_men_n177_), .B1(f), .Y(men_men_n945_));
  OAI210     u0917(.A0(men_men_n945_), .A1(men_men_n468_), .B0(men_men_n924_), .Y(men_men_n946_));
  NO2        u0918(.A(men_men_n448_), .B(men_men_n71_), .Y(men_men_n947_));
  OAI210     u0919(.A0(men_men_n865_), .A1(men_men_n947_), .B0(men_men_n720_), .Y(men_men_n948_));
  AN4        u0920(.A(men_men_n948_), .B(men_men_n946_), .C(men_men_n944_), .D(men_men_n934_), .Y(men_men_n949_));
  NA4        u0921(.A(men_men_n949_), .B(men_men_n932_), .C(men_men_n911_), .D(men_men_n858_), .Y(men12));
  NO2        u0922(.A(men_men_n463_), .B(c), .Y(men_men_n951_));
  NO4        u0923(.A(men_men_n453_), .B(men_men_n254_), .C(men_men_n603_), .D(men_men_n218_), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n952_), .B(men_men_n951_), .Y(men_men_n953_));
  NA2        u0925(.A(men_men_n562_), .B(men_men_n947_), .Y(men_men_n954_));
  NO2        u0926(.A(men_men_n463_), .B(men_men_n117_), .Y(men_men_n955_));
  NO2        u0927(.A(men_men_n868_), .B(men_men_n358_), .Y(men_men_n956_));
  NO2        u0928(.A(men_men_n674_), .B(men_men_n385_), .Y(men_men_n957_));
  AOI220     u0929(.A0(men_men_n957_), .A1(men_men_n560_), .B0(men_men_n956_), .B1(men_men_n955_), .Y(men_men_n958_));
  NA4        u0930(.A(men_men_n958_), .B(men_men_n954_), .C(men_men_n953_), .D(men_men_n452_), .Y(men_men_n959_));
  AOI210     u0931(.A0(men_men_n238_), .A1(men_men_n342_), .B0(men_men_n204_), .Y(men_men_n960_));
  OR2        u0932(.A(men_men_n960_), .B(men_men_n952_), .Y(men_men_n961_));
  AOI210     u0933(.A0(men_men_n339_), .A1(men_men_n397_), .B0(men_men_n218_), .Y(men_men_n962_));
  OAI210     u0934(.A0(men_men_n962_), .A1(men_men_n961_), .B0(men_men_n411_), .Y(men_men_n963_));
  NO2        u0935(.A(men_men_n653_), .B(men_men_n265_), .Y(men_men_n964_));
  NO2        u0936(.A(men_men_n611_), .B(men_men_n860_), .Y(men_men_n965_));
  AOI220     u0937(.A0(men_men_n965_), .A1(men_men_n585_), .B0(men_men_n838_), .B1(men_men_n964_), .Y(men_men_n966_));
  NO2        u0938(.A(men_men_n152_), .B(men_men_n241_), .Y(men_men_n967_));
  NA3        u0939(.A(men_men_n967_), .B(men_men_n244_), .C(i), .Y(men_men_n968_));
  NA3        u0940(.A(men_men_n968_), .B(men_men_n966_), .C(men_men_n963_), .Y(men_men_n969_));
  OR2        u0941(.A(men_men_n327_), .B(men_men_n955_), .Y(men_men_n970_));
  NA2        u0942(.A(men_men_n970_), .B(men_men_n359_), .Y(men_men_n971_));
  NO3        u0943(.A(men_men_n134_), .B(men_men_n153_), .C(men_men_n218_), .Y(men_men_n972_));
  NA2        u0944(.A(men_men_n972_), .B(men_men_n547_), .Y(men_men_n973_));
  NA4        u0945(.A(men_men_n454_), .B(men_men_n446_), .C(men_men_n183_), .D(u), .Y(men_men_n974_));
  NA3        u0946(.A(men_men_n974_), .B(men_men_n973_), .C(men_men_n971_), .Y(men_men_n975_));
  NO3        u0947(.A(men_men_n679_), .B(men_men_n93_), .C(men_men_n45_), .Y(men_men_n976_));
  NO4        u0948(.A(men_men_n976_), .B(men_men_n975_), .C(men_men_n969_), .D(men_men_n959_), .Y(men_men_n977_));
  NO2        u0949(.A(men_men_n375_), .B(men_men_n374_), .Y(men_men_n978_));
  NA2        u0950(.A(men_men_n608_), .B(men_men_n73_), .Y(men_men_n979_));
  NA2        u0951(.A(men_men_n572_), .B(men_men_n146_), .Y(men_men_n980_));
  NOi21      u0952(.An(men_men_n34_), .B(men_men_n667_), .Y(men_men_n981_));
  AOI220     u0953(.A0(men_men_n981_), .A1(men_men_n980_), .B0(men_men_n979_), .B1(men_men_n978_), .Y(men_men_n982_));
  OAI210     u0954(.A0(men_men_n253_), .A1(men_men_n45_), .B0(men_men_n982_), .Y(men_men_n983_));
  NA2        u0955(.A(men_men_n444_), .B(men_men_n267_), .Y(men_men_n984_));
  NO3        u0956(.A(men_men_n839_), .B(men_men_n91_), .C(men_men_n416_), .Y(men_men_n985_));
  NAi31      u0957(.An(men_men_n985_), .B(men_men_n984_), .C(men_men_n324_), .Y(men_men_n986_));
  NO2        u0958(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n987_));
  NO2        u0959(.A(men_men_n518_), .B(men_men_n301_), .Y(men_men_n988_));
  INV        u0960(.A(men_men_n988_), .Y(men_men_n989_));
  NO2        u0961(.A(men_men_n989_), .B(men_men_n146_), .Y(men_men_n990_));
  NA2        u0962(.A(men_men_n645_), .B(men_men_n368_), .Y(men_men_n991_));
  OAI210     u0963(.A0(men_men_n754_), .A1(men_men_n991_), .B0(men_men_n372_), .Y(men_men_n992_));
  NO4        u0964(.A(men_men_n992_), .B(men_men_n990_), .C(men_men_n986_), .D(men_men_n983_), .Y(men_men_n993_));
  NA2        u0965(.A(men_men_n351_), .B(u), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n164_), .B(i), .Y(men_men_n995_));
  NA2        u0967(.A(men_men_n46_), .B(i), .Y(men_men_n996_));
  OAI220     u0968(.A0(men_men_n996_), .A1(men_men_n203_), .B0(men_men_n995_), .B1(men_men_n93_), .Y(men_men_n997_));
  AOI210     u0969(.A0(men_men_n427_), .A1(men_men_n37_), .B0(men_men_n997_), .Y(men_men_n998_));
  NO2        u0970(.A(men_men_n146_), .B(men_men_n86_), .Y(men_men_n999_));
  OR2        u0971(.A(men_men_n999_), .B(men_men_n571_), .Y(men_men_n1000_));
  NA2        u0972(.A(men_men_n572_), .B(men_men_n389_), .Y(men_men_n1001_));
  AOI210     u0973(.A0(men_men_n1001_), .A1(n), .B0(men_men_n1000_), .Y(men_men_n1002_));
  OAI220     u0974(.A0(men_men_n1002_), .A1(men_men_n994_), .B0(men_men_n998_), .B1(men_men_n336_), .Y(men_men_n1003_));
  NO2        u0975(.A(men_men_n674_), .B(men_men_n512_), .Y(men_men_n1004_));
  NA3        u0976(.A(men_men_n347_), .B(men_men_n642_), .C(i), .Y(men_men_n1005_));
  OAI210     u0977(.A0(men_men_n448_), .A1(men_men_n313_), .B0(men_men_n1005_), .Y(men_men_n1006_));
  OAI220     u0978(.A0(men_men_n1006_), .A1(men_men_n1004_), .B0(men_men_n691_), .B1(men_men_n779_), .Y(men_men_n1007_));
  OR3        u0979(.A(men_men_n313_), .B(men_men_n443_), .C(f), .Y(men_men_n1008_));
  NA3        u0980(.A(men_men_n328_), .B(men_men_n119_), .C(u), .Y(men_men_n1009_));
  AOI210     u0981(.A0(men_men_n688_), .A1(men_men_n1009_), .B0(m), .Y(men_men_n1010_));
  OAI210     u0982(.A0(men_men_n1010_), .A1(men_men_n956_), .B0(men_men_n327_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n707_), .B(men_men_n899_), .Y(men_men_n1012_));
  NA2        u0984(.A(men_men_n862_), .B(men_men_n449_), .Y(men_men_n1013_));
  INV        u0985(.A(men_men_n1008_), .Y(men_men_n1014_));
  AOI220     u0986(.A0(men_men_n1014_), .A1(men_men_n260_), .B0(men_men_n1013_), .B1(men_men_n1012_), .Y(men_men_n1015_));
  NA3        u0987(.A(men_men_n1015_), .B(men_men_n1011_), .C(men_men_n1007_), .Y(men_men_n1016_));
  NO2        u0988(.A(men_men_n385_), .B(men_men_n92_), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n1017_), .B(men_men_n242_), .Y(men_men_n1018_));
  NA2        u0990(.A(men_men_n678_), .B(men_men_n90_), .Y(men_men_n1019_));
  NO2        u0991(.A(men_men_n471_), .B(men_men_n218_), .Y(men_men_n1020_));
  AOI220     u0992(.A0(men_men_n1020_), .A1(men_men_n390_), .B0(men_men_n970_), .B1(men_men_n222_), .Y(men_men_n1021_));
  NA3        u0993(.A(men_men_n1021_), .B(men_men_n1019_), .C(men_men_n1018_), .Y(men_men_n1022_));
  OAI210     u0994(.A0(men_men_n1013_), .A1(men_men_n965_), .B0(men_men_n560_), .Y(men_men_n1023_));
  OAI210     u0995(.A0(men_men_n375_), .A1(men_men_n374_), .B0(men_men_n110_), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n1024_), .B(men_men_n552_), .Y(men_men_n1025_));
  NA2        u0997(.A(men_men_n1010_), .B(men_men_n955_), .Y(men_men_n1026_));
  NO3        u0998(.A(men_men_n913_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1027_));
  AOI220     u0999(.A0(men_men_n1027_), .A1(men_men_n640_), .B0(men_men_n658_), .B1(men_men_n547_), .Y(men_men_n1028_));
  NA4        u1000(.A(men_men_n1028_), .B(men_men_n1026_), .C(men_men_n1025_), .D(men_men_n1023_), .Y(men_men_n1029_));
  NO4        u1001(.A(men_men_n1029_), .B(men_men_n1022_), .C(men_men_n1016_), .D(men_men_n1003_), .Y(men_men_n1030_));
  NAi31      u1002(.An(men_men_n143_), .B(men_men_n429_), .C(n), .Y(men_men_n1031_));
  NO3        u1003(.A(men_men_n127_), .B(men_men_n345_), .C(men_men_n869_), .Y(men_men_n1032_));
  NO2        u1004(.A(men_men_n1032_), .B(men_men_n1031_), .Y(men_men_n1033_));
  NO3        u1005(.A(men_men_n275_), .B(men_men_n143_), .C(men_men_n416_), .Y(men_men_n1034_));
  AOI210     u1006(.A0(men_men_n1034_), .A1(men_men_n513_), .B0(men_men_n1033_), .Y(men_men_n1035_));
  NA2        u1007(.A(men_men_n507_), .B(i), .Y(men_men_n1036_));
  NA2        u1008(.A(men_men_n1036_), .B(men_men_n1035_), .Y(men_men_n1037_));
  NA2        u1009(.A(men_men_n235_), .B(men_men_n173_), .Y(men_men_n1038_));
  NO3        u1010(.A(men_men_n310_), .B(men_men_n454_), .C(men_men_n177_), .Y(men_men_n1039_));
  NOi31      u1011(.An(men_men_n1038_), .B(men_men_n1039_), .C(men_men_n218_), .Y(men_men_n1040_));
  NAi21      u1012(.An(men_men_n572_), .B(men_men_n1020_), .Y(men_men_n1041_));
  NA2        u1013(.A(men_men_n447_), .B(men_men_n899_), .Y(men_men_n1042_));
  NO3        u1014(.A(men_men_n448_), .B(men_men_n313_), .C(men_men_n75_), .Y(men_men_n1043_));
  AOI220     u1015(.A0(men_men_n1043_), .A1(men_men_n1042_), .B0(men_men_n496_), .B1(u), .Y(men_men_n1044_));
  NA2        u1016(.A(men_men_n1044_), .B(men_men_n1041_), .Y(men_men_n1045_));
  NO2        u1017(.A(men_men_n675_), .B(men_men_n385_), .Y(men_men_n1046_));
  NA2        u1018(.A(men_men_n960_), .B(men_men_n951_), .Y(men_men_n1047_));
  NO3        u1019(.A(men_men_n561_), .B(men_men_n150_), .C(men_men_n217_), .Y(men_men_n1048_));
  OAI210     u1020(.A0(men_men_n1048_), .A1(men_men_n541_), .B0(men_men_n386_), .Y(men_men_n1049_));
  OAI220     u1021(.A0(men_men_n957_), .A1(men_men_n965_), .B0(men_men_n562_), .B1(men_men_n437_), .Y(men_men_n1050_));
  NA4        u1022(.A(men_men_n1050_), .B(men_men_n1049_), .C(men_men_n1047_), .D(men_men_n634_), .Y(men_men_n1051_));
  OAI210     u1023(.A0(men_men_n960_), .A1(men_men_n952_), .B0(men_men_n1038_), .Y(men_men_n1052_));
  NA3        u1024(.A(men_men_n1001_), .B(men_men_n501_), .C(men_men_n46_), .Y(men_men_n1053_));
  INV        u1025(.A(men_men_n335_), .Y(men_men_n1054_));
  NA4        u1026(.A(men_men_n1054_), .B(men_men_n1053_), .C(men_men_n1052_), .D(men_men_n276_), .Y(men_men_n1055_));
  OR3        u1027(.A(men_men_n1055_), .B(men_men_n1051_), .C(men_men_n1046_), .Y(men_men_n1056_));
  NO4        u1028(.A(men_men_n1056_), .B(men_men_n1045_), .C(men_men_n1040_), .D(men_men_n1037_), .Y(men_men_n1057_));
  NA4        u1029(.A(men_men_n1057_), .B(men_men_n1030_), .C(men_men_n993_), .D(men_men_n977_), .Y(men13));
  NA2        u1030(.A(men_men_n46_), .B(men_men_n89_), .Y(men_men_n1059_));
  AN2        u1031(.A(c), .B(b), .Y(men_men_n1060_));
  NA3        u1032(.A(men_men_n252_), .B(men_men_n1060_), .C(m), .Y(men_men_n1061_));
  NA2        u1033(.A(d), .B(f), .Y(men_men_n1062_));
  NO4        u1034(.A(men_men_n1062_), .B(men_men_n1061_), .C(men_men_n1059_), .D(men_men_n604_), .Y(men_men_n1063_));
  NA2        u1035(.A(men_men_n267_), .B(men_men_n1060_), .Y(men_men_n1064_));
  NO4        u1036(.A(men_men_n1064_), .B(men_men_n1062_), .C(men_men_n995_), .D(a), .Y(men_men_n1065_));
  NAi32      u1037(.An(d), .Bn(c), .C(e), .Y(men_men_n1066_));
  NA2        u1038(.A(men_men_n142_), .B(men_men_n45_), .Y(men_men_n1067_));
  NO4        u1039(.A(men_men_n1067_), .B(men_men_n1066_), .C(men_men_n611_), .D(men_men_n309_), .Y(men_men_n1068_));
  NA2        u1040(.A(men_men_n682_), .B(men_men_n229_), .Y(men_men_n1069_));
  NA2        u1041(.A(men_men_n419_), .B(men_men_n217_), .Y(men_men_n1070_));
  AN2        u1042(.A(d), .B(c), .Y(men_men_n1071_));
  NA2        u1043(.A(men_men_n1071_), .B(men_men_n117_), .Y(men_men_n1072_));
  NO4        u1044(.A(men_men_n1072_), .B(men_men_n1070_), .C(men_men_n178_), .D(men_men_n169_), .Y(men_men_n1073_));
  AN2        u1045(.A(men_men_n1073_), .B(men_men_n1069_), .Y(men_men_n1074_));
  OR4        u1046(.A(men_men_n1074_), .B(men_men_n1068_), .C(men_men_n1065_), .D(men_men_n1063_), .Y(men_men_n1075_));
  NAi32      u1047(.An(f), .Bn(e), .C(c), .Y(men_men_n1076_));
  NO2        u1048(.A(men_men_n1076_), .B(men_men_n147_), .Y(men_men_n1077_));
  NA2        u1049(.A(men_men_n1077_), .B(u), .Y(men_men_n1078_));
  OR3        u1050(.A(men_men_n229_), .B(men_men_n178_), .C(men_men_n169_), .Y(men_men_n1079_));
  NO2        u1051(.A(men_men_n1079_), .B(men_men_n1078_), .Y(men_men_n1080_));
  NO2        u1052(.A(j), .B(men_men_n45_), .Y(men_men_n1081_));
  NA2        u1053(.A(men_men_n644_), .B(men_men_n1081_), .Y(men_men_n1082_));
  NO2        u1054(.A(men_men_n783_), .B(men_men_n113_), .Y(men_men_n1083_));
  NOi41      u1055(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1084_));
  NA2        u1056(.A(men_men_n1084_), .B(men_men_n1083_), .Y(men_men_n1085_));
  NO2        u1057(.A(men_men_n1085_), .B(men_men_n1078_), .Y(men_men_n1086_));
  OR3        u1058(.A(e), .B(d), .C(c), .Y(men_men_n1087_));
  NA3        u1059(.A(k), .B(j), .C(i), .Y(men_men_n1088_));
  NO3        u1060(.A(men_men_n1088_), .B(men_men_n309_), .C(men_men_n92_), .Y(men_men_n1089_));
  NOi21      u1061(.An(men_men_n1089_), .B(men_men_n1087_), .Y(men_men_n1090_));
  OR3        u1062(.A(men_men_n1090_), .B(men_men_n1086_), .C(men_men_n1080_), .Y(men_men_n1091_));
  NA3        u1063(.A(men_men_n479_), .B(men_men_n338_), .C(men_men_n56_), .Y(men_men_n1092_));
  NO2        u1064(.A(men_men_n1092_), .B(men_men_n1082_), .Y(men_men_n1093_));
  NO3        u1065(.A(men_men_n1092_), .B(men_men_n607_), .C(men_men_n461_), .Y(men_men_n1094_));
  NO2        u1066(.A(f), .B(c), .Y(men_men_n1095_));
  NOi21      u1067(.An(men_men_n1095_), .B(men_men_n453_), .Y(men_men_n1096_));
  NA2        u1068(.A(men_men_n1096_), .B(men_men_n59_), .Y(men_men_n1097_));
  OR2        u1069(.A(k), .B(i), .Y(men_men_n1098_));
  NO3        u1070(.A(men_men_n1098_), .B(men_men_n248_), .C(l), .Y(men_men_n1099_));
  NOi31      u1071(.An(men_men_n1099_), .B(men_men_n1097_), .C(j), .Y(men_men_n1100_));
  OR3        u1072(.A(men_men_n1100_), .B(men_men_n1094_), .C(men_men_n1093_), .Y(men_men_n1101_));
  OR3        u1073(.A(men_men_n1101_), .B(men_men_n1091_), .C(men_men_n1075_), .Y(men02));
  OR2        u1074(.A(l), .B(k), .Y(men_men_n1103_));
  OR3        u1075(.A(h), .B(u), .C(f), .Y(men_men_n1104_));
  OR3        u1076(.A(n), .B(m), .C(i), .Y(men_men_n1105_));
  NO4        u1077(.A(men_men_n1105_), .B(men_men_n1104_), .C(men_men_n1103_), .D(men_men_n1087_), .Y(men_men_n1106_));
  NOi31      u1078(.An(e), .B(d), .C(c), .Y(men_men_n1107_));
  AOI210     u1079(.A0(men_men_n1089_), .A1(men_men_n1107_), .B0(men_men_n1068_), .Y(men_men_n1108_));
  AN3        u1080(.A(u), .B(f), .C(c), .Y(men_men_n1109_));
  NA2        u1081(.A(men_men_n1109_), .B(men_men_n479_), .Y(men_men_n1110_));
  OR2        u1082(.A(men_men_n1088_), .B(men_men_n309_), .Y(men_men_n1111_));
  OR2        u1083(.A(men_men_n1111_), .B(men_men_n1110_), .Y(men_men_n1112_));
  NO3        u1084(.A(men_men_n1092_), .B(men_men_n1067_), .C(men_men_n607_), .Y(men_men_n1113_));
  NO2        u1085(.A(men_men_n1113_), .B(men_men_n1080_), .Y(men_men_n1114_));
  NA3        u1086(.A(l), .B(k), .C(j), .Y(men_men_n1115_));
  NA2        u1087(.A(i), .B(h), .Y(men_men_n1116_));
  NO3        u1088(.A(men_men_n1116_), .B(men_men_n1115_), .C(men_men_n134_), .Y(men_men_n1117_));
  NO3        u1089(.A(men_men_n144_), .B(men_men_n287_), .C(men_men_n218_), .Y(men_men_n1118_));
  NA2        u1090(.A(men_men_n1118_), .B(men_men_n1117_), .Y(men_men_n1119_));
  NA3        u1091(.A(c), .B(b), .C(a), .Y(men_men_n1120_));
  NO3        u1092(.A(men_men_n1120_), .B(men_men_n923_), .C(men_men_n217_), .Y(men_men_n1121_));
  NO4        u1093(.A(men_men_n1088_), .B(men_men_n301_), .C(men_men_n49_), .D(men_men_n113_), .Y(men_men_n1122_));
  AOI210     u1094(.A0(men_men_n1122_), .A1(men_men_n1121_), .B0(men_men_n1093_), .Y(men_men_n1123_));
  AN4        u1095(.A(men_men_n1123_), .B(men_men_n1119_), .C(men_men_n1114_), .D(men_men_n1112_), .Y(men_men_n1124_));
  NO2        u1096(.A(men_men_n1072_), .B(men_men_n1070_), .Y(men_men_n1125_));
  NA2        u1097(.A(men_men_n1085_), .B(men_men_n1079_), .Y(men_men_n1126_));
  AOI210     u1098(.A0(men_men_n1126_), .A1(men_men_n1125_), .B0(men_men_n1063_), .Y(men_men_n1127_));
  NAi41      u1099(.An(men_men_n1106_), .B(men_men_n1127_), .C(men_men_n1124_), .D(men_men_n1108_), .Y(men03));
  INV        u1100(.A(men_men_n376_), .Y(men_men_n1129_));
  NO2        u1101(.A(men_men_n1129_), .B(men_men_n1024_), .Y(men_men_n1130_));
  NOi41      u1102(.An(men_men_n827_), .B(men_men_n874_), .C(men_men_n863_), .D(men_men_n733_), .Y(men_men_n1131_));
  OAI220     u1103(.A0(men_men_n1131_), .A1(men_men_n707_), .B0(men_men_n1130_), .B1(men_men_n608_), .Y(men_men_n1132_));
  NOi31      u1104(.An(i), .B(k), .C(j), .Y(men_men_n1133_));
  NA4        u1105(.A(men_men_n1133_), .B(men_men_n1107_), .C(men_men_n347_), .D(men_men_n338_), .Y(men_men_n1134_));
  OAI210     u1106(.A0(men_men_n839_), .A1(men_men_n430_), .B0(men_men_n1134_), .Y(men_men_n1135_));
  NOi31      u1107(.An(m), .B(n), .C(f), .Y(men_men_n1136_));
  NA2        u1108(.A(men_men_n1136_), .B(men_men_n51_), .Y(men_men_n1137_));
  NO2        u1109(.A(men_men_n906_), .B(men_men_n436_), .Y(men_men_n1138_));
  NA2        u1110(.A(men_men_n522_), .B(l), .Y(men_men_n1139_));
  NOi31      u1111(.An(men_men_n885_), .B(men_men_n1061_), .C(men_men_n1139_), .Y(men_men_n1140_));
  NO3        u1112(.A(men_men_n1140_), .B(men_men_n1138_), .C(men_men_n1135_), .Y(men_men_n1141_));
  NO2        u1113(.A(men_men_n287_), .B(a), .Y(men_men_n1142_));
  INV        u1114(.A(men_men_n1068_), .Y(men_men_n1143_));
  NO2        u1115(.A(men_men_n1116_), .B(men_men_n499_), .Y(men_men_n1144_));
  NO2        u1116(.A(men_men_n89_), .B(u), .Y(men_men_n1145_));
  AOI210     u1117(.A0(men_men_n1145_), .A1(men_men_n1144_), .B0(men_men_n1099_), .Y(men_men_n1146_));
  OR2        u1118(.A(men_men_n1146_), .B(men_men_n1097_), .Y(men_men_n1147_));
  NA3        u1119(.A(men_men_n1147_), .B(men_men_n1143_), .C(men_men_n1141_), .Y(men_men_n1148_));
  NO4        u1120(.A(men_men_n1148_), .B(men_men_n1132_), .C(men_men_n840_), .D(men_men_n584_), .Y(men_men_n1149_));
  NA2        u1121(.A(c), .B(b), .Y(men_men_n1150_));
  NO2        u1122(.A(men_men_n719_), .B(men_men_n1150_), .Y(men_men_n1151_));
  OAI210     u1123(.A0(men_men_n883_), .A1(men_men_n854_), .B0(men_men_n423_), .Y(men_men_n1152_));
  OAI210     u1124(.A0(men_men_n1152_), .A1(men_men_n884_), .B0(men_men_n1151_), .Y(men_men_n1153_));
  NAi21      u1125(.An(men_men_n431_), .B(men_men_n1151_), .Y(men_men_n1154_));
  NA3        u1126(.A(men_men_n437_), .B(men_men_n577_), .C(f), .Y(men_men_n1155_));
  OAI210     u1127(.A0(men_men_n566_), .A1(men_men_n39_), .B0(men_men_n1142_), .Y(men_men_n1156_));
  NA3        u1128(.A(men_men_n1156_), .B(men_men_n1155_), .C(men_men_n1154_), .Y(men_men_n1157_));
  INV        u1129(.A(men_men_n120_), .Y(men_men_n1158_));
  OAI210     u1130(.A0(men_men_n1158_), .A1(men_men_n291_), .B0(u), .Y(men_men_n1159_));
  NAi21      u1131(.An(f), .B(d), .Y(men_men_n1160_));
  NO2        u1132(.A(men_men_n1160_), .B(men_men_n1120_), .Y(men_men_n1161_));
  INV        u1133(.A(men_men_n1161_), .Y(men_men_n1162_));
  AOI210     u1134(.A0(men_men_n1159_), .A1(men_men_n297_), .B0(men_men_n1162_), .Y(men_men_n1163_));
  AOI210     u1135(.A0(men_men_n1163_), .A1(men_men_n114_), .B0(men_men_n1157_), .Y(men_men_n1164_));
  NA2        u1136(.A(men_men_n482_), .B(men_men_n481_), .Y(men_men_n1165_));
  NO2        u1137(.A(men_men_n184_), .B(men_men_n241_), .Y(men_men_n1166_));
  NA2        u1138(.A(men_men_n1166_), .B(m), .Y(men_men_n1167_));
  NA3        u1139(.A(men_men_n940_), .B(men_men_n1139_), .C(men_men_n485_), .Y(men_men_n1168_));
  OAI210     u1140(.A0(men_men_n1168_), .A1(men_men_n314_), .B0(men_men_n483_), .Y(men_men_n1169_));
  AOI210     u1141(.A0(men_men_n1169_), .A1(men_men_n1165_), .B0(men_men_n1167_), .Y(men_men_n1170_));
  NA2        u1142(.A(men_men_n579_), .B(men_men_n418_), .Y(men_men_n1171_));
  NA2        u1143(.A(men_men_n160_), .B(men_men_n33_), .Y(men_men_n1172_));
  AOI210     u1144(.A0(men_men_n991_), .A1(men_men_n1172_), .B0(men_men_n218_), .Y(men_men_n1173_));
  OAI210     u1145(.A0(men_men_n1173_), .A1(men_men_n457_), .B0(men_men_n1161_), .Y(men_men_n1174_));
  NO2        u1146(.A(men_men_n379_), .B(men_men_n378_), .Y(men_men_n1175_));
  AOI210     u1147(.A0(men_men_n1166_), .A1(men_men_n439_), .B0(men_men_n985_), .Y(men_men_n1176_));
  NAi41      u1148(.An(men_men_n1175_), .B(men_men_n1176_), .C(men_men_n1174_), .D(men_men_n1171_), .Y(men_men_n1177_));
  NO2        u1149(.A(men_men_n1177_), .B(men_men_n1170_), .Y(men_men_n1178_));
  NA4        u1150(.A(men_men_n1178_), .B(men_men_n1164_), .C(men_men_n1153_), .D(men_men_n1149_), .Y(men00));
  AOI210     u1151(.A0(men_men_n300_), .A1(men_men_n218_), .B0(men_men_n279_), .Y(men_men_n1180_));
  NO2        u1152(.A(men_men_n1180_), .B(men_men_n598_), .Y(men_men_n1181_));
  AOI210     u1153(.A0(men_men_n920_), .A1(men_men_n967_), .B0(men_men_n1135_), .Y(men_men_n1182_));
  NO2        u1154(.A(men_men_n1113_), .B(men_men_n985_), .Y(men_men_n1183_));
  NA3        u1155(.A(men_men_n1183_), .B(men_men_n1182_), .C(men_men_n1025_), .Y(men_men_n1184_));
  NA2        u1156(.A(men_men_n524_), .B(f), .Y(men_men_n1185_));
  OAI210     u1157(.A0(men_men_n1032_), .A1(men_men_n40_), .B0(men_men_n660_), .Y(men_men_n1186_));
  NA3        u1158(.A(men_men_n1186_), .B(men_men_n259_), .C(n), .Y(men_men_n1187_));
  AOI210     u1159(.A0(men_men_n1187_), .A1(men_men_n1185_), .B0(men_men_n1072_), .Y(men_men_n1188_));
  NO4        u1160(.A(men_men_n1188_), .B(men_men_n1184_), .C(men_men_n1181_), .D(men_men_n1091_), .Y(men_men_n1189_));
  NA3        u1161(.A(men_men_n168_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1190_));
  NA3        u1162(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1191_));
  NOi31      u1163(.An(n), .B(m), .C(i), .Y(men_men_n1192_));
  NA3        u1164(.A(men_men_n1192_), .B(men_men_n663_), .C(men_men_n51_), .Y(men_men_n1193_));
  OAI210     u1165(.A0(men_men_n1191_), .A1(men_men_n1190_), .B0(men_men_n1193_), .Y(men_men_n1194_));
  INV        u1166(.A(men_men_n597_), .Y(men_men_n1195_));
  NO4        u1167(.A(men_men_n1195_), .B(men_men_n1194_), .C(men_men_n1175_), .D(men_men_n943_), .Y(men_men_n1196_));
  NO4        u1168(.A(men_men_n502_), .B(men_men_n361_), .C(men_men_n1150_), .D(men_men_n59_), .Y(men_men_n1197_));
  NA3        u1169(.A(men_men_n391_), .B(men_men_n225_), .C(u), .Y(men_men_n1198_));
  OA220      u1170(.A0(men_men_n1198_), .A1(men_men_n1191_), .B0(men_men_n392_), .B1(men_men_n137_), .Y(men_men_n1199_));
  NO2        u1171(.A(h), .B(u), .Y(men_men_n1200_));
  NA4        u1172(.A(men_men_n513_), .B(men_men_n479_), .C(men_men_n1200_), .D(men_men_n1060_), .Y(men_men_n1201_));
  NA2        u1173(.A(men_men_n972_), .B(men_men_n596_), .Y(men_men_n1202_));
  NA3        u1174(.A(men_men_n1202_), .B(men_men_n1201_), .C(men_men_n1199_), .Y(men_men_n1203_));
  NO3        u1175(.A(men_men_n1203_), .B(men_men_n1197_), .C(men_men_n269_), .Y(men_men_n1204_));
  INV        u1176(.A(men_men_n599_), .Y(men_men_n1205_));
  NA2        u1177(.A(men_men_n1205_), .B(men_men_n155_), .Y(men_men_n1206_));
  NA3        u1178(.A(men_men_n181_), .B(men_men_n113_), .C(u), .Y(men_men_n1207_));
  NA3        u1179(.A(men_men_n479_), .B(men_men_n40_), .C(f), .Y(men_men_n1208_));
  NOi31      u1180(.An(men_men_n892_), .B(men_men_n1208_), .C(men_men_n1207_), .Y(men_men_n1209_));
  NO2        u1181(.A(men_men_n278_), .B(men_men_n75_), .Y(men_men_n1210_));
  NO3        u1182(.A(men_men_n436_), .B(men_men_n850_), .C(n), .Y(men_men_n1211_));
  AOI210     u1183(.A0(men_men_n1211_), .A1(men_men_n1210_), .B0(men_men_n1106_), .Y(men_men_n1212_));
  NA2        u1184(.A(men_men_n1212_), .B(men_men_n74_), .Y(men_men_n1213_));
  NO4        u1185(.A(men_men_n1213_), .B(men_men_n1209_), .C(men_men_n1206_), .D(men_men_n534_), .Y(men_men_n1214_));
  AN3        u1186(.A(men_men_n1214_), .B(men_men_n1204_), .C(men_men_n1196_), .Y(men_men_n1215_));
  NA2        u1187(.A(men_men_n552_), .B(men_men_n102_), .Y(men_men_n1216_));
  NA3        u1188(.A(men_men_n1136_), .B(men_men_n623_), .C(men_men_n478_), .Y(men_men_n1217_));
  NA4        u1189(.A(men_men_n1217_), .B(men_men_n580_), .C(men_men_n1216_), .D(men_men_n246_), .Y(men_men_n1218_));
  OAI210     u1190(.A0(men_men_n477_), .A1(men_men_n121_), .B0(men_men_n886_), .Y(men_men_n1219_));
  AOI220     u1191(.A0(men_men_n1219_), .A1(men_men_n1168_), .B0(men_men_n579_), .B1(men_men_n418_), .Y(men_men_n1220_));
  NO2        u1192(.A(men_men_n221_), .B(men_men_n218_), .Y(men_men_n1221_));
  NA2        u1193(.A(n), .B(e), .Y(men_men_n1222_));
  NO2        u1194(.A(men_men_n1222_), .B(men_men_n147_), .Y(men_men_n1223_));
  AOI220     u1195(.A0(men_men_n1223_), .A1(men_men_n277_), .B0(men_men_n867_), .B1(men_men_n1221_), .Y(men_men_n1224_));
  OAI210     u1196(.A0(men_men_n362_), .A1(men_men_n315_), .B0(men_men_n459_), .Y(men_men_n1225_));
  NA3        u1197(.A(men_men_n1225_), .B(men_men_n1224_), .C(men_men_n1220_), .Y(men_men_n1226_));
  AOI210     u1198(.A0(men_men_n1223_), .A1(men_men_n871_), .B0(men_men_n840_), .Y(men_men_n1227_));
  AOI220     u1199(.A0(men_men_n981_), .A1(men_men_n596_), .B0(men_men_n663_), .B1(men_men_n249_), .Y(men_men_n1228_));
  NO2        u1200(.A(men_men_n68_), .B(h), .Y(men_men_n1229_));
  NO3        u1201(.A(men_men_n1072_), .B(men_men_n1070_), .C(men_men_n746_), .Y(men_men_n1230_));
  NO2        u1202(.A(men_men_n1103_), .B(men_men_n134_), .Y(men_men_n1231_));
  AN2        u1203(.A(men_men_n1231_), .B(men_men_n1118_), .Y(men_men_n1232_));
  OAI210     u1204(.A0(men_men_n1232_), .A1(men_men_n1230_), .B0(men_men_n1229_), .Y(men_men_n1233_));
  NA4        u1205(.A(men_men_n1233_), .B(men_men_n1228_), .C(men_men_n1227_), .D(men_men_n887_), .Y(men_men_n1234_));
  NO3        u1206(.A(men_men_n1234_), .B(men_men_n1226_), .C(men_men_n1218_), .Y(men_men_n1235_));
  NA2        u1207(.A(men_men_n855_), .B(men_men_n778_), .Y(men_men_n1236_));
  NA4        u1208(.A(men_men_n1236_), .B(men_men_n1235_), .C(men_men_n1215_), .D(men_men_n1189_), .Y(men01));
  AN2        u1209(.A(men_men_n1049_), .B(men_men_n1047_), .Y(men_men_n1238_));
  NO4        u1210(.A(men_men_n823_), .B(men_men_n816_), .C(men_men_n493_), .D(men_men_n285_), .Y(men_men_n1239_));
  NA2        u1211(.A(men_men_n402_), .B(i), .Y(men_men_n1240_));
  NA3        u1212(.A(men_men_n1240_), .B(men_men_n1239_), .C(men_men_n1238_), .Y(men_men_n1241_));
  NA2        u1213(.A(men_men_n572_), .B(men_men_n274_), .Y(men_men_n1242_));
  NA2        u1214(.A(men_men_n988_), .B(men_men_n1242_), .Y(men_men_n1243_));
  NA3        u1215(.A(men_men_n1243_), .B(men_men_n936_), .C(men_men_n337_), .Y(men_men_n1244_));
  NA2        u1216(.A(men_men_n45_), .B(f), .Y(men_men_n1245_));
  NA2        u1217(.A(men_men_n726_), .B(men_men_n97_), .Y(men_men_n1246_));
  NO2        u1218(.A(men_men_n1246_), .B(men_men_n1245_), .Y(men_men_n1247_));
  NA2        u1219(.A(men_men_n1247_), .B(men_men_n649_), .Y(men_men_n1248_));
  INV        u1220(.A(men_men_n119_), .Y(men_men_n1249_));
  OA220      u1221(.A0(men_men_n1249_), .A1(men_men_n606_), .B0(men_men_n676_), .B1(men_men_n376_), .Y(men_men_n1250_));
  NAi41      u1222(.An(men_men_n163_), .B(men_men_n1250_), .C(men_men_n1248_), .D(men_men_n919_), .Y(men_men_n1251_));
  NO3        u1223(.A(men_men_n804_), .B(men_men_n690_), .C(men_men_n527_), .Y(men_men_n1252_));
  OR2        u1224(.A(men_men_n198_), .B(men_men_n196_), .Y(men_men_n1253_));
  NA3        u1225(.A(men_men_n1253_), .B(men_men_n1252_), .C(men_men_n140_), .Y(men_men_n1254_));
  NO4        u1226(.A(men_men_n1254_), .B(men_men_n1251_), .C(men_men_n1244_), .D(men_men_n1241_), .Y(men_men_n1255_));
  INV        u1227(.A(men_men_n1198_), .Y(men_men_n1256_));
  OAI210     u1228(.A0(men_men_n1256_), .A1(men_men_n303_), .B0(men_men_n547_), .Y(men_men_n1257_));
  NA2        u1229(.A(men_men_n555_), .B(men_men_n404_), .Y(men_men_n1258_));
  NOi21      u1230(.An(men_men_n581_), .B(men_men_n603_), .Y(men_men_n1259_));
  NA2        u1231(.A(men_men_n1259_), .B(men_men_n1258_), .Y(men_men_n1260_));
  AOI210     u1232(.A0(men_men_n207_), .A1(men_men_n91_), .B0(men_men_n217_), .Y(men_men_n1261_));
  OAI210     u1233(.A0(men_men_n830_), .A1(men_men_n437_), .B0(men_men_n1261_), .Y(men_men_n1262_));
  AN3        u1234(.A(m), .B(l), .C(k), .Y(men_men_n1263_));
  OAI210     u1235(.A0(men_men_n364_), .A1(men_men_n34_), .B0(men_men_n1263_), .Y(men_men_n1264_));
  NA2        u1236(.A(men_men_n206_), .B(men_men_n34_), .Y(men_men_n1265_));
  AO210      u1237(.A0(men_men_n1265_), .A1(men_men_n1264_), .B0(men_men_n336_), .Y(men_men_n1266_));
  NA4        u1238(.A(men_men_n1266_), .B(men_men_n1262_), .C(men_men_n1260_), .D(men_men_n1257_), .Y(men_men_n1267_));
  INV        u1239(.A(men_men_n618_), .Y(men_men_n1268_));
  OAI210     u1240(.A0(men_men_n1249_), .A1(men_men_n615_), .B0(men_men_n1268_), .Y(men_men_n1269_));
  NA2        u1241(.A(men_men_n284_), .B(men_men_n198_), .Y(men_men_n1270_));
  NA2        u1242(.A(men_men_n1270_), .B(men_men_n681_), .Y(men_men_n1271_));
  NO3        u1243(.A(men_men_n839_), .B(men_men_n207_), .C(men_men_n416_), .Y(men_men_n1272_));
  NO2        u1244(.A(men_men_n1272_), .B(men_men_n985_), .Y(men_men_n1273_));
  OAI210     u1245(.A0(men_men_n1247_), .A1(men_men_n330_), .B0(men_men_n691_), .Y(men_men_n1274_));
  NA4        u1246(.A(men_men_n1274_), .B(men_men_n1273_), .C(men_men_n1271_), .D(men_men_n807_), .Y(men_men_n1275_));
  NO3        u1247(.A(men_men_n1275_), .B(men_men_n1269_), .C(men_men_n1267_), .Y(men_men_n1276_));
  NA2        u1248(.A(men_men_n519_), .B(men_men_n58_), .Y(men_men_n1277_));
  NO2        u1249(.A(men_men_n210_), .B(men_men_n112_), .Y(men_men_n1278_));
  NO2        u1250(.A(men_men_n1278_), .B(men_men_n1194_), .Y(men_men_n1279_));
  NA3        u1251(.A(men_men_n1279_), .B(men_men_n1277_), .C(men_men_n777_), .Y(men_men_n1280_));
  NO2        u1252(.A(men_men_n995_), .B(men_men_n237_), .Y(men_men_n1281_));
  NO2        u1253(.A(men_men_n996_), .B(men_men_n574_), .Y(men_men_n1282_));
  OAI210     u1254(.A0(men_men_n1282_), .A1(men_men_n1281_), .B0(men_men_n345_), .Y(men_men_n1283_));
  NA2        u1255(.A(men_men_n591_), .B(men_men_n589_), .Y(men_men_n1284_));
  NO3        u1256(.A(men_men_n81_), .B(men_men_n301_), .C(men_men_n45_), .Y(men_men_n1285_));
  NA2        u1257(.A(men_men_n1285_), .B(men_men_n571_), .Y(men_men_n1286_));
  NA2        u1258(.A(men_men_n1286_), .B(men_men_n1284_), .Y(men_men_n1287_));
  OR2        u1259(.A(men_men_n1198_), .B(men_men_n1191_), .Y(men_men_n1288_));
  NA2        u1260(.A(men_men_n1285_), .B(men_men_n833_), .Y(men_men_n1289_));
  NA3        u1261(.A(men_men_n1289_), .B(men_men_n1288_), .C(men_men_n394_), .Y(men_men_n1290_));
  NOi41      u1262(.An(men_men_n1283_), .B(men_men_n1290_), .C(men_men_n1287_), .D(men_men_n1280_), .Y(men_men_n1291_));
  NO2        u1263(.A(men_men_n133_), .B(men_men_n45_), .Y(men_men_n1292_));
  NO2        u1264(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1293_));
  AO220      u1265(.A0(men_men_n1293_), .A1(men_men_n637_), .B0(men_men_n1292_), .B1(men_men_n724_), .Y(men_men_n1294_));
  NA2        u1266(.A(men_men_n1294_), .B(men_men_n345_), .Y(men_men_n1295_));
  NO3        u1267(.A(men_men_n1116_), .B(men_men_n178_), .C(men_men_n89_), .Y(men_men_n1296_));
  NA2        u1268(.A(men_men_n1285_), .B(men_men_n999_), .Y(men_men_n1297_));
  NA2        u1269(.A(men_men_n1297_), .B(men_men_n1295_), .Y(men_men_n1298_));
  NO2        u1270(.A(men_men_n628_), .B(men_men_n627_), .Y(men_men_n1299_));
  NO4        u1271(.A(men_men_n1116_), .B(men_men_n1299_), .C(men_men_n176_), .D(men_men_n89_), .Y(men_men_n1300_));
  NO3        u1272(.A(men_men_n1300_), .B(men_men_n1298_), .C(men_men_n652_), .Y(men_men_n1301_));
  NA4        u1273(.A(men_men_n1301_), .B(men_men_n1291_), .C(men_men_n1276_), .D(men_men_n1255_), .Y(men06));
  NO2        u1274(.A(men_men_n417_), .B(men_men_n578_), .Y(men_men_n1303_));
  INV        u1275(.A(men_men_n753_), .Y(men_men_n1304_));
  NA2        u1276(.A(men_men_n1304_), .B(men_men_n1303_), .Y(men_men_n1305_));
  NO2        u1277(.A(men_men_n229_), .B(men_men_n103_), .Y(men_men_n1306_));
  OAI210     u1278(.A0(men_men_n1306_), .A1(men_men_n1296_), .B0(men_men_n390_), .Y(men_men_n1307_));
  NO3        u1279(.A(men_men_n619_), .B(men_men_n828_), .C(men_men_n620_), .Y(men_men_n1308_));
  OR2        u1280(.A(men_men_n1308_), .B(men_men_n906_), .Y(men_men_n1309_));
  NA4        u1281(.A(men_men_n1309_), .B(men_men_n1307_), .C(men_men_n1305_), .D(men_men_n1283_), .Y(men_men_n1310_));
  NO3        u1282(.A(men_men_n1310_), .B(men_men_n1287_), .C(men_men_n258_), .Y(men_men_n1311_));
  NO2        u1283(.A(men_men_n301_), .B(men_men_n45_), .Y(men_men_n1312_));
  AOI210     u1284(.A0(men_men_n1312_), .A1(men_men_n1000_), .B0(men_men_n1281_), .Y(men_men_n1313_));
  AOI210     u1285(.A0(men_men_n1312_), .A1(men_men_n575_), .B0(men_men_n1294_), .Y(men_men_n1314_));
  AOI210     u1286(.A0(men_men_n1314_), .A1(men_men_n1313_), .B0(men_men_n342_), .Y(men_men_n1315_));
  OAI210     u1287(.A0(men_men_n91_), .A1(men_men_n40_), .B0(men_men_n689_), .Y(men_men_n1316_));
  NA2        u1288(.A(men_men_n1316_), .B(men_men_n656_), .Y(men_men_n1317_));
  NO2        u1289(.A(men_men_n530_), .B(men_men_n173_), .Y(men_men_n1318_));
  NOi21      u1290(.An(men_men_n139_), .B(men_men_n45_), .Y(men_men_n1319_));
  NO2        u1291(.A(men_men_n624_), .B(men_men_n1137_), .Y(men_men_n1320_));
  OAI210     u1292(.A0(men_men_n472_), .A1(men_men_n251_), .B0(men_men_n930_), .Y(men_men_n1321_));
  NO4        u1293(.A(men_men_n1321_), .B(men_men_n1320_), .C(men_men_n1319_), .D(men_men_n1318_), .Y(men_men_n1322_));
  NO2        u1294(.A(men_men_n375_), .B(men_men_n138_), .Y(men_men_n1323_));
  AOI210     u1295(.A0(men_men_n1323_), .A1(men_men_n609_), .B0(men_men_n618_), .Y(men_men_n1324_));
  NA3        u1296(.A(men_men_n1324_), .B(men_men_n1322_), .C(men_men_n1317_), .Y(men_men_n1325_));
  NO2        u1297(.A(men_men_n769_), .B(men_men_n374_), .Y(men_men_n1326_));
  NO3        u1298(.A(men_men_n691_), .B(men_men_n779_), .C(men_men_n649_), .Y(men_men_n1327_));
  NOi21      u1299(.An(men_men_n1326_), .B(men_men_n1327_), .Y(men_men_n1328_));
  AN2        u1300(.A(men_men_n981_), .B(men_men_n659_), .Y(men_men_n1329_));
  NO4        u1301(.A(men_men_n1329_), .B(men_men_n1328_), .C(men_men_n1325_), .D(men_men_n1315_), .Y(men_men_n1330_));
  NO2        u1302(.A(men_men_n822_), .B(men_men_n280_), .Y(men_men_n1331_));
  OAI220     u1303(.A0(men_men_n753_), .A1(men_men_n47_), .B0(men_men_n229_), .B1(men_men_n630_), .Y(men_men_n1332_));
  OAI210     u1304(.A0(men_men_n280_), .A1(c), .B0(men_men_n655_), .Y(men_men_n1333_));
  AOI220     u1305(.A0(men_men_n1333_), .A1(men_men_n1332_), .B0(men_men_n1331_), .B1(men_men_n270_), .Y(men_men_n1334_));
  NO3        u1306(.A(men_men_n248_), .B(men_men_n103_), .C(men_men_n287_), .Y(men_men_n1335_));
  OAI220     u1307(.A0(men_men_n716_), .A1(men_men_n251_), .B0(men_men_n526_), .B1(men_men_n530_), .Y(men_men_n1336_));
  OAI210     u1308(.A0(l), .A1(i), .B0(k), .Y(men_men_n1337_));
  NO3        u1309(.A(men_men_n1337_), .B(men_men_n617_), .C(j), .Y(men_men_n1338_));
  NOi21      u1310(.An(men_men_n1338_), .B(men_men_n685_), .Y(men_men_n1339_));
  NO4        u1311(.A(men_men_n1339_), .B(men_men_n1336_), .C(men_men_n1335_), .D(men_men_n1138_), .Y(men_men_n1340_));
  NA4        u1312(.A(men_men_n814_), .B(men_men_n813_), .C(men_men_n447_), .D(men_men_n899_), .Y(men_men_n1341_));
  NAi31      u1313(.An(men_men_n769_), .B(men_men_n1341_), .C(men_men_n206_), .Y(men_men_n1342_));
  NA4        u1314(.A(men_men_n1342_), .B(men_men_n1340_), .C(men_men_n1334_), .D(men_men_n1228_), .Y(men_men_n1343_));
  NOi31      u1315(.An(men_men_n1308_), .B(men_men_n476_), .C(men_men_n403_), .Y(men_men_n1344_));
  OR3        u1316(.A(men_men_n1344_), .B(men_men_n803_), .C(men_men_n558_), .Y(men_men_n1345_));
  OR3        u1317(.A(men_men_n378_), .B(men_men_n229_), .C(men_men_n630_), .Y(men_men_n1346_));
  AOI210     u1318(.A0(men_men_n591_), .A1(men_men_n459_), .B0(men_men_n380_), .Y(men_men_n1347_));
  NA3        u1319(.A(men_men_n1347_), .B(men_men_n1346_), .C(men_men_n1345_), .Y(men_men_n1348_));
  AN2        u1320(.A(men_men_n952_), .B(men_men_n951_), .Y(men_men_n1349_));
  NO4        u1321(.A(men_men_n1349_), .B(men_men_n897_), .C(men_men_n515_), .D(men_men_n496_), .Y(men_men_n1350_));
  NA2        u1322(.A(men_men_n1350_), .B(men_men_n1289_), .Y(men_men_n1351_));
  NAi21      u1323(.An(j), .B(i), .Y(men_men_n1352_));
  NO4        u1324(.A(men_men_n1299_), .B(men_men_n1352_), .C(men_men_n453_), .D(men_men_n239_), .Y(men_men_n1353_));
  NO4        u1325(.A(men_men_n1353_), .B(men_men_n1351_), .C(men_men_n1348_), .D(men_men_n1343_), .Y(men_men_n1354_));
  NA4        u1326(.A(men_men_n1354_), .B(men_men_n1330_), .C(men_men_n1311_), .D(men_men_n1301_), .Y(men07));
  NOi21      u1327(.An(j), .B(k), .Y(men_men_n1356_));
  NA4        u1328(.A(men_men_n181_), .B(men_men_n109_), .C(men_men_n1356_), .D(f), .Y(men_men_n1357_));
  NAi32      u1329(.An(m), .Bn(b), .C(n), .Y(men_men_n1358_));
  NO3        u1330(.A(men_men_n1358_), .B(u), .C(f), .Y(men_men_n1359_));
  OAI210     u1331(.A0(men_men_n325_), .A1(men_men_n498_), .B0(men_men_n1359_), .Y(men_men_n1360_));
  NAi21      u1332(.An(f), .B(c), .Y(men_men_n1361_));
  OR2        u1333(.A(e), .B(d), .Y(men_men_n1362_));
  OAI220     u1334(.A0(men_men_n1362_), .A1(men_men_n1361_), .B0(men_men_n643_), .B1(men_men_n326_), .Y(men_men_n1363_));
  NA3        u1335(.A(men_men_n1363_), .B(men_men_n1081_), .C(men_men_n181_), .Y(men_men_n1364_));
  NOi31      u1336(.An(n), .B(m), .C(b), .Y(men_men_n1365_));
  NO3        u1337(.A(men_men_n134_), .B(men_men_n461_), .C(h), .Y(men_men_n1366_));
  NA3        u1338(.A(men_men_n1364_), .B(men_men_n1360_), .C(men_men_n1357_), .Y(men_men_n1367_));
  NOi41      u1339(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1368_));
  NO2        u1340(.A(k), .B(i), .Y(men_men_n1369_));
  NA3        u1341(.A(men_men_n1369_), .B(men_men_n918_), .C(men_men_n181_), .Y(men_men_n1370_));
  NO2        u1342(.A(men_men_n1088_), .B(men_men_n309_), .Y(men_men_n1371_));
  NA2        u1343(.A(men_men_n559_), .B(men_men_n82_), .Y(men_men_n1372_));
  NA2        u1344(.A(men_men_n1229_), .B(men_men_n295_), .Y(men_men_n1373_));
  NA3        u1345(.A(men_men_n1373_), .B(men_men_n1372_), .C(men_men_n1370_), .Y(men_men_n1374_));
  NO2        u1346(.A(men_men_n1374_), .B(men_men_n1367_), .Y(men_men_n1375_));
  NO3        u1347(.A(e), .B(d), .C(c), .Y(men_men_n1376_));
  NO2        u1348(.A(men_men_n134_), .B(men_men_n218_), .Y(men_men_n1377_));
  NA2        u1349(.A(men_men_n1377_), .B(men_men_n1376_), .Y(men_men_n1378_));
  NO2        u1350(.A(men_men_n1378_), .B(c), .Y(men_men_n1379_));
  OR2        u1351(.A(h), .B(f), .Y(men_men_n1380_));
  NO3        u1352(.A(n), .B(m), .C(i), .Y(men_men_n1381_));
  OAI210     u1353(.A0(c), .A1(men_men_n158_), .B0(men_men_n1381_), .Y(men_men_n1382_));
  NO2        u1354(.A(i), .B(u), .Y(men_men_n1383_));
  OR3        u1355(.A(men_men_n1383_), .B(men_men_n1358_), .C(men_men_n72_), .Y(men_men_n1384_));
  OAI220     u1356(.A0(men_men_n1384_), .A1(men_men_n498_), .B0(men_men_n1382_), .B1(men_men_n1380_), .Y(men_men_n1385_));
  NA3        u1357(.A(men_men_n713_), .B(men_men_n699_), .C(men_men_n113_), .Y(men_men_n1386_));
  NO2        u1358(.A(men_men_n1386_), .B(men_men_n45_), .Y(men_men_n1387_));
  NO2        u1359(.A(l), .B(k), .Y(men_men_n1388_));
  NOi41      u1360(.An(men_men_n564_), .B(men_men_n1388_), .C(men_men_n491_), .D(men_men_n453_), .Y(men_men_n1389_));
  NO3        u1361(.A(men_men_n453_), .B(d), .C(c), .Y(men_men_n1390_));
  NO4        u1362(.A(men_men_n1389_), .B(men_men_n1387_), .C(men_men_n1385_), .D(men_men_n1379_), .Y(men_men_n1391_));
  NO2        u1363(.A(men_men_n148_), .B(h), .Y(men_men_n1392_));
  NO2        u1364(.A(men_men_n1098_), .B(l), .Y(men_men_n1393_));
  NO2        u1365(.A(u), .B(c), .Y(men_men_n1394_));
  NA3        u1366(.A(men_men_n1394_), .B(men_men_n144_), .C(men_men_n189_), .Y(men_men_n1395_));
  NO2        u1367(.A(men_men_n1395_), .B(men_men_n1393_), .Y(men_men_n1396_));
  NA2        u1368(.A(men_men_n1396_), .B(men_men_n181_), .Y(men_men_n1397_));
  NO2        u1369(.A(men_men_n463_), .B(a), .Y(men_men_n1398_));
  NA3        u1370(.A(men_men_n1398_), .B(k), .C(men_men_n114_), .Y(men_men_n1399_));
  NO2        u1371(.A(i), .B(h), .Y(men_men_n1400_));
  NA2        u1372(.A(men_men_n1400_), .B(men_men_n225_), .Y(men_men_n1401_));
  AOI210     u1373(.A0(men_men_n1160_), .A1(h), .B0(men_men_n424_), .Y(men_men_n1402_));
  NA2        u1374(.A(men_men_n141_), .B(men_men_n225_), .Y(men_men_n1403_));
  AOI210     u1375(.A0(men_men_n259_), .A1(men_men_n117_), .B0(men_men_n547_), .Y(men_men_n1404_));
  OAI220     u1376(.A0(men_men_n1404_), .A1(men_men_n1401_), .B0(men_men_n1403_), .B1(men_men_n1402_), .Y(men_men_n1405_));
  NO2        u1377(.A(men_men_n775_), .B(men_men_n190_), .Y(men_men_n1406_));
  NOi31      u1378(.An(m), .B(n), .C(b), .Y(men_men_n1407_));
  NOi31      u1379(.An(f), .B(d), .C(c), .Y(men_men_n1408_));
  NA2        u1380(.A(men_men_n1408_), .B(men_men_n1407_), .Y(men_men_n1409_));
  INV        u1381(.A(men_men_n1409_), .Y(men_men_n1410_));
  NO3        u1382(.A(men_men_n1410_), .B(men_men_n1406_), .C(men_men_n1405_), .Y(men_men_n1411_));
  NA2        u1383(.A(men_men_n1109_), .B(men_men_n479_), .Y(men_men_n1412_));
  NO4        u1384(.A(men_men_n1412_), .B(men_men_n1083_), .C(men_men_n453_), .D(men_men_n45_), .Y(men_men_n1413_));
  OAI210     u1385(.A0(men_men_n184_), .A1(men_men_n542_), .B0(men_men_n1084_), .Y(men_men_n1414_));
  NO3        u1386(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1415_));
  INV        u1387(.A(men_men_n1414_), .Y(men_men_n1416_));
  NO2        u1388(.A(men_men_n1416_), .B(men_men_n1413_), .Y(men_men_n1417_));
  AN4        u1389(.A(men_men_n1417_), .B(men_men_n1411_), .C(men_men_n1399_), .D(men_men_n1397_), .Y(men_men_n1418_));
  NA2        u1390(.A(men_men_n1365_), .B(men_men_n387_), .Y(men_men_n1419_));
  NO2        u1391(.A(men_men_n1419_), .B(men_men_n1069_), .Y(men_men_n1420_));
  NA2        u1392(.A(men_men_n1390_), .B(men_men_n219_), .Y(men_men_n1421_));
  NO2        u1393(.A(men_men_n190_), .B(b), .Y(men_men_n1422_));
  AOI220     u1394(.A0(men_men_n1192_), .A1(men_men_n1422_), .B0(men_men_n1117_), .B1(men_men_n1412_), .Y(men_men_n1423_));
  NO2        u1395(.A(i), .B(men_men_n217_), .Y(men_men_n1424_));
  NA4        u1396(.A(men_men_n1166_), .B(men_men_n1424_), .C(men_men_n104_), .D(m), .Y(men_men_n1425_));
  NAi41      u1397(.An(men_men_n1420_), .B(men_men_n1425_), .C(men_men_n1423_), .D(men_men_n1421_), .Y(men_men_n1426_));
  NO4        u1398(.A(men_men_n134_), .B(u), .C(f), .D(e), .Y(men_men_n1427_));
  NA3        u1399(.A(men_men_n1369_), .B(men_men_n296_), .C(h), .Y(men_men_n1428_));
  OR2        u1400(.A(e), .B(a), .Y(men_men_n1429_));
  NA2        u1401(.A(men_men_n30_), .B(h), .Y(men_men_n1430_));
  NO2        u1402(.A(men_men_n1430_), .B(men_men_n1105_), .Y(men_men_n1431_));
  NOi41      u1403(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1432_));
  NA2        u1404(.A(men_men_n1432_), .B(men_men_n114_), .Y(men_men_n1433_));
  NA2        u1405(.A(men_men_n1368_), .B(men_men_n1388_), .Y(men_men_n1434_));
  NA2        u1406(.A(men_men_n1434_), .B(men_men_n1433_), .Y(men_men_n1435_));
  NA2        u1407(.A(men_men_n1136_), .B(men_men_n416_), .Y(men_men_n1436_));
  NO2        u1408(.A(men_men_n1436_), .B(men_men_n446_), .Y(men_men_n1437_));
  AO210      u1409(.A0(men_men_n1437_), .A1(men_men_n117_), .B0(men_men_n1435_), .Y(men_men_n1438_));
  NO3        u1410(.A(men_men_n1438_), .B(men_men_n1431_), .C(men_men_n1426_), .Y(men_men_n1439_));
  NA4        u1411(.A(men_men_n1439_), .B(men_men_n1418_), .C(men_men_n1391_), .D(men_men_n1375_), .Y(men_men_n1440_));
  NO2        u1412(.A(men_men_n1150_), .B(men_men_n111_), .Y(men_men_n1441_));
  NA2        u1413(.A(men_men_n387_), .B(men_men_n56_), .Y(men_men_n1442_));
  NA2        u1414(.A(men_men_n219_), .B(men_men_n181_), .Y(men_men_n1443_));
  AOI210     u1415(.A0(men_men_n1443_), .A1(men_men_n1207_), .B0(men_men_n1442_), .Y(men_men_n1444_));
  NO2        u1416(.A(men_men_n399_), .B(j), .Y(men_men_n1445_));
  NA3        u1417(.A(men_men_n1415_), .B(men_men_n1362_), .C(men_men_n1136_), .Y(men_men_n1446_));
  NAi41      u1418(.An(men_men_n1400_), .B(men_men_n1096_), .C(men_men_n169_), .D(men_men_n151_), .Y(men_men_n1447_));
  NA2        u1419(.A(men_men_n1447_), .B(men_men_n1446_), .Y(men_men_n1448_));
  NA3        u1420(.A(u), .B(men_men_n1445_), .C(men_men_n160_), .Y(men_men_n1449_));
  INV        u1421(.A(men_men_n1449_), .Y(men_men_n1450_));
  NO3        u1422(.A(men_men_n769_), .B(men_men_n176_), .C(men_men_n419_), .Y(men_men_n1451_));
  NO3        u1423(.A(men_men_n1451_), .B(men_men_n1450_), .C(men_men_n1448_), .Y(men_men_n1452_));
  NO2        u1424(.A(men_men_n1562_), .B(men_men_n1076_), .Y(men_men_n1453_));
  OR2        u1425(.A(n), .B(i), .Y(men_men_n1454_));
  OAI210     u1426(.A0(men_men_n1454_), .A1(men_men_n1095_), .B0(men_men_n49_), .Y(men_men_n1455_));
  AOI220     u1427(.A0(men_men_n1455_), .A1(men_men_n1200_), .B0(men_men_n843_), .B1(men_men_n197_), .Y(men_men_n1456_));
  INV        u1428(.A(men_men_n1456_), .Y(men_men_n1457_));
  OAI220     u1429(.A0(men_men_n682_), .A1(u), .B0(men_men_n229_), .B1(c), .Y(men_men_n1458_));
  AOI210     u1430(.A0(men_men_n1422_), .A1(men_men_n41_), .B0(men_men_n1458_), .Y(men_men_n1459_));
  NO2        u1431(.A(men_men_n134_), .B(l), .Y(men_men_n1460_));
  NO2        u1432(.A(men_men_n229_), .B(k), .Y(men_men_n1461_));
  OAI210     u1433(.A0(men_men_n1461_), .A1(men_men_n1400_), .B0(men_men_n1460_), .Y(men_men_n1462_));
  OAI220     u1434(.A0(men_men_n1462_), .A1(men_men_n31_), .B0(men_men_n1459_), .B1(men_men_n178_), .Y(men_men_n1463_));
  NO3        u1435(.A(men_men_n1463_), .B(men_men_n1457_), .C(men_men_n1453_), .Y(men_men_n1464_));
  NO3        u1436(.A(men_men_n1120_), .B(men_men_n1362_), .C(men_men_n49_), .Y(men_men_n1465_));
  NO2        u1437(.A(men_men_n1105_), .B(h), .Y(men_men_n1466_));
  NA3        u1438(.A(men_men_n1466_), .B(d), .C(men_men_n1070_), .Y(men_men_n1467_));
  NO2        u1439(.A(men_men_n1467_), .B(c), .Y(men_men_n1468_));
  NA3        u1440(.A(men_men_n1441_), .B(men_men_n479_), .C(f), .Y(men_men_n1469_));
  NA2        u1441(.A(men_men_n181_), .B(men_men_n113_), .Y(men_men_n1470_));
  NO2        u1442(.A(men_men_n1356_), .B(men_men_n42_), .Y(men_men_n1471_));
  AOI210     u1443(.A0(men_men_n114_), .A1(men_men_n40_), .B0(men_men_n1471_), .Y(men_men_n1472_));
  NO2        u1444(.A(men_men_n1472_), .B(men_men_n1469_), .Y(men_men_n1473_));
  AOI210     u1445(.A0(men_men_n542_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1474_));
  NA2        u1446(.A(men_men_n1474_), .B(men_men_n1398_), .Y(men_men_n1475_));
  NO2        u1447(.A(men_men_n1352_), .B(men_men_n176_), .Y(men_men_n1476_));
  NOi21      u1448(.An(d), .B(f), .Y(men_men_n1477_));
  NO3        u1449(.A(men_men_n1408_), .B(men_men_n1477_), .C(men_men_n40_), .Y(men_men_n1478_));
  NA2        u1450(.A(men_men_n1478_), .B(men_men_n1476_), .Y(men_men_n1479_));
  NO2        u1451(.A(men_men_n1362_), .B(f), .Y(men_men_n1480_));
  NA2        u1452(.A(men_men_n1398_), .B(men_men_n1471_), .Y(men_men_n1481_));
  NO2        u1453(.A(men_men_n301_), .B(c), .Y(men_men_n1482_));
  NA2        u1454(.A(men_men_n1482_), .B(men_men_n559_), .Y(men_men_n1483_));
  NA4        u1455(.A(men_men_n1483_), .B(men_men_n1481_), .C(men_men_n1479_), .D(men_men_n1475_), .Y(men_men_n1484_));
  NO3        u1456(.A(men_men_n1484_), .B(men_men_n1473_), .C(men_men_n1468_), .Y(men_men_n1485_));
  NA4        u1457(.A(men_men_n1485_), .B(men_men_n1464_), .C(men_men_n1452_), .D(men_men_n1563_), .Y(men_men_n1486_));
  NO3        u1458(.A(men_men_n1109_), .B(men_men_n1095_), .C(men_men_n40_), .Y(men_men_n1487_));
  NO2        u1459(.A(men_men_n479_), .B(men_men_n301_), .Y(men_men_n1488_));
  OAI210     u1460(.A0(men_men_n1488_), .A1(men_men_n1487_), .B0(men_men_n1371_), .Y(men_men_n1489_));
  OAI210     u1461(.A0(men_men_n1427_), .A1(men_men_n1365_), .B0(men_men_n903_), .Y(men_men_n1490_));
  NO2        u1462(.A(men_men_n1066_), .B(men_men_n134_), .Y(men_men_n1491_));
  NA2        u1463(.A(men_men_n1491_), .B(men_men_n636_), .Y(men_men_n1492_));
  NA3        u1464(.A(men_men_n1492_), .B(men_men_n1490_), .C(men_men_n1489_), .Y(men_men_n1493_));
  NA2        u1465(.A(men_men_n1394_), .B(men_men_n1477_), .Y(men_men_n1494_));
  NO2        u1466(.A(men_men_n1494_), .B(m), .Y(men_men_n1495_));
  NO2        u1467(.A(men_men_n152_), .B(men_men_n183_), .Y(men_men_n1496_));
  OAI210     u1468(.A0(men_men_n1496_), .A1(men_men_n111_), .B0(men_men_n1407_), .Y(men_men_n1497_));
  INV        u1469(.A(men_men_n1497_), .Y(men_men_n1498_));
  NO3        u1470(.A(men_men_n1498_), .B(men_men_n1495_), .C(men_men_n1493_), .Y(men_men_n1499_));
  NO2        u1471(.A(men_men_n1361_), .B(e), .Y(men_men_n1500_));
  NA2        u1472(.A(men_men_n1500_), .B(men_men_n414_), .Y(men_men_n1501_));
  NA2        u1473(.A(men_men_n1145_), .B(men_men_n645_), .Y(men_men_n1502_));
  OR3        u1474(.A(men_men_n1461_), .B(men_men_n1229_), .C(men_men_n134_), .Y(men_men_n1503_));
  OAI220     u1475(.A0(men_men_n1503_), .A1(men_men_n1501_), .B0(men_men_n1502_), .B1(men_men_n455_), .Y(men_men_n1504_));
  INV        u1476(.A(men_men_n1504_), .Y(men_men_n1505_));
  NO2        u1477(.A(men_men_n183_), .B(c), .Y(men_men_n1506_));
  NA2        u1478(.A(men_men_n1506_), .B(men_men_n181_), .Y(men_men_n1507_));
  AOI220     u1479(.A0(men_men_n1507_), .A1(men_men_n1097_), .B0(men_men_n549_), .B1(men_men_n374_), .Y(men_men_n1508_));
  NA2        u1480(.A(men_men_n557_), .B(u), .Y(men_men_n1509_));
  AOI210     u1481(.A0(men_men_n1509_), .A1(men_men_n1390_), .B0(men_men_n1465_), .Y(men_men_n1510_));
  NO2        u1482(.A(men_men_n1429_), .B(f), .Y(men_men_n1511_));
  AOI210     u1483(.A0(men_men_n1145_), .A1(a), .B0(men_men_n1511_), .Y(men_men_n1512_));
  OAI220     u1484(.A0(men_men_n1512_), .A1(men_men_n69_), .B0(men_men_n1510_), .B1(men_men_n217_), .Y(men_men_n1513_));
  AOI210     u1485(.A0(men_men_n923_), .A1(men_men_n426_), .B0(men_men_n105_), .Y(men_men_n1514_));
  OR2        u1486(.A(men_men_n1514_), .B(men_men_n557_), .Y(men_men_n1515_));
  NO2        u1487(.A(men_men_n1515_), .B(men_men_n176_), .Y(men_men_n1516_));
  NA4        u1488(.A(men_men_n1118_), .B(men_men_n1115_), .C(men_men_n225_), .D(men_men_n68_), .Y(men_men_n1517_));
  NA2        u1489(.A(men_men_n1366_), .B(men_men_n184_), .Y(men_men_n1518_));
  NO2        u1490(.A(men_men_n49_), .B(l), .Y(men_men_n1519_));
  OAI210     u1491(.A0(men_men_n1429_), .A1(men_men_n882_), .B0(men_men_n498_), .Y(men_men_n1520_));
  OAI210     u1492(.A0(men_men_n1520_), .A1(men_men_n1121_), .B0(men_men_n1519_), .Y(men_men_n1521_));
  NO2        u1493(.A(men_men_n254_), .B(u), .Y(men_men_n1522_));
  NO2        u1494(.A(m), .B(i), .Y(men_men_n1523_));
  BUFFER     u1495(.A(men_men_n1523_), .Y(men_men_n1524_));
  AOI220     u1496(.A0(men_men_n1524_), .A1(men_men_n1392_), .B0(men_men_n1096_), .B1(men_men_n1522_), .Y(men_men_n1525_));
  NA4        u1497(.A(men_men_n1525_), .B(men_men_n1521_), .C(men_men_n1518_), .D(men_men_n1517_), .Y(men_men_n1526_));
  NO4        u1498(.A(men_men_n1526_), .B(men_men_n1516_), .C(men_men_n1513_), .D(men_men_n1508_), .Y(men_men_n1527_));
  NA3        u1499(.A(men_men_n1527_), .B(men_men_n1505_), .C(men_men_n1499_), .Y(men_men_n1528_));
  NA3        u1500(.A(men_men_n987_), .B(men_men_n141_), .C(men_men_n46_), .Y(men_men_n1529_));
  AOI210     u1501(.A0(men_men_n149_), .A1(c), .B0(men_men_n1529_), .Y(men_men_n1530_));
  INV        u1502(.A(men_men_n187_), .Y(men_men_n1531_));
  NA2        u1503(.A(men_men_n1531_), .B(men_men_n1466_), .Y(men_men_n1532_));
  OR2        u1504(.A(men_men_n135_), .B(men_men_n1419_), .Y(men_men_n1533_));
  NO2        u1505(.A(men_men_n72_), .B(c), .Y(men_men_n1534_));
  NA2        u1506(.A(men_men_n1476_), .B(men_men_n1534_), .Y(men_men_n1535_));
  NA3        u1507(.A(men_men_n1535_), .B(men_men_n1533_), .C(men_men_n1532_), .Y(men_men_n1536_));
  NO2        u1508(.A(men_men_n1536_), .B(men_men_n1530_), .Y(men_men_n1537_));
  NA2        u1509(.A(men_men_n158_), .B(men_men_n56_), .Y(men_men_n1538_));
  NO2        u1510(.A(men_men_n1538_), .B(men_men_n1470_), .Y(men_men_n1539_));
  NOi21      u1511(.An(men_men_n1366_), .B(e), .Y(men_men_n1540_));
  NO2        u1512(.A(men_men_n1540_), .B(men_men_n1539_), .Y(men_men_n1541_));
  AN2        u1513(.A(men_men_n1118_), .B(men_men_n1103_), .Y(men_men_n1542_));
  AOI220     u1514(.A0(men_men_n1523_), .A1(men_men_n654_), .B0(men_men_n1081_), .B1(men_men_n161_), .Y(men_men_n1543_));
  NOi31      u1515(.An(men_men_n30_), .B(men_men_n1543_), .C(n), .Y(men_men_n1544_));
  AOI210     u1516(.A0(men_men_n1542_), .A1(men_men_n1192_), .B0(men_men_n1544_), .Y(men_men_n1545_));
  NA2        u1517(.A(men_men_n59_), .B(a), .Y(men_men_n1546_));
  NO2        u1518(.A(men_men_n1369_), .B(men_men_n119_), .Y(men_men_n1547_));
  OAI220     u1519(.A0(men_men_n1547_), .A1(men_men_n1419_), .B0(men_men_n1436_), .B1(men_men_n1546_), .Y(men_men_n1548_));
  INV        u1520(.A(men_men_n1548_), .Y(men_men_n1549_));
  NA4        u1521(.A(men_men_n1549_), .B(men_men_n1545_), .C(men_men_n1541_), .D(men_men_n1537_), .Y(men_men_n1550_));
  OR4        u1522(.A(men_men_n1550_), .B(men_men_n1528_), .C(men_men_n1486_), .D(men_men_n1440_), .Y(men04));
  NOi31      u1523(.An(men_men_n1427_), .B(men_men_n1428_), .C(men_men_n1072_), .Y(men_men_n1552_));
  NA2        u1524(.A(men_men_n1480_), .B(men_men_n843_), .Y(men_men_n1553_));
  NO3        u1525(.A(men_men_n1553_), .B(men_men_n1061_), .C(men_men_n499_), .Y(men_men_n1554_));
  OR3        u1526(.A(men_men_n1554_), .B(men_men_n1552_), .C(men_men_n1086_), .Y(men_men_n1555_));
  INV        u1527(.A(men_men_n1209_), .Y(men_men_n1556_));
  NA2        u1528(.A(men_men_n1556_), .B(men_men_n1233_), .Y(men_men_n1557_));
  NO4        u1529(.A(men_men_n1557_), .B(men_men_n1555_), .C(men_men_n1094_), .D(men_men_n1075_), .Y(men_men_n1558_));
  NA4        u1530(.A(men_men_n1558_), .B(men_men_n1147_), .C(men_men_n1134_), .D(men_men_n1124_), .Y(men05));
  INV        u1531(.A(men_men_n181_), .Y(men_men_n1562_));
  INV        u1532(.A(men_men_n1444_), .Y(men_men_n1563_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule