//Benchmark atmr_misex3_1774_0.5

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1597_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, men_men_n1605_, men_men_n1606_, men_men_n1607_, men_men_n1608_, men_men_n1609_, men_men_n1610_, men_men_n1611_, men_men_n1612_, men_men_n1613_, men_men_n1614_, men_men_n1615_, men_men_n1616_, men_men_n1617_, men_men_n1618_, men_men_n1619_, men_men_n1620_, men_men_n1621_, men_men_n1622_, men_men_n1623_, men_men_n1624_, men_men_n1625_, men_men_n1626_, men_men_n1627_, men_men_n1628_, men_men_n1629_, men_men_n1630_, men_men_n1631_, men_men_n1632_, men_men_n1633_, men_men_n1634_, men_men_n1635_, men_men_n1636_, men_men_n1637_, men_men_n1638_, men_men_n1639_, men_men_n1640_, men_men_n1641_, men_men_n1642_, men_men_n1643_, men_men_n1644_, men_men_n1645_, men_men_n1646_, men_men_n1647_, men_men_n1648_, men_men_n1649_, men_men_n1650_, men_men_n1651_, men_men_n1652_, men_men_n1653_, men_men_n1654_, men_men_n1655_, men_men_n1657_, men_men_n1658_, men_men_n1659_, men_men_n1660_, men_men_n1661_, men_men_n1662_, men_men_n1663_, men_men_n1664_, men_men_n1668_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  ZERO       o00(.Y(ori10));
  ZERO       o01(.Y(ori11));
  ZERO       o02(.Y(ori08));
  ZERO       o03(.Y(ori09));
  ZERO       o04(.Y(ori12));
  ZERO       o05(.Y(ori13));
  ZERO       o06(.Y(ori02));
  ZERO       o07(.Y(ori03));
  ZERO       o08(.Y(ori00));
  ZERO       o09(.Y(ori01));
  ZERO       o10(.Y(ori06));
  ZERO       o11(.Y(ori07));
  ONE        o12(.Y(ori04));
  ZERO       o13(.Y(ori05));
  NO2        m0000(.A(d), .B(c), .Y(mai_mai_n29_));
  AN2        m0001(.A(f), .B(e), .Y(mai_mai_n30_));
  NA3        m0002(.A(mai_mai_n30_), .B(mai_mai_n29_), .C(a), .Y(mai_mai_n31_));
  NOi32      m0003(.An(m), .Bn(l), .C(n), .Y(mai_mai_n32_));
  NOi32      m0004(.An(i), .Bn(g), .C(h), .Y(mai_mai_n33_));
  NA2        m0005(.A(mai_mai_n33_), .B(mai_mai_n32_), .Y(mai_mai_n34_));
  NOi32      m0006(.An(j), .Bn(g), .C(k), .Y(mai_mai_n35_));
  NA2        m0007(.A(mai_mai_n35_), .B(m), .Y(mai_mai_n36_));
  NO2        m0008(.A(mai_mai_n36_), .B(n), .Y(mai_mai_n37_));
  INV        m0009(.A(h), .Y(mai_mai_n38_));
  NAi21      m0010(.An(j), .B(l), .Y(mai_mai_n39_));
  NAi32      m0011(.An(n), .Bn(g), .C(m), .Y(mai_mai_n40_));
  NO3        m0012(.A(mai_mai_n40_), .B(mai_mai_n39_), .C(mai_mai_n38_), .Y(mai_mai_n41_));
  NAi31      m0013(.An(n), .B(m), .C(l), .Y(mai_mai_n42_));
  INV        m0014(.A(i), .Y(mai_mai_n43_));
  AN2        m0015(.A(h), .B(g), .Y(mai_mai_n44_));
  NO2        m0016(.A(mai_mai_n1058_), .B(mai_mai_n42_), .Y(mai_mai_n45_));
  NAi21      m0017(.An(n), .B(m), .Y(mai_mai_n46_));
  NOi32      m0018(.An(k), .Bn(h), .C(l), .Y(mai_mai_n47_));
  NOi32      m0019(.An(k), .Bn(h), .C(g), .Y(mai_mai_n48_));
  AOI210     m0020(.A0(mai_mai_n46_), .A1(mai_mai_n34_), .B0(mai_mai_n31_), .Y(mai_mai_n49_));
  INV        m0021(.A(c), .Y(mai_mai_n50_));
  INV        m0022(.A(d), .Y(mai_mai_n51_));
  NAi21      m0023(.An(i), .B(h), .Y(mai_mai_n52_));
  NA2        m0024(.A(g), .B(f), .Y(mai_mai_n53_));
  NAi21      m0025(.An(i), .B(j), .Y(mai_mai_n54_));
  NAi32      m0026(.An(n), .Bn(k), .C(m), .Y(mai_mai_n55_));
  NO2        m0027(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  NAi31      m0028(.An(l), .B(m), .C(k), .Y(mai_mai_n57_));
  NAi21      m0029(.An(e), .B(h), .Y(mai_mai_n58_));
  NAi41      m0030(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n59_));
  NA2        m0031(.A(mai_mai_n56_), .B(g), .Y(mai_mai_n60_));
  INV        m0032(.A(m), .Y(mai_mai_n61_));
  NA2        m0033(.A(k), .B(mai_mai_n61_), .Y(mai_mai_n62_));
  AN4        m0034(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n63_));
  NA2        m0035(.A(h), .B(mai_mai_n63_), .Y(mai_mai_n64_));
  NAi32      m0036(.An(m), .Bn(k), .C(j), .Y(mai_mai_n65_));
  NOi32      m0037(.An(h), .Bn(g), .C(f), .Y(mai_mai_n66_));
  NA2        m0038(.A(mai_mai_n66_), .B(mai_mai_n63_), .Y(mai_mai_n67_));
  OA220      m0039(.A0(mai_mai_n67_), .A1(mai_mai_n65_), .B0(mai_mai_n64_), .B1(mai_mai_n62_), .Y(mai_mai_n68_));
  NA2        m0040(.A(mai_mai_n68_), .B(mai_mai_n60_), .Y(mai_mai_n69_));
  INV        m0041(.A(n), .Y(mai_mai_n70_));
  INV        m0042(.A(j), .Y(mai_mai_n71_));
  NA3        m0043(.A(m), .B(mai_mai_n71_), .C(g), .Y(mai_mai_n72_));
  NO2        m0044(.A(mai_mai_n72_), .B(f), .Y(mai_mai_n73_));
  NAi32      m0045(.An(g), .Bn(f), .C(h), .Y(mai_mai_n74_));
  NAi31      m0046(.An(j), .B(m), .C(l), .Y(mai_mai_n75_));
  NO2        m0047(.A(mai_mai_n75_), .B(mai_mai_n74_), .Y(mai_mai_n76_));
  NAi31      m0048(.An(k), .B(j), .C(g), .Y(mai_mai_n77_));
  NO2        m0049(.A(mai_mai_n77_), .B(f), .Y(mai_mai_n78_));
  NOi21      m0050(.An(g), .B(i), .Y(mai_mai_n79_));
  AOI220     m0051(.A0(m), .A1(mai_mai_n79_), .B0(m), .B1(g), .Y(mai_mai_n80_));
  NO2        m0052(.A(mai_mai_n80_), .B(f), .Y(mai_mai_n81_));
  NO4        m0053(.A(mai_mai_n81_), .B(mai_mai_n78_), .C(mai_mai_n76_), .D(mai_mai_n73_), .Y(mai_mai_n82_));
  NAi41      m0054(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n83_));
  AN2        m0055(.A(e), .B(b), .Y(mai_mai_n84_));
  NOi31      m0056(.An(c), .B(h), .C(f), .Y(mai_mai_n85_));
  NA2        m0057(.A(mai_mai_n85_), .B(mai_mai_n84_), .Y(mai_mai_n86_));
  NO3        m0058(.A(mai_mai_n86_), .B(mai_mai_n83_), .C(g), .Y(mai_mai_n87_));
  NOi21      m0059(.An(i), .B(h), .Y(mai_mai_n88_));
  NA3        m0060(.A(mai_mai_n88_), .B(g), .C(m), .Y(mai_mai_n89_));
  INV        m0061(.A(l), .Y(mai_mai_n90_));
  NOi21      m0062(.An(m), .B(n), .Y(mai_mai_n91_));
  AN2        m0063(.A(k), .B(h), .Y(mai_mai_n92_));
  NO2        m0064(.A(mai_mai_n89_), .B(n), .Y(mai_mai_n93_));
  INV        m0065(.A(b), .Y(mai_mai_n94_));
  NA2        m0066(.A(l), .B(j), .Y(mai_mai_n95_));
  AN2        m0067(.A(k), .B(i), .Y(mai_mai_n96_));
  NA2        m0068(.A(g), .B(e), .Y(mai_mai_n97_));
  NA2        m0069(.A(c), .B(mai_mai_n91_), .Y(mai_mai_n98_));
  NO3        m0070(.A(mai_mai_n98_), .B(mai_mai_n97_), .C(mai_mai_n94_), .Y(mai_mai_n99_));
  NO3        m0071(.A(mai_mai_n99_), .B(mai_mai_n93_), .C(mai_mai_n87_), .Y(mai_mai_n100_));
  OAI210     m0072(.A0(mai_mai_n82_), .A1(n), .B0(mai_mai_n100_), .Y(mai_mai_n101_));
  NOi31      m0073(.An(k), .B(m), .C(j), .Y(mai_mai_n102_));
  NA3        m0074(.A(mai_mai_n102_), .B(h), .C(mai_mai_n63_), .Y(mai_mai_n103_));
  NOi31      m0075(.An(k), .B(m), .C(i), .Y(mai_mai_n104_));
  NA3        m0076(.A(mai_mai_n104_), .B(mai_mai_n66_), .C(mai_mai_n63_), .Y(mai_mai_n105_));
  NA2        m0077(.A(mai_mai_n105_), .B(mai_mai_n103_), .Y(mai_mai_n106_));
  NAi21      m0078(.An(g), .B(h), .Y(mai_mai_n107_));
  NAi21      m0079(.An(m), .B(n), .Y(mai_mai_n108_));
  NAi21      m0080(.An(j), .B(k), .Y(mai_mai_n109_));
  NO3        m0081(.A(mai_mai_n109_), .B(mai_mai_n108_), .C(mai_mai_n107_), .Y(mai_mai_n110_));
  NAi41      m0082(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n111_));
  NAi31      m0083(.An(j), .B(k), .C(h), .Y(mai_mai_n112_));
  NO3        m0084(.A(mai_mai_n112_), .B(mai_mai_n111_), .C(mai_mai_n108_), .Y(mai_mai_n113_));
  AOI210     m0085(.A0(mai_mai_n110_), .A1(b), .B0(mai_mai_n113_), .Y(mai_mai_n114_));
  NO2        m0086(.A(k), .B(j), .Y(mai_mai_n115_));
  INV        m0087(.A(mai_mai_n108_), .Y(mai_mai_n116_));
  AN2        m0088(.A(k), .B(j), .Y(mai_mai_n117_));
  NAi21      m0089(.An(c), .B(b), .Y(mai_mai_n118_));
  NA2        m0090(.A(f), .B(d), .Y(mai_mai_n119_));
  NO3        m0091(.A(mai_mai_n119_), .B(mai_mai_n118_), .C(mai_mai_n107_), .Y(mai_mai_n120_));
  NA2        m0092(.A(h), .B(c), .Y(mai_mai_n121_));
  NA2        m0093(.A(mai_mai_n120_), .B(mai_mai_n116_), .Y(mai_mai_n122_));
  NA2        m0094(.A(d), .B(b), .Y(mai_mai_n123_));
  NAi21      m0095(.An(e), .B(f), .Y(mai_mai_n124_));
  NO2        m0096(.A(mai_mai_n124_), .B(mai_mai_n123_), .Y(mai_mai_n125_));
  NAi21      m0097(.An(e), .B(g), .Y(mai_mai_n126_));
  NAi21      m0098(.An(c), .B(d), .Y(mai_mai_n127_));
  NAi31      m0099(.An(l), .B(k), .C(h), .Y(mai_mai_n128_));
  NO2        m0100(.A(mai_mai_n108_), .B(mai_mai_n128_), .Y(mai_mai_n129_));
  NA2        m0101(.A(mai_mai_n129_), .B(mai_mai_n125_), .Y(mai_mai_n130_));
  NAi41      m0102(.An(mai_mai_n106_), .B(mai_mai_n130_), .C(mai_mai_n122_), .D(mai_mai_n114_), .Y(mai_mai_n131_));
  NOi21      m0103(.An(h), .B(i), .Y(mai_mai_n132_));
  NOi21      m0104(.An(k), .B(m), .Y(mai_mai_n133_));
  NA3        m0105(.A(mai_mai_n133_), .B(mai_mai_n132_), .C(n), .Y(mai_mai_n134_));
  NOi21      m0106(.An(b), .B(mai_mai_n134_), .Y(mai_mai_n135_));
  NA2        m0107(.A(b), .B(h), .Y(mai_mai_n136_));
  INV        m0108(.A(mai_mai_n46_), .Y(mai_mai_n137_));
  NA2        m0109(.A(mai_mai_n137_), .B(g), .Y(mai_mai_n138_));
  NOi32      m0110(.An(n), .Bn(k), .C(m), .Y(mai_mai_n139_));
  NA2        m0111(.A(l), .B(i), .Y(mai_mai_n140_));
  NA2        m0112(.A(mai_mai_n140_), .B(mai_mai_n139_), .Y(mai_mai_n141_));
  OAI210     m0113(.A0(mai_mai_n141_), .A1(mai_mai_n136_), .B0(mai_mai_n138_), .Y(mai_mai_n142_));
  NA2        m0114(.A(j), .B(h), .Y(mai_mai_n143_));
  OR3        m0115(.A(n), .B(m), .C(k), .Y(mai_mai_n144_));
  NO2        m0116(.A(mai_mai_n144_), .B(mai_mai_n143_), .Y(mai_mai_n145_));
  NAi32      m0117(.An(m), .Bn(k), .C(n), .Y(mai_mai_n146_));
  NO2        m0118(.A(mai_mai_n146_), .B(mai_mai_n143_), .Y(mai_mai_n147_));
  AOI220     m0119(.A0(mai_mai_n147_), .A1(b), .B0(mai_mai_n145_), .B1(c), .Y(mai_mai_n148_));
  NO2        m0120(.A(n), .B(m), .Y(mai_mai_n149_));
  NA2        m0121(.A(mai_mai_n149_), .B(mai_mai_n47_), .Y(mai_mai_n150_));
  NAi21      m0122(.An(f), .B(e), .Y(mai_mai_n151_));
  NA2        m0123(.A(d), .B(c), .Y(mai_mai_n152_));
  NAi31      m0124(.An(m), .B(n), .C(b), .Y(mai_mai_n153_));
  NA2        m0125(.A(k), .B(i), .Y(mai_mai_n154_));
  NAi21      m0126(.An(h), .B(f), .Y(mai_mai_n155_));
  NO2        m0127(.A(mai_mai_n155_), .B(mai_mai_n154_), .Y(mai_mai_n156_));
  NO2        m0128(.A(mai_mai_n153_), .B(mai_mai_n127_), .Y(mai_mai_n157_));
  NA2        m0129(.A(mai_mai_n157_), .B(mai_mai_n156_), .Y(mai_mai_n158_));
  NO2        m0130(.A(c), .B(c), .Y(mai_mai_n159_));
  NO3        m0131(.A(n), .B(m), .C(j), .Y(mai_mai_n160_));
  NA2        m0132(.A(mai_mai_n160_), .B(mai_mai_n92_), .Y(mai_mai_n161_));
  AO210      m0133(.A0(mai_mai_n161_), .A1(mai_mai_n150_), .B0(mai_mai_n159_), .Y(mai_mai_n162_));
  NA3        m0134(.A(mai_mai_n162_), .B(mai_mai_n158_), .C(mai_mai_n148_), .Y(mai_mai_n163_));
  OR4        m0135(.A(mai_mai_n163_), .B(mai_mai_n142_), .C(mai_mai_n135_), .D(mai_mai_n131_), .Y(mai_mai_n164_));
  NO4        m0136(.A(mai_mai_n164_), .B(mai_mai_n101_), .C(mai_mai_n69_), .D(mai_mai_n49_), .Y(mai_mai_n165_));
  NAi31      m0137(.An(n), .B(h), .C(g), .Y(mai_mai_n166_));
  NO2        m0138(.A(mai_mai_n166_), .B(mai_mai_n1051_), .Y(mai_mai_n167_));
  NA3        m0139(.A(m), .B(mai_mai_n71_), .C(g), .Y(mai_mai_n168_));
  NO2        m0140(.A(mai_mai_n168_), .B(n), .Y(mai_mai_n169_));
  NOi21      m0141(.An(k), .B(j), .Y(mai_mai_n170_));
  NA4        m0142(.A(mai_mai_n170_), .B(mai_mai_n91_), .C(i), .D(g), .Y(mai_mai_n171_));
  AN2        m0143(.A(i), .B(g), .Y(mai_mai_n172_));
  NA3        m0144(.A(k), .B(mai_mai_n172_), .C(mai_mai_n91_), .Y(mai_mai_n173_));
  NA2        m0145(.A(mai_mai_n173_), .B(mai_mai_n171_), .Y(mai_mai_n174_));
  INV        m0146(.A(f), .Y(mai_mai_n175_));
  INV        m0147(.A(g), .Y(mai_mai_n176_));
  NOi31      m0148(.An(i), .B(j), .C(h), .Y(mai_mai_n177_));
  NOi21      m0149(.An(l), .B(m), .Y(mai_mai_n178_));
  NA2        m0150(.A(mai_mai_n178_), .B(mai_mai_n177_), .Y(mai_mai_n179_));
  NO3        m0151(.A(mai_mai_n179_), .B(mai_mai_n176_), .C(mai_mai_n175_), .Y(mai_mai_n180_));
  NA2        m0152(.A(mai_mai_n180_), .B(n), .Y(mai_mai_n181_));
  INV        m0153(.A(mai_mai_n181_), .Y(mai_mai_n182_));
  NOi21      m0154(.An(n), .B(m), .Y(mai_mai_n183_));
  NOi32      m0155(.An(l), .Bn(i), .C(j), .Y(mai_mai_n184_));
  NA2        m0156(.A(mai_mai_n184_), .B(mai_mai_n183_), .Y(mai_mai_n185_));
  OA220      m0157(.A0(mai_mai_n185_), .A1(mai_mai_n86_), .B0(mai_mai_n65_), .B1(mai_mai_n64_), .Y(mai_mai_n186_));
  NAi21      m0158(.An(j), .B(h), .Y(mai_mai_n187_));
  NOi31      m0159(.An(k), .B(n), .C(m), .Y(mai_mai_n188_));
  NOi31      m0160(.An(mai_mai_n188_), .B(mai_mai_n152_), .C(mai_mai_n151_), .Y(mai_mai_n189_));
  INV        m0161(.A(mai_mai_n189_), .Y(mai_mai_n190_));
  NAi31      m0162(.An(f), .B(e), .C(c), .Y(mai_mai_n191_));
  NO4        m0163(.A(mai_mai_n191_), .B(mai_mai_n144_), .C(mai_mai_n143_), .D(mai_mai_n51_), .Y(mai_mai_n192_));
  NAi32      m0164(.An(m), .Bn(i), .C(k), .Y(mai_mai_n193_));
  NO3        m0165(.A(mai_mai_n193_), .B(mai_mai_n74_), .C(n), .Y(mai_mai_n194_));
  NA2        m0166(.A(k), .B(h), .Y(mai_mai_n195_));
  NO2        m0167(.A(mai_mai_n194_), .B(mai_mai_n192_), .Y(mai_mai_n196_));
  NAi21      m0168(.An(n), .B(a), .Y(mai_mai_n197_));
  NO2        m0169(.A(mai_mai_n197_), .B(mai_mai_n123_), .Y(mai_mai_n198_));
  NAi41      m0170(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n199_));
  NO2        m0171(.A(mai_mai_n199_), .B(e), .Y(mai_mai_n200_));
  OAI210     m0172(.A0(m), .A1(mai_mai_n200_), .B0(mai_mai_n198_), .Y(mai_mai_n201_));
  AN4        m0173(.A(mai_mai_n201_), .B(mai_mai_n196_), .C(mai_mai_n190_), .D(mai_mai_n186_), .Y(mai_mai_n202_));
  OR2        m0174(.A(h), .B(g), .Y(mai_mai_n203_));
  NO2        m0175(.A(mai_mai_n203_), .B(mai_mai_n83_), .Y(mai_mai_n204_));
  NA2        m0176(.A(mai_mai_n204_), .B(b), .Y(mai_mai_n205_));
  NAi41      m0177(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n206_));
  NO2        m0178(.A(mai_mai_n206_), .B(mai_mai_n175_), .Y(mai_mai_n207_));
  NA2        m0179(.A(mai_mai_n133_), .B(mai_mai_n88_), .Y(mai_mai_n208_));
  NAi21      m0180(.An(mai_mai_n208_), .B(mai_mai_n207_), .Y(mai_mai_n209_));
  NO2        m0181(.A(n), .B(a), .Y(mai_mai_n210_));
  NAi31      m0182(.An(mai_mai_n199_), .B(mai_mai_n210_), .C(mai_mai_n84_), .Y(mai_mai_n211_));
  AN2        m0183(.A(mai_mai_n211_), .B(mai_mai_n209_), .Y(mai_mai_n212_));
  NAi21      m0184(.An(h), .B(i), .Y(mai_mai_n213_));
  NA2        m0185(.A(mai_mai_n149_), .B(k), .Y(mai_mai_n214_));
  NO2        m0186(.A(mai_mai_n214_), .B(mai_mai_n213_), .Y(mai_mai_n215_));
  NA2        m0187(.A(mai_mai_n215_), .B(c), .Y(mai_mai_n216_));
  NA3        m0188(.A(mai_mai_n216_), .B(mai_mai_n212_), .C(mai_mai_n205_), .Y(mai_mai_n217_));
  NOi21      m0189(.An(g), .B(e), .Y(mai_mai_n218_));
  NO2        m0190(.A(mai_mai_n59_), .B(mai_mai_n61_), .Y(mai_mai_n219_));
  NO2        m0191(.A(mai_mai_n55_), .B(mai_mai_n95_), .Y(mai_mai_n220_));
  NOi41      m0192(.An(mai_mai_n202_), .B(mai_mai_n219_), .C(mai_mai_n217_), .D(mai_mai_n182_), .Y(mai_mai_n221_));
  NO4        m0193(.A(mai_mai_n167_), .B(mai_mai_n45_), .C(mai_mai_n41_), .D(mai_mai_n37_), .Y(mai_mai_n222_));
  INV        m0194(.A(mai_mai_n222_), .Y(mai_mai_n223_));
  NAi21      m0195(.An(h), .B(g), .Y(mai_mai_n224_));
  OR3        m0196(.A(mai_mai_n224_), .B(mai_mai_n185_), .C(e), .Y(mai_mai_n225_));
  NO2        m0197(.A(mai_mai_n208_), .B(f), .Y(mai_mai_n226_));
  NA2        m0198(.A(mai_mai_n226_), .B(mai_mai_n63_), .Y(mai_mai_n227_));
  NAi31      m0199(.An(g), .B(k), .C(h), .Y(mai_mai_n228_));
  NO3        m0200(.A(mai_mai_n108_), .B(mai_mai_n228_), .C(l), .Y(mai_mai_n229_));
  NAi31      m0201(.An(e), .B(d), .C(a), .Y(mai_mai_n230_));
  NA2        m0202(.A(mai_mai_n229_), .B(b), .Y(mai_mai_n231_));
  NA3        m0203(.A(mai_mai_n231_), .B(mai_mai_n227_), .C(mai_mai_n225_), .Y(mai_mai_n232_));
  NA4        m0204(.A(mai_mai_n133_), .B(mai_mai_n66_), .C(mai_mai_n63_), .D(mai_mai_n95_), .Y(mai_mai_n233_));
  NA3        m0205(.A(mai_mai_n133_), .B(mai_mai_n132_), .C(mai_mai_n70_), .Y(mai_mai_n234_));
  NO2        m0206(.A(mai_mai_n234_), .B(mai_mai_n159_), .Y(mai_mai_n235_));
  NOi21      m0207(.An(mai_mai_n233_), .B(mai_mai_n235_), .Y(mai_mai_n236_));
  NA3        m0208(.A(e), .B(c), .C(b), .Y(mai_mai_n237_));
  INV        m0209(.A(mai_mai_n46_), .Y(mai_mai_n238_));
  NA2        m0210(.A(g), .B(mai_mai_n238_), .Y(mai_mai_n239_));
  NAi21      m0211(.An(l), .B(k), .Y(mai_mai_n240_));
  NO2        m0212(.A(mai_mai_n240_), .B(mai_mai_n46_), .Y(mai_mai_n241_));
  NA2        m0213(.A(h), .B(l), .Y(mai_mai_n242_));
  NO2        m0214(.A(mai_mai_n242_), .B(mai_mai_n59_), .Y(mai_mai_n243_));
  INV        m0215(.A(mai_mai_n243_), .Y(mai_mai_n244_));
  NAi32      m0216(.An(j), .Bn(h), .C(i), .Y(mai_mai_n245_));
  NAi21      m0217(.An(m), .B(l), .Y(mai_mai_n246_));
  NO3        m0218(.A(mai_mai_n246_), .B(mai_mai_n245_), .C(mai_mai_n70_), .Y(mai_mai_n247_));
  NA2        m0219(.A(h), .B(g), .Y(mai_mai_n248_));
  NA2        m0220(.A(mai_mai_n247_), .B(b), .Y(mai_mai_n249_));
  NA4        m0221(.A(mai_mai_n249_), .B(mai_mai_n244_), .C(mai_mai_n239_), .D(mai_mai_n236_), .Y(mai_mai_n250_));
  NO2        m0222(.A(f), .B(d), .Y(mai_mai_n251_));
  NO2        m0223(.A(mai_mai_n86_), .B(mai_mai_n83_), .Y(mai_mai_n252_));
  NAi32      m0224(.An(n), .Bn(m), .C(l), .Y(mai_mai_n253_));
  NO2        m0225(.A(mai_mai_n253_), .B(mai_mai_n245_), .Y(mai_mai_n254_));
  NA2        m0226(.A(mai_mai_n252_), .B(mai_mai_n51_), .Y(mai_mai_n255_));
  NO4        m0227(.A(mai_mai_n252_), .B(mai_mai_n250_), .C(mai_mai_n232_), .D(mai_mai_n223_), .Y(mai_mai_n256_));
  NA2        m0228(.A(mai_mai_n215_), .B(c), .Y(mai_mai_n257_));
  NAi21      m0229(.An(m), .B(k), .Y(mai_mai_n258_));
  INV        m0230(.A(mai_mai_n258_), .Y(mai_mai_n259_));
  NAi41      m0231(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n260_));
  NO2        m0232(.A(mai_mai_n260_), .B(mai_mai_n126_), .Y(mai_mai_n261_));
  NA2        m0233(.A(mai_mai_n261_), .B(mai_mai_n259_), .Y(mai_mai_n262_));
  NO4        m0234(.A(i), .B(mai_mai_n126_), .C(mai_mai_n59_), .D(mai_mai_n61_), .Y(mai_mai_n263_));
  NAi31      m0235(.An(d), .B(e), .C(b), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n108_), .B(mai_mai_n264_), .Y(mai_mai_n265_));
  NA2        m0237(.A(mai_mai_n265_), .B(mai_mai_n96_), .Y(mai_mai_n266_));
  NAi41      m0238(.An(mai_mai_n263_), .B(mai_mai_n266_), .C(mai_mai_n262_), .D(mai_mai_n257_), .Y(mai_mai_n267_));
  NO4        m0239(.A(mai_mai_n260_), .B(mai_mai_n65_), .C(mai_mai_n58_), .D(mai_mai_n176_), .Y(mai_mai_n268_));
  OR2        m0240(.A(n), .B(mai_mai_n168_), .Y(mai_mai_n269_));
  NOi31      m0241(.An(l), .B(n), .C(m), .Y(mai_mai_n270_));
  NA2        m0242(.A(mai_mai_n270_), .B(mai_mai_n177_), .Y(mai_mai_n271_));
  NO2        m0243(.A(mai_mai_n271_), .B(mai_mai_n159_), .Y(mai_mai_n272_));
  NAi32      m0244(.An(mai_mai_n272_), .Bn(mai_mai_n268_), .C(mai_mai_n269_), .Y(mai_mai_n273_));
  NAi32      m0245(.An(m), .Bn(j), .C(k), .Y(mai_mai_n274_));
  NAi41      m0246(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n275_));
  NOi31      m0247(.An(j), .B(m), .C(k), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n102_), .B(mai_mai_n276_), .Y(mai_mai_n277_));
  AN3        m0249(.A(h), .B(g), .C(f), .Y(mai_mai_n278_));
  NAi31      m0250(.An(mai_mai_n277_), .B(mai_mai_n278_), .C(b), .Y(mai_mai_n279_));
  OR2        m0251(.A(mai_mai_n1050_), .B(mai_mai_n166_), .Y(mai_mai_n280_));
  NO2        m0252(.A(mai_mai_n246_), .B(mai_mai_n245_), .Y(mai_mai_n281_));
  NO2        m0253(.A(mai_mai_n179_), .B(g), .Y(mai_mai_n282_));
  AOI220     m0254(.A0(b), .A1(mai_mai_n282_), .B0(mai_mai_n207_), .B1(mai_mai_n281_), .Y(mai_mai_n283_));
  NA3        m0255(.A(mai_mai_n283_), .B(mai_mai_n280_), .C(mai_mai_n279_), .Y(mai_mai_n284_));
  NA3        m0256(.A(h), .B(g), .C(f), .Y(mai_mai_n285_));
  NO2        m0257(.A(mai_mai_n285_), .B(mai_mai_n62_), .Y(mai_mai_n286_));
  NA2        m0258(.A(h), .B(e), .Y(mai_mai_n287_));
  AOI220     m0259(.A0(h), .A1(mai_mai_n91_), .B0(b), .B1(mai_mai_n286_), .Y(mai_mai_n288_));
  NA3        m0260(.A(g), .B(mai_mai_n240_), .C(mai_mai_n91_), .Y(mai_mai_n289_));
  BUFFER     m0261(.A(mai_mai_n289_), .Y(mai_mai_n290_));
  AN2        m0262(.A(l), .B(j), .Y(mai_mai_n291_));
  INV        m0263(.A(mai_mai_n258_), .Y(mai_mai_n292_));
  NO3        m0264(.A(mai_mai_n260_), .B(mai_mai_n58_), .C(mai_mai_n176_), .Y(mai_mai_n293_));
  NA3        m0265(.A(mai_mai_n173_), .B(mai_mai_n171_), .C(mai_mai_n34_), .Y(mai_mai_n294_));
  AOI220     m0266(.A0(mai_mai_n294_), .A1(b), .B0(mai_mai_n293_), .B1(mai_mai_n292_), .Y(mai_mai_n295_));
  NA4        m0267(.A(m), .B(mai_mai_n71_), .C(g), .D(mai_mai_n175_), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n48_), .B(mai_mai_n91_), .Y(mai_mai_n297_));
  NO2        m0269(.A(mai_mai_n297_), .B(d), .Y(mai_mai_n298_));
  NA2        m0270(.A(mai_mai_n298_), .B(b), .Y(mai_mai_n299_));
  NA4        m0271(.A(mai_mai_n299_), .B(mai_mai_n295_), .C(mai_mai_n290_), .D(mai_mai_n288_), .Y(mai_mai_n300_));
  NO4        m0272(.A(mai_mai_n300_), .B(mai_mai_n284_), .C(mai_mai_n273_), .D(mai_mai_n267_), .Y(mai_mai_n301_));
  NA4        m0273(.A(mai_mai_n301_), .B(mai_mai_n256_), .C(mai_mai_n221_), .D(mai_mai_n165_), .Y(mai10));
  NA3        m0274(.A(m), .B(k), .C(i), .Y(mai_mai_n303_));
  NOi32      m0275(.An(k), .Bn(h), .C(j), .Y(mai_mai_n304_));
  NA2        m0276(.A(mai_mai_n304_), .B(mai_mai_n183_), .Y(mai_mai_n305_));
  NA2        m0277(.A(mai_mai_n134_), .B(mai_mai_n305_), .Y(mai_mai_n306_));
  NA2        m0278(.A(mai_mai_n306_), .B(c), .Y(mai_mai_n307_));
  AN2        m0279(.A(j), .B(h), .Y(mai_mai_n308_));
  NO3        m0280(.A(n), .B(m), .C(k), .Y(mai_mai_n309_));
  NA2        m0281(.A(mai_mai_n309_), .B(mai_mai_n308_), .Y(mai_mai_n310_));
  NO3        m0282(.A(mai_mai_n310_), .B(mai_mai_n127_), .C(mai_mai_n175_), .Y(mai_mai_n311_));
  OR2        m0283(.A(m), .B(k), .Y(mai_mai_n312_));
  NO2        m0284(.A(mai_mai_n143_), .B(mai_mai_n312_), .Y(mai_mai_n313_));
  NA4        m0285(.A(n), .B(f), .C(c), .D(mai_mai_n94_), .Y(mai_mai_n314_));
  NOi21      m0286(.An(mai_mai_n313_), .B(mai_mai_n314_), .Y(mai_mai_n315_));
  NAi21      m0287(.An(i), .B(g), .Y(mai_mai_n316_));
  NAi31      m0288(.An(k), .B(m), .C(j), .Y(mai_mai_n317_));
  NO3        m0289(.A(mai_mai_n317_), .B(mai_mai_n316_), .C(n), .Y(mai_mai_n318_));
  BUFFER     m0290(.A(mai_mai_n318_), .Y(mai_mai_n319_));
  NO3        m0291(.A(mai_mai_n319_), .B(mai_mai_n315_), .C(mai_mai_n311_), .Y(mai_mai_n320_));
  NO2        m0292(.A(mai_mai_n314_), .B(mai_mai_n246_), .Y(mai_mai_n321_));
  AOI220     m0293(.A0(d), .A1(mai_mai_n254_), .B0(mai_mai_n321_), .B1(mai_mai_n177_), .Y(mai_mai_n322_));
  NA3        m0294(.A(mai_mai_n322_), .B(mai_mai_n320_), .C(mai_mai_n307_), .Y(mai_mai_n323_));
  INV        m0295(.A(mai_mai_n168_), .Y(mai_mai_n324_));
  AN2        m0296(.A(g), .B(e), .Y(mai_mai_n325_));
  NA3        m0297(.A(mai_mai_n325_), .B(m), .C(i), .Y(mai_mai_n326_));
  NA2        m0298(.A(mai_mai_n72_), .B(mai_mai_n326_), .Y(mai_mai_n327_));
  INV        m0299(.A(mai_mai_n80_), .Y(mai_mai_n328_));
  NO3        m0300(.A(mai_mai_n328_), .B(mai_mai_n327_), .C(mai_mai_n324_), .Y(mai_mai_n329_));
  NOi32      m0301(.An(h), .Bn(e), .C(g), .Y(mai_mai_n330_));
  NA2        m0302(.A(mai_mai_n330_), .B(m), .Y(mai_mai_n331_));
  NA3        m0303(.A(m), .B(h), .C(e), .Y(mai_mai_n332_));
  AN3        m0304(.A(h), .B(g), .C(e), .Y(mai_mai_n333_));
  NA2        m0305(.A(mai_mai_n333_), .B(m), .Y(mai_mai_n334_));
  AN3        m0306(.A(mai_mai_n334_), .B(mai_mai_n332_), .C(mai_mai_n331_), .Y(mai_mai_n335_));
  AOI210     m0307(.A0(mai_mai_n335_), .A1(mai_mai_n329_), .B0(n), .Y(mai_mai_n336_));
  NA3        m0308(.A(mai_mai_n35_), .B(m), .C(e), .Y(mai_mai_n337_));
  NO2        m0309(.A(mai_mai_n337_), .B(n), .Y(mai_mai_n338_));
  NO2        m0310(.A(b), .B(n), .Y(mai_mai_n339_));
  OAI210     m0311(.A0(mai_mai_n48_), .A1(mai_mai_n47_), .B0(m), .Y(mai_mai_n340_));
  NO2        m0312(.A(mai_mai_n340_), .B(mai_mai_n124_), .Y(mai_mai_n341_));
  NA2        m0313(.A(mai_mai_n341_), .B(mai_mai_n339_), .Y(mai_mai_n342_));
  INV        m0314(.A(mai_mai_n342_), .Y(mai_mai_n343_));
  NO4        m0315(.A(mai_mai_n343_), .B(mai_mai_n338_), .C(mai_mai_n336_), .D(mai_mai_n323_), .Y(mai_mai_n344_));
  NO3        m0316(.A(mai_mai_n230_), .B(i), .C(c), .Y(mai_mai_n345_));
  NOi21      m0317(.An(a), .B(n), .Y(mai_mai_n346_));
  NA3        m0318(.A(i), .B(g), .C(f), .Y(mai_mai_n347_));
  OR2        m0319(.A(mai_mai_n347_), .B(mai_mai_n57_), .Y(mai_mai_n348_));
  NA3        m0320(.A(m), .B(h), .C(mai_mai_n151_), .Y(mai_mai_n349_));
  AOI210     m0321(.A0(mai_mai_n349_), .A1(mai_mai_n348_), .B0(n), .Y(mai_mai_n350_));
  AOI210     m0322(.A0(mai_mai_n345_), .A1(mai_mai_n241_), .B0(mai_mai_n350_), .Y(mai_mai_n351_));
  OR2        m0323(.A(n), .B(m), .Y(mai_mai_n352_));
  NO2        m0324(.A(mai_mai_n352_), .B(mai_mai_n128_), .Y(mai_mai_n353_));
  OAI210     m0325(.A0(mai_mai_n353_), .A1(mai_mai_n145_), .B0(d), .Y(mai_mai_n354_));
  INV        m0326(.A(mai_mai_n46_), .Y(mai_mai_n355_));
  NAi21      m0327(.An(k), .B(j), .Y(mai_mai_n356_));
  NA3        m0328(.A(i), .B(g), .C(mai_mai_n355_), .Y(mai_mai_n357_));
  NAi21      m0329(.An(e), .B(d), .Y(mai_mai_n358_));
  NO2        m0330(.A(mai_mai_n358_), .B(mai_mai_n50_), .Y(mai_mai_n359_));
  NO2        m0331(.A(mai_mai_n214_), .B(mai_mai_n175_), .Y(mai_mai_n360_));
  NA2        m0332(.A(mai_mai_n360_), .B(mai_mai_n359_), .Y(mai_mai_n361_));
  NA4        m0333(.A(mai_mai_n361_), .B(mai_mai_n357_), .C(mai_mai_n297_), .D(mai_mai_n354_), .Y(mai_mai_n362_));
  NO2        m0334(.A(mai_mai_n271_), .B(mai_mai_n175_), .Y(mai_mai_n363_));
  NA2        m0335(.A(mai_mai_n363_), .B(mai_mai_n359_), .Y(mai_mai_n364_));
  NOi31      m0336(.An(n), .B(m), .C(k), .Y(mai_mai_n365_));
  AOI220     m0337(.A0(mai_mai_n365_), .A1(mai_mai_n308_), .B0(mai_mai_n183_), .B1(mai_mai_n47_), .Y(mai_mai_n366_));
  NAi31      m0338(.An(g), .B(f), .C(c), .Y(mai_mai_n367_));
  OR3        m0339(.A(mai_mai_n367_), .B(mai_mai_n366_), .C(e), .Y(mai_mai_n368_));
  NA3        m0340(.A(mai_mai_n368_), .B(mai_mai_n364_), .C(mai_mai_n255_), .Y(mai_mai_n369_));
  NOi41      m0341(.An(mai_mai_n351_), .B(mai_mai_n369_), .C(mai_mai_n362_), .D(mai_mai_n219_), .Y(mai_mai_n370_));
  NA2        m0342(.A(a), .B(mai_mai_n91_), .Y(mai_mai_n371_));
  AN2        m0343(.A(e), .B(d), .Y(mai_mai_n372_));
  NO2        m0344(.A(mai_mai_n53_), .B(e), .Y(mai_mai_n373_));
  AOI210     m0345(.A0(h), .A1(f), .B0(mai_mai_n373_), .Y(mai_mai_n374_));
  AOI210     m0346(.A0(mai_mai_n374_), .A1(mai_mai_n228_), .B0(mai_mai_n371_), .Y(mai_mai_n375_));
  NO2        m0347(.A(mai_mai_n174_), .B(mai_mai_n169_), .Y(mai_mai_n376_));
  NO2        m0348(.A(n), .B(mai_mai_n168_), .Y(mai_mai_n377_));
  NA2        m0349(.A(mai_mai_n222_), .B(mai_mai_n376_), .Y(mai_mai_n378_));
  NO4        m0350(.A(mai_mai_n155_), .B(mai_mai_n83_), .C(mai_mai_n50_), .D(b), .Y(mai_mai_n379_));
  NA2        m0351(.A(c), .B(mai_mai_n129_), .Y(mai_mai_n380_));
  NA2        m0352(.A(l), .B(k), .Y(mai_mai_n381_));
  AOI210     m0353(.A0(mai_mai_n193_), .A1(mai_mai_n274_), .B0(mai_mai_n70_), .Y(mai_mai_n382_));
  OR3        m0354(.A(mai_mai_n1055_), .B(mai_mai_n121_), .C(mai_mai_n111_), .Y(mai_mai_n383_));
  NA3        m0355(.A(mai_mai_n233_), .B(mai_mai_n105_), .C(mai_mai_n103_), .Y(mai_mai_n384_));
  NO4        m0356(.A(n), .B(mai_mai_n77_), .C(mai_mai_n90_), .D(e), .Y(mai_mai_n385_));
  NO3        m0357(.A(n), .B(mai_mai_n75_), .C(mai_mai_n107_), .Y(mai_mai_n386_));
  NO4        m0358(.A(mai_mai_n386_), .B(mai_mai_n385_), .C(mai_mai_n384_), .D(mai_mai_n263_), .Y(mai_mai_n387_));
  NA3        m0359(.A(mai_mai_n387_), .B(mai_mai_n383_), .C(mai_mai_n380_), .Y(mai_mai_n388_));
  NO4        m0360(.A(mai_mai_n388_), .B(mai_mai_n379_), .C(mai_mai_n378_), .D(mai_mai_n375_), .Y(mai_mai_n389_));
  NA2        m0361(.A(mai_mai_n56_), .B(g), .Y(mai_mai_n390_));
  NO2        m0362(.A(mai_mai_n155_), .B(mai_mai_n50_), .Y(mai_mai_n391_));
  NAi31      m0363(.An(j), .B(l), .C(i), .Y(mai_mai_n392_));
  OAI210     m0364(.A0(mai_mai_n392_), .A1(mai_mai_n108_), .B0(mai_mai_n83_), .Y(mai_mai_n393_));
  NA3        m0365(.A(mai_mai_n393_), .B(mai_mai_n391_), .C(b), .Y(mai_mai_n394_));
  NO2        m0366(.A(mai_mai_n1050_), .B(mai_mai_n166_), .Y(mai_mai_n395_));
  INV        m0367(.A(mai_mai_n297_), .Y(mai_mai_n396_));
  NO3        m0368(.A(mai_mai_n396_), .B(mai_mai_n395_), .C(mai_mai_n252_), .Y(mai_mai_n397_));
  NA4        m0369(.A(mai_mai_n397_), .B(mai_mai_n394_), .C(mai_mai_n390_), .D(mai_mai_n202_), .Y(mai_mai_n398_));
  OAI210     m0370(.A0(mai_mai_n104_), .A1(mai_mai_n102_), .B0(n), .Y(mai_mai_n399_));
  NO2        m0371(.A(mai_mai_n399_), .B(mai_mai_n107_), .Y(mai_mai_n400_));
  AO210      m0372(.A0(mai_mai_n247_), .A1(mai_mai_n176_), .B0(mai_mai_n204_), .Y(mai_mai_n401_));
  OA210      m0373(.A0(mai_mai_n401_), .A1(mai_mai_n400_), .B0(c), .Y(mai_mai_n402_));
  XO2        m0374(.A(i), .B(h), .Y(mai_mai_n403_));
  NA3        m0375(.A(mai_mai_n403_), .B(mai_mai_n133_), .C(n), .Y(mai_mai_n404_));
  NAi41      m0376(.An(mai_mai_n247_), .B(mai_mai_n404_), .C(mai_mai_n366_), .D(mai_mai_n305_), .Y(mai_mai_n405_));
  AN2        m0377(.A(mai_mai_n405_), .B(mai_mai_n373_), .Y(mai_mai_n406_));
  AOI210     m0378(.A0(mai_mai_n234_), .A1(mai_mai_n161_), .B0(c), .Y(mai_mai_n407_));
  NOi21      m0379(.An(mai_mai_n68_), .B(mai_mai_n407_), .Y(mai_mai_n408_));
  NA3        m0380(.A(mai_mai_n1061_), .B(m), .C(g), .Y(mai_mai_n409_));
  NA2        m0381(.A(mai_mai_n188_), .B(mai_mai_n88_), .Y(mai_mai_n410_));
  AOI210     m0382(.A0(mai_mai_n410_), .A1(mai_mai_n150_), .B0(c), .Y(mai_mai_n411_));
  NA2        m0383(.A(mai_mai_n289_), .B(mai_mai_n34_), .Y(mai_mai_n412_));
  NOi31      m0384(.An(mai_mai_n409_), .B(mai_mai_n412_), .C(mai_mai_n411_), .Y(mai_mai_n413_));
  AO220      m0385(.A0(mai_mai_n238_), .A1(g), .B0(mai_mai_n137_), .B1(g), .Y(mai_mai_n414_));
  NA3        m0386(.A(mai_mai_n35_), .B(m), .C(f), .Y(mai_mai_n415_));
  NO2        m0387(.A(mai_mai_n415_), .B(n), .Y(mai_mai_n416_));
  NO2        m0388(.A(mai_mai_n416_), .B(mai_mai_n243_), .Y(mai_mai_n417_));
  NAi41      m0389(.An(mai_mai_n414_), .B(mai_mai_n417_), .C(mai_mai_n413_), .D(mai_mai_n408_), .Y(mai_mai_n418_));
  NO4        m0390(.A(mai_mai_n418_), .B(mai_mai_n406_), .C(mai_mai_n402_), .D(mai_mai_n398_), .Y(mai_mai_n419_));
  NA4        m0391(.A(mai_mai_n419_), .B(mai_mai_n389_), .C(mai_mai_n370_), .D(mai_mai_n344_), .Y(mai11));
  NA2        m0392(.A(j), .B(g), .Y(mai_mai_n421_));
  NAi31      m0393(.An(i), .B(m), .C(l), .Y(mai_mai_n422_));
  NA3        m0394(.A(m), .B(k), .C(j), .Y(mai_mai_n423_));
  OAI220     m0395(.A0(mai_mai_n423_), .A1(mai_mai_n107_), .B0(mai_mai_n422_), .B1(mai_mai_n421_), .Y(mai_mai_n424_));
  NOi32      m0396(.An(e), .Bn(b), .C(f), .Y(mai_mai_n425_));
  NA2        m0397(.A(j), .B(mai_mai_n91_), .Y(mai_mai_n426_));
  NA2        m0398(.A(mai_mai_n44_), .B(j), .Y(mai_mai_n427_));
  OAI220     m0399(.A0(mai_mai_n427_), .A1(n), .B0(mai_mai_n426_), .B1(mai_mai_n176_), .Y(mai_mai_n428_));
  NAi31      m0400(.An(d), .B(e), .C(a), .Y(mai_mai_n429_));
  NO2        m0401(.A(mai_mai_n429_), .B(n), .Y(mai_mai_n430_));
  AOI220     m0402(.A0(mai_mai_n430_), .A1(mai_mai_n81_), .B0(mai_mai_n428_), .B1(mai_mai_n425_), .Y(mai_mai_n431_));
  NA2        m0403(.A(j), .B(i), .Y(mai_mai_n432_));
  NAi31      m0404(.An(n), .B(m), .C(k), .Y(mai_mai_n433_));
  NO3        m0405(.A(mai_mai_n433_), .B(mai_mai_n432_), .C(mai_mai_n90_), .Y(mai_mai_n434_));
  OR2        m0406(.A(n), .B(c), .Y(mai_mai_n435_));
  INV        m0407(.A(mai_mai_n435_), .Y(mai_mai_n436_));
  NOi32      m0408(.An(g), .Bn(f), .C(i), .Y(mai_mai_n437_));
  AOI220     m0409(.A0(mai_mai_n437_), .A1(m), .B0(mai_mai_n424_), .B1(f), .Y(mai_mai_n438_));
  NO2        m0410(.A(mai_mai_n228_), .B(mai_mai_n46_), .Y(mai_mai_n439_));
  NO2        m0411(.A(mai_mai_n438_), .B(n), .Y(mai_mai_n440_));
  AOI210     m0412(.A0(mai_mai_n434_), .A1(g), .B0(mai_mai_n440_), .Y(mai_mai_n441_));
  NA2        m0413(.A(mai_mai_n117_), .B(mai_mai_n33_), .Y(mai_mai_n442_));
  OAI220     m0414(.A0(mai_mai_n442_), .A1(m), .B0(mai_mai_n427_), .B1(mai_mai_n193_), .Y(mai_mai_n443_));
  NAi32      m0415(.An(e), .Bn(b), .C(c), .Y(mai_mai_n444_));
  OAI220     m0416(.A0(mai_mai_n317_), .A1(mai_mai_n316_), .B0(mai_mai_n422_), .B1(mai_mai_n421_), .Y(mai_mai_n445_));
  NO2        m0417(.A(d), .B(n), .Y(mai_mai_n446_));
  NA3        m0418(.A(mai_mai_n446_), .B(mai_mai_n445_), .C(e), .Y(mai_mai_n447_));
  NO3        m0419(.A(i), .B(mai_mai_n46_), .C(mai_mai_n176_), .Y(mai_mai_n448_));
  OAI210     m0420(.A0(mai_mai_n448_), .A1(mai_mai_n318_), .B0(a), .Y(mai_mai_n449_));
  NA2        m0421(.A(mai_mai_n449_), .B(mai_mai_n447_), .Y(mai_mai_n450_));
  NA2        m0422(.A(mai_mai_n445_), .B(f), .Y(mai_mai_n451_));
  NO2        m0423(.A(d), .B(mai_mai_n46_), .Y(mai_mai_n452_));
  NO3        m0424(.A(mai_mai_n146_), .B(mai_mai_n143_), .C(g), .Y(mai_mai_n453_));
  AOI220     m0425(.A0(mai_mai_n453_), .A1(c), .B0(g), .B1(mai_mai_n452_), .Y(mai_mai_n454_));
  OAI210     m0426(.A0(mai_mai_n451_), .A1(n), .B0(mai_mai_n454_), .Y(mai_mai_n455_));
  NO2        m0427(.A(mai_mai_n123_), .B(c), .Y(mai_mai_n456_));
  NA3        m0428(.A(mai_mai_n456_), .B(h), .C(mai_mai_n365_), .Y(mai_mai_n457_));
  NA3        m0429(.A(f), .B(d), .C(b), .Y(mai_mai_n458_));
  NO4        m0430(.A(mai_mai_n458_), .B(mai_mai_n146_), .C(mai_mai_n143_), .D(g), .Y(mai_mai_n459_));
  NAi21      m0431(.An(mai_mai_n459_), .B(mai_mai_n457_), .Y(mai_mai_n460_));
  NO4        m0432(.A(mai_mai_n460_), .B(mai_mai_n455_), .C(mai_mai_n450_), .D(mai_mai_n443_), .Y(mai_mai_n461_));
  AN3        m0433(.A(mai_mai_n461_), .B(mai_mai_n441_), .C(mai_mai_n431_), .Y(mai_mai_n462_));
  INV        m0434(.A(k), .Y(mai_mai_n463_));
  NA4        m0435(.A(a), .B(h), .C(mai_mai_n151_), .D(mai_mai_n91_), .Y(mai_mai_n464_));
  NAi31      m0436(.An(h), .B(g), .C(f), .Y(mai_mai_n465_));
  OR3        m0437(.A(mai_mai_n465_), .B(mai_mai_n230_), .C(mai_mai_n46_), .Y(mai_mai_n466_));
  NA4        m0438(.A(h), .B(c), .C(mai_mai_n91_), .D(e), .Y(mai_mai_n467_));
  AN2        m0439(.A(mai_mai_n467_), .B(mai_mai_n466_), .Y(mai_mai_n468_));
  NO2        m0440(.A(mai_mai_n59_), .B(mai_mai_n61_), .Y(mai_mai_n469_));
  NO3        m0441(.A(mai_mai_n465_), .B(mai_mai_n435_), .C(mai_mai_n61_), .Y(mai_mai_n470_));
  OR2        m0442(.A(mai_mai_n470_), .B(mai_mai_n469_), .Y(mai_mai_n471_));
  NAi31      m0443(.An(mai_mai_n471_), .B(mai_mai_n468_), .C(mai_mai_n464_), .Y(mai_mai_n472_));
  NAi31      m0444(.An(f), .B(h), .C(g), .Y(mai_mai_n473_));
  NO4        m0445(.A(k), .B(mai_mai_n473_), .C(mai_mai_n59_), .D(mai_mai_n61_), .Y(mai_mai_n474_));
  NOi41      m0446(.An(b), .B(mai_mai_n285_), .C(mai_mai_n55_), .D(mai_mai_n95_), .Y(mai_mai_n475_));
  OR2        m0447(.A(mai_mai_n475_), .B(mai_mai_n474_), .Y(mai_mai_n476_));
  NO2        m0448(.A(n), .B(c), .Y(mai_mai_n477_));
  NA3        m0449(.A(mai_mai_n477_), .B(a), .C(m), .Y(mai_mai_n478_));
  AOI210     m0450(.A0(mai_mai_n33_), .A1(mai_mai_n91_), .B0(mai_mai_n476_), .Y(mai_mai_n479_));
  OAI210     m0451(.A0(mai_mai_n209_), .A1(mai_mai_n71_), .B0(mai_mai_n479_), .Y(mai_mai_n480_));
  NO2        m0452(.A(mai_mai_n472_), .B(mai_mai_n480_), .Y(mai_mai_n481_));
  NO3        m0453(.A(mai_mai_n258_), .B(mai_mai_n52_), .C(n), .Y(mai_mai_n482_));
  NA2        m0454(.A(k), .B(mai_mai_n91_), .Y(mai_mai_n483_));
  AOI210     m0455(.A0(mai_mai_n91_), .A1(g), .B0(mai_mai_n482_), .Y(mai_mai_n484_));
  NO2        m0456(.A(mai_mai_n484_), .B(mai_mai_n71_), .Y(mai_mai_n485_));
  NA3        m0457(.A(d), .B(mai_mai_n276_), .C(mai_mai_n44_), .Y(mai_mai_n486_));
  AOI220     m0458(.A0(e), .A1(mai_mai_n313_), .B0(e), .B1(mai_mai_n145_), .Y(mai_mai_n487_));
  NA2        m0459(.A(g), .B(mai_mai_n220_), .Y(mai_mai_n488_));
  NAi21      m0460(.An(k), .B(h), .Y(mai_mai_n489_));
  NOi31      m0461(.An(m), .B(n), .C(k), .Y(mai_mai_n490_));
  NA2        m0462(.A(j), .B(mai_mai_n490_), .Y(mai_mai_n491_));
  NAi21      m0463(.An(mai_mai_n491_), .B(g), .Y(mai_mai_n492_));
  NO2        m0464(.A(mai_mai_n230_), .B(mai_mai_n46_), .Y(mai_mai_n493_));
  INV        m0465(.A(mai_mai_n46_), .Y(mai_mai_n494_));
  AOI220     m0466(.A0(mai_mai_n494_), .A1(g), .B0(mai_mai_n493_), .B1(g), .Y(mai_mai_n495_));
  NA3        m0467(.A(mai_mai_n495_), .B(mai_mai_n492_), .C(mai_mai_n488_), .Y(mai_mai_n496_));
  NO2        m0468(.A(k), .B(mai_mai_n176_), .Y(mai_mai_n497_));
  INV        m0469(.A(n), .Y(mai_mai_n498_));
  NAi31      m0470(.An(mai_mai_n1057_), .B(mai_mai_n498_), .C(mai_mai_n497_), .Y(mai_mai_n499_));
  NO2        m0471(.A(mai_mai_n427_), .B(mai_mai_n146_), .Y(mai_mai_n500_));
  NA2        m0472(.A(mai_mai_n403_), .B(mai_mai_n133_), .Y(mai_mai_n501_));
  NO3        m0473(.A(mai_mai_n314_), .B(mai_mai_n501_), .C(mai_mai_n71_), .Y(mai_mai_n502_));
  AOI210     m0474(.A0(c), .A1(mai_mai_n500_), .B0(mai_mai_n502_), .Y(mai_mai_n503_));
  NA3        m0475(.A(mai_mai_n403_), .B(mai_mai_n133_), .C(mai_mai_n176_), .Y(mai_mai_n504_));
  INV        m0476(.A(mai_mai_n504_), .Y(mai_mai_n505_));
  NAi31      m0477(.An(m), .B(n), .C(k), .Y(mai_mai_n506_));
  OAI210     m0478(.A0(mai_mai_n111_), .A1(mai_mai_n506_), .B0(mai_mai_n211_), .Y(mai_mai_n507_));
  OAI210     m0479(.A0(mai_mai_n507_), .A1(mai_mai_n505_), .B0(j), .Y(mai_mai_n508_));
  NA3        m0480(.A(mai_mai_n508_), .B(mai_mai_n503_), .C(mai_mai_n499_), .Y(mai_mai_n509_));
  NO4        m0481(.A(mai_mai_n509_), .B(mai_mai_n496_), .C(mai_mai_n313_), .D(mai_mai_n485_), .Y(mai_mai_n510_));
  NA2        m0482(.A(mai_mai_n1061_), .B(h), .Y(mai_mai_n511_));
  NAi31      m0483(.An(g), .B(h), .C(f), .Y(mai_mai_n512_));
  OR3        m0484(.A(mai_mai_n512_), .B(mai_mai_n230_), .C(n), .Y(mai_mai_n513_));
  NA3        m0485(.A(mai_mai_n330_), .B(c), .C(mai_mai_n70_), .Y(mai_mai_n514_));
  OAI210     m0486(.A0(n), .A1(mai_mai_n74_), .B0(mai_mai_n514_), .Y(mai_mai_n515_));
  NOi21      m0487(.An(mai_mai_n513_), .B(mai_mai_n515_), .Y(mai_mai_n516_));
  AOI210     m0488(.A0(mai_mai_n516_), .A1(mai_mai_n511_), .B0(mai_mai_n423_), .Y(mai_mai_n517_));
  NAi21      m0489(.An(h), .B(j), .Y(mai_mai_n518_));
  OAI220     m0490(.A0(mai_mai_n518_), .A1(mai_mai_n83_), .B0(mai_mai_n410_), .B1(mai_mai_n71_), .Y(mai_mai_n519_));
  OAI210     m0491(.A0(mai_mai_n519_), .A1(mai_mai_n313_), .B0(c), .Y(mai_mai_n520_));
  OR2        m0492(.A(mai_mai_n489_), .B(mai_mai_n59_), .Y(mai_mai_n521_));
  NA2        m0493(.A(h), .B(mai_mai_n35_), .Y(mai_mai_n522_));
  NA2        m0494(.A(m), .B(mai_mai_n44_), .Y(mai_mai_n523_));
  OAI220     m0495(.A0(mai_mai_n523_), .A1(n), .B0(mai_mai_n522_), .B1(mai_mai_n371_), .Y(mai_mai_n524_));
  INV        m0496(.A(mai_mai_n46_), .Y(mai_mai_n525_));
  AOI210     m0497(.A0(g), .A1(mai_mai_n525_), .B0(mai_mai_n524_), .Y(mai_mai_n526_));
  NA3        m0498(.A(mai_mai_n526_), .B(mai_mai_n521_), .C(mai_mai_n520_), .Y(mai_mai_n527_));
  NA2        m0499(.A(mai_mai_n265_), .B(mai_mai_n117_), .Y(mai_mai_n528_));
  AOI220     m0500(.A0(mai_mai_n1056_), .A1(mai_mai_n425_), .B0(b), .B1(mai_mai_n91_), .Y(mai_mai_n529_));
  OA210      m0501(.A0(mai_mai_n529_), .A1(mai_mai_n442_), .B0(mai_mai_n289_), .Y(mai_mai_n530_));
  NA2        m0502(.A(mai_mai_n528_), .B(mai_mai_n530_), .Y(mai_mai_n531_));
  NA2        m0503(.A(mai_mai_n215_), .B(j), .Y(mai_mai_n532_));
  NO2        m0504(.A(mai_mai_n143_), .B(i), .Y(mai_mai_n533_));
  NO4        m0505(.A(mai_mai_n423_), .B(n), .C(mai_mai_n107_), .D(mai_mai_n175_), .Y(mai_mai_n534_));
  INV        m0506(.A(mai_mai_n534_), .Y(mai_mai_n535_));
  NA4        m0507(.A(mai_mai_n535_), .B(mai_mai_n532_), .C(mai_mai_n409_), .D(mai_mai_n320_), .Y(mai_mai_n536_));
  NO4        m0508(.A(mai_mai_n536_), .B(mai_mai_n531_), .C(mai_mai_n527_), .D(mai_mai_n517_), .Y(mai_mai_n537_));
  NA4        m0509(.A(mai_mai_n537_), .B(mai_mai_n510_), .C(mai_mai_n481_), .D(mai_mai_n462_), .Y(mai08));
  NO2        m0510(.A(k), .B(h), .Y(mai_mai_n539_));
  AO210      m0511(.A0(mai_mai_n213_), .A1(mai_mai_n356_), .B0(mai_mai_n539_), .Y(mai_mai_n540_));
  NO2        m0512(.A(mai_mai_n540_), .B(mai_mai_n246_), .Y(mai_mai_n541_));
  AOI210     m0513(.A0(c), .A1(mai_mai_n541_), .B0(mai_mai_n386_), .Y(mai_mai_n542_));
  NA2        m0514(.A(b), .B(mai_mai_n282_), .Y(mai_mai_n543_));
  NA4        m0515(.A(mai_mai_n178_), .B(mai_mai_n117_), .C(mai_mai_n43_), .D(h), .Y(mai_mai_n544_));
  NA4        m0516(.A(l), .B(mai_mai_n88_), .C(mai_mai_n61_), .D(mai_mai_n176_), .Y(mai_mai_n545_));
  OAI210     m0517(.A0(mai_mai_n544_), .A1(g), .B0(mai_mai_n545_), .Y(mai_mai_n546_));
  NA2        m0518(.A(mai_mai_n546_), .B(b), .Y(mai_mai_n547_));
  NA4        m0519(.A(mai_mai_n547_), .B(mai_mai_n543_), .C(mai_mai_n542_), .D(mai_mai_n283_), .Y(mai_mai_n548_));
  AN2        m0520(.A(mai_mai_n430_), .B(mai_mai_n78_), .Y(mai_mai_n549_));
  NO4        m0521(.A(mai_mai_n143_), .B(mai_mai_n312_), .C(mai_mai_n90_), .D(g), .Y(mai_mai_n550_));
  AOI210     m0522(.A0(mai_mai_n550_), .A1(b), .B0(mai_mai_n416_), .Y(mai_mai_n551_));
  NO2        m0523(.A(mai_mai_n36_), .B(mai_mai_n175_), .Y(mai_mai_n552_));
  NA2        m0524(.A(e), .B(mai_mai_n281_), .Y(mai_mai_n553_));
  NAi31      m0525(.An(mai_mai_n549_), .B(mai_mai_n553_), .C(mai_mai_n551_), .Y(mai_mai_n554_));
  INV        m0526(.A(mai_mai_n34_), .Y(mai_mai_n555_));
  NA2        m0527(.A(mai_mai_n444_), .B(mai_mai_n111_), .Y(mai_mai_n556_));
  NO2        m0528(.A(mai_mai_n381_), .B(mai_mai_n108_), .Y(mai_mai_n557_));
  AOI210     m0529(.A0(mai_mai_n557_), .A1(mai_mai_n556_), .B0(mai_mai_n555_), .Y(mai_mai_n558_));
  NO3        m0530(.A(mai_mai_n258_), .B(mai_mai_n107_), .C(mai_mai_n39_), .Y(mai_mai_n559_));
  NAi21      m0531(.An(mai_mai_n559_), .B(mai_mai_n545_), .Y(mai_mai_n560_));
  NA2        m0532(.A(mai_mai_n540_), .B(mai_mai_n112_), .Y(mai_mai_n561_));
  AOI220     m0533(.A0(mai_mai_n561_), .A1(mai_mai_n321_), .B0(mai_mai_n560_), .B1(mai_mai_n63_), .Y(mai_mai_n562_));
  OAI210     m0534(.A0(mai_mai_n558_), .A1(mai_mai_n71_), .B0(mai_mai_n562_), .Y(mai_mai_n563_));
  NA2        m0535(.A(b), .B(mai_mai_n41_), .Y(mai_mai_n564_));
  NA2        m0536(.A(mai_mai_n270_), .B(mai_mai_n304_), .Y(mai_mai_n565_));
  NA2        m0537(.A(l), .B(mai_mai_n183_), .Y(mai_mai_n566_));
  NO2        m0538(.A(mai_mai_n566_), .B(mai_mai_n264_), .Y(mai_mai_n567_));
  AOI210     m0539(.A0(mai_mai_n567_), .A1(i), .B0(mai_mai_n385_), .Y(mai_mai_n568_));
  NA3        m0540(.A(m), .B(l), .C(k), .Y(mai_mai_n569_));
  AOI210     m0541(.A0(mai_mai_n514_), .A1(mai_mai_n513_), .B0(mai_mai_n569_), .Y(mai_mai_n570_));
  NOi21      m0542(.An(g), .B(mai_mai_n426_), .Y(mai_mai_n571_));
  NA4        m0543(.A(mai_mai_n91_), .B(l), .C(k), .D(mai_mai_n71_), .Y(mai_mai_n572_));
  NA3        m0544(.A(c), .B(mai_mai_n325_), .C(i), .Y(mai_mai_n573_));
  NO2        m0545(.A(mai_mai_n573_), .B(mai_mai_n572_), .Y(mai_mai_n574_));
  NO3        m0546(.A(mai_mai_n574_), .B(mai_mai_n571_), .C(mai_mai_n570_), .Y(mai_mai_n575_));
  NA4        m0547(.A(mai_mai_n575_), .B(mai_mai_n568_), .C(mai_mai_n565_), .D(mai_mai_n564_), .Y(mai_mai_n576_));
  NO4        m0548(.A(mai_mai_n576_), .B(mai_mai_n563_), .C(mai_mai_n554_), .D(mai_mai_n548_), .Y(mai_mai_n577_));
  NA2        m0549(.A(e), .B(mai_mai_n313_), .Y(mai_mai_n578_));
  NA2        m0550(.A(mai_mai_n494_), .B(g), .Y(mai_mai_n579_));
  AO210      m0551(.A0(mai_mai_n579_), .A1(mai_mai_n466_), .B0(mai_mai_n432_), .Y(mai_mai_n580_));
  AOI210     m0552(.A0(g), .A1(mai_mai_n91_), .B0(mai_mai_n396_), .Y(mai_mai_n581_));
  NA4        m0553(.A(mai_mai_n581_), .B(mai_mai_n580_), .C(mai_mai_n578_), .D(mai_mai_n212_), .Y(mai_mai_n582_));
  NA2        m0554(.A(l), .B(mai_mai_n61_), .Y(mai_mai_n583_));
  NO3        m0555(.A(mai_mai_n143_), .B(n), .C(i), .Y(mai_mai_n584_));
  NOi21      m0556(.An(h), .B(j), .Y(mai_mai_n585_));
  NA2        m0557(.A(mai_mai_n585_), .B(f), .Y(mai_mai_n586_));
  NO2        m0558(.A(mai_mai_n586_), .B(mai_mai_n206_), .Y(mai_mai_n587_));
  NO3        m0559(.A(mai_mai_n587_), .B(mai_mai_n584_), .C(mai_mai_n533_), .Y(mai_mai_n588_));
  OAI210     m0560(.A0(mai_mai_n588_), .A1(mai_mai_n583_), .B0(mai_mai_n468_), .Y(mai_mai_n589_));
  AOI210     m0561(.A0(mai_mai_n582_), .A1(l), .B0(mai_mai_n589_), .Y(mai_mai_n590_));
  NO2        m0562(.A(j), .B(i), .Y(mai_mai_n591_));
  NA2        m0563(.A(mai_mai_n591_), .B(mai_mai_n32_), .Y(mai_mai_n592_));
  NO3        m0564(.A(mai_mai_n127_), .B(mai_mai_n46_), .C(a), .Y(mai_mai_n593_));
  NO2        m0565(.A(mai_mai_n435_), .B(mai_mai_n61_), .Y(mai_mai_n594_));
  OAI210     m0566(.A0(mai_mai_n594_), .A1(mai_mai_n593_), .B0(g), .Y(mai_mai_n595_));
  OAI210     m0567(.A0(mai_mai_n579_), .A1(i), .B0(mai_mai_n595_), .Y(mai_mai_n596_));
  NA2        m0568(.A(k), .B(j), .Y(mai_mai_n597_));
  NO3        m0569(.A(mai_mai_n246_), .B(mai_mai_n597_), .C(mai_mai_n38_), .Y(mai_mai_n598_));
  AN2        m0570(.A(mai_mai_n598_), .B(mai_mai_n79_), .Y(mai_mai_n599_));
  NO3        m0571(.A(mai_mai_n143_), .B(mai_mai_n312_), .C(mai_mai_n90_), .Y(mai_mai_n600_));
  AOI210     m0572(.A0(mai_mai_n600_), .A1(mai_mai_n207_), .B0(mai_mai_n254_), .Y(mai_mai_n601_));
  NA2        m0573(.A(mai_mai_n76_), .B(mai_mai_n70_), .Y(mai_mai_n602_));
  NA2        m0574(.A(mai_mai_n602_), .B(mai_mai_n601_), .Y(mai_mai_n603_));
  NO2        m0575(.A(mai_mai_n246_), .B(mai_mai_n112_), .Y(mai_mai_n604_));
  AOI220     m0576(.A0(mai_mai_n604_), .A1(e), .B0(mai_mai_n559_), .B1(b), .Y(mai_mai_n605_));
  OAI210     m0577(.A0(g), .A1(g), .B0(mai_mai_n525_), .Y(mai_mai_n606_));
  NA2        m0578(.A(mai_mai_n606_), .B(mai_mai_n605_), .Y(mai_mai_n607_));
  OR4        m0579(.A(mai_mai_n607_), .B(mai_mai_n603_), .C(mai_mai_n599_), .D(mai_mai_n596_), .Y(mai_mai_n608_));
  NA3        m0580(.A(mai_mai_n178_), .B(mai_mai_n356_), .C(mai_mai_n33_), .Y(mai_mai_n609_));
  OAI220     m0581(.A0(mai_mai_n544_), .A1(mai_mai_n1063_), .B0(n), .B1(mai_mai_n36_), .Y(mai_mai_n610_));
  AOI210     m0582(.A0(g), .A1(mai_mai_n219_), .B0(mai_mai_n610_), .Y(mai_mai_n611_));
  NO2        m0583(.A(mai_mai_n75_), .B(mai_mai_n1058_), .Y(mai_mai_n612_));
  NA2        m0584(.A(mai_mai_n612_), .B(mai_mai_n498_), .Y(mai_mai_n613_));
  NA3        m0585(.A(mai_mai_n613_), .B(mai_mai_n611_), .C(mai_mai_n609_), .Y(mai_mai_n614_));
  NA2        m0586(.A(g), .B(mai_mai_n493_), .Y(mai_mai_n615_));
  NO2        m0587(.A(n), .B(mai_mai_n61_), .Y(mai_mai_n616_));
  AOI210     m0588(.A0(g), .A1(mai_mai_n616_), .B0(mai_mai_n272_), .Y(mai_mai_n617_));
  OAI210     m0589(.A0(mai_mai_n569_), .A1(mai_mai_n512_), .B0(mai_mai_n415_), .Y(mai_mai_n618_));
  NA2        m0590(.A(mai_mai_n70_), .B(mai_mai_n618_), .Y(mai_mai_n619_));
  NA3        m0591(.A(mai_mai_n619_), .B(mai_mai_n617_), .C(mai_mai_n615_), .Y(mai_mai_n620_));
  NO3        m0592(.A(mai_mai_n620_), .B(mai_mai_n614_), .C(mai_mai_n608_), .Y(mai_mai_n621_));
  NO3        m0593(.A(mai_mai_n277_), .B(mai_mai_n248_), .C(mai_mai_n90_), .Y(mai_mai_n622_));
  INV        m0594(.A(mai_mai_n622_), .Y(mai_mai_n623_));
  NO2        m0595(.A(mai_mai_n592_), .B(mai_mai_n230_), .Y(mai_mai_n624_));
  INV        m0596(.A(mai_mai_n624_), .Y(mai_mai_n625_));
  NA4        m0597(.A(mai_mai_n625_), .B(mai_mai_n623_), .C(mai_mai_n544_), .D(mai_mai_n322_), .Y(mai_mai_n626_));
  OR2        m0598(.A(mai_mai_n512_), .B(mai_mai_n75_), .Y(mai_mai_n627_));
  INV        m0599(.A(n), .Y(mai_mai_n628_));
  NO2        m0600(.A(n), .B(mai_mai_n627_), .Y(mai_mai_n629_));
  NOi21      m0601(.An(l), .B(mai_mai_n134_), .Y(mai_mai_n630_));
  AOI210     m0602(.A0(mai_mai_n622_), .A1(c), .B0(mai_mai_n630_), .Y(mai_mai_n631_));
  OAI210     m0603(.A0(mai_mai_n544_), .A1(mai_mai_n314_), .B0(mai_mai_n631_), .Y(mai_mai_n632_));
  AOI210     m0604(.A0(mai_mai_n604_), .A1(c), .B0(mai_mai_n541_), .Y(mai_mai_n633_));
  AOI210     m0605(.A0(mai_mai_n337_), .A1(mai_mai_n331_), .B0(n), .Y(mai_mai_n634_));
  NA2        m0606(.A(mai_mai_n567_), .B(mai_mai_n33_), .Y(mai_mai_n635_));
  NAi21      m0607(.An(mai_mai_n572_), .B(mai_mai_n345_), .Y(mai_mai_n636_));
  NO2        m0608(.A(mai_mai_n224_), .B(i), .Y(mai_mai_n637_));
  NA2        m0609(.A(mai_mai_n550_), .B(b), .Y(mai_mai_n638_));
  OAI210     m0610(.A0(mai_mai_n470_), .A1(mai_mai_n469_), .B0(mai_mai_n291_), .Y(mai_mai_n639_));
  AN3        m0611(.A(mai_mai_n639_), .B(mai_mai_n638_), .C(mai_mai_n636_), .Y(mai_mai_n640_));
  NAi41      m0612(.An(mai_mai_n634_), .B(mai_mai_n640_), .C(mai_mai_n635_), .D(mai_mai_n633_), .Y(mai_mai_n641_));
  NO4        m0613(.A(mai_mai_n641_), .B(mai_mai_n632_), .C(mai_mai_n629_), .D(mai_mai_n626_), .Y(mai_mai_n642_));
  NA4        m0614(.A(mai_mai_n642_), .B(mai_mai_n621_), .C(mai_mai_n590_), .D(mai_mai_n577_), .Y(mai09));
  INV        m0615(.A(g), .Y(mai_mai_n644_));
  NO2        m0616(.A(g), .B(h), .Y(mai_mai_n645_));
  NA2        m0617(.A(mai_mai_n645_), .B(mai_mai_n644_), .Y(mai_mai_n646_));
  NA2        m0618(.A(mai_mai_n353_), .B(e), .Y(mai_mai_n647_));
  NO2        m0619(.A(mai_mai_n647_), .B(c), .Y(mai_mai_n648_));
  AOI210     m0620(.A0(mai_mai_n646_), .A1(mai_mai_n91_), .B0(mai_mai_n648_), .Y(mai_mai_n649_));
  NA3        m0621(.A(m), .B(l), .C(i), .Y(mai_mai_n650_));
  OAI220     m0622(.A0(mai_mai_n465_), .A1(mai_mai_n650_), .B0(mai_mai_n285_), .B1(mai_mai_n422_), .Y(mai_mai_n651_));
  NA4        m0623(.A(m), .B(mai_mai_n71_), .C(g), .D(f), .Y(mai_mai_n652_));
  NAi31      m0624(.An(mai_mai_n651_), .B(mai_mai_n652_), .C(mai_mai_n348_), .Y(mai_mai_n653_));
  NA3        m0625(.A(mai_mai_n627_), .B(mai_mai_n451_), .C(mai_mai_n415_), .Y(mai_mai_n654_));
  OA210      m0626(.A0(mai_mai_n654_), .A1(n), .B0(mai_mai_n628_), .Y(mai_mai_n655_));
  INV        m0627(.A(mai_mai_n275_), .Y(mai_mai_n656_));
  NO2        m0628(.A(mai_mai_n104_), .B(mai_mai_n102_), .Y(mai_mai_n657_));
  AOI210     m0629(.A0(m), .A1(mai_mai_n657_), .B0(mai_mai_n473_), .Y(mai_mai_n658_));
  NA2        m0630(.A(mai_mai_n278_), .B(m), .Y(mai_mai_n659_));
  OAI210     m0631(.A0(mai_mai_n168_), .A1(mai_mai_n175_), .B0(mai_mai_n659_), .Y(mai_mai_n660_));
  AOI220     m0632(.A0(mai_mai_n660_), .A1(mai_mai_n210_), .B0(mai_mai_n658_), .B1(mai_mai_n656_), .Y(mai_mai_n661_));
  NA3        m0633(.A(mai_mai_n1052_), .B(mai_mai_n157_), .C(mai_mai_n30_), .Y(mai_mai_n662_));
  NA4        m0634(.A(mai_mai_n662_), .B(mai_mai_n661_), .C(mai_mai_n487_), .D(mai_mai_n68_), .Y(mai_mai_n663_));
  INV        m0635(.A(mai_mai_n392_), .Y(mai_mai_n664_));
  NA2        m0636(.A(mai_mai_n664_), .B(mai_mai_n157_), .Y(mai_mai_n665_));
  NA2        m0637(.A(f), .B(m), .Y(mai_mai_n666_));
  NA4        m0638(.A(g), .B(mai_mai_n477_), .C(a), .D(m), .Y(mai_mai_n667_));
  INV        m0639(.A(mai_mai_n667_), .Y(mai_mai_n668_));
  INV        m0640(.A(mai_mai_n668_), .Y(mai_mai_n669_));
  NO3        m0641(.A(n), .B(mai_mai_n61_), .C(mai_mai_n176_), .Y(mai_mai_n670_));
  INV        m0642(.A(mai_mai_n670_), .Y(mai_mai_n671_));
  NAi41      m0643(.An(mai_mai_n384_), .B(mai_mai_n671_), .C(mai_mai_n669_), .D(mai_mai_n665_), .Y(mai_mai_n672_));
  NO3        m0644(.A(mai_mai_n108_), .B(mai_mai_n264_), .C(mai_mai_n128_), .Y(mai_mai_n673_));
  NO2        m0645(.A(mai_mai_n506_), .B(mai_mai_n264_), .Y(mai_mai_n674_));
  AN2        m0646(.A(mai_mai_n674_), .B(i), .Y(mai_mai_n675_));
  NO3        m0647(.A(mai_mai_n675_), .B(mai_mai_n673_), .C(mai_mai_n194_), .Y(mai_mai_n676_));
  OAI220     m0648(.A0(mai_mai_n659_), .A1(n), .B0(n), .B1(mai_mai_n348_), .Y(mai_mai_n677_));
  NA3        m0649(.A(mai_mai_n133_), .B(mai_mai_n88_), .C(g), .Y(mai_mai_n678_));
  OAI220     m0650(.A0(n), .A1(mai_mai_n340_), .B0(mai_mai_n275_), .B1(mai_mai_n678_), .Y(mai_mai_n679_));
  NOi41      m0651(.An(mai_mai_n186_), .B(mai_mai_n679_), .C(mai_mai_n677_), .D(mai_mai_n252_), .Y(mai_mai_n680_));
  NA2        m0652(.A(c), .B(mai_mai_n94_), .Y(mai_mai_n681_));
  NA3        m0653(.A(e), .B(mai_mai_n405_), .C(f), .Y(mai_mai_n682_));
  OR2        m0654(.A(mai_mai_n512_), .B(mai_mai_n433_), .Y(mai_mai_n683_));
  NA4        m0655(.A(mai_mai_n683_), .B(mai_mai_n682_), .C(mai_mai_n680_), .D(mai_mai_n676_), .Y(mai_mai_n684_));
  NO4        m0656(.A(mai_mai_n684_), .B(mai_mai_n672_), .C(mai_mai_n663_), .D(mai_mai_n655_), .Y(mai_mai_n685_));
  OR2        m0657(.A(n), .B(mai_mai_n61_), .Y(mai_mai_n686_));
  INV        m0658(.A(g), .Y(mai_mai_n687_));
  AOI210     m0659(.A0(mai_mai_n687_), .A1(mai_mai_n242_), .B0(mai_mai_n686_), .Y(mai_mai_n688_));
  AOI210     m0660(.A0(n), .A1(n), .B0(mai_mai_n652_), .Y(mai_mai_n689_));
  NO2        m0661(.A(mai_mai_n112_), .B(mai_mai_n108_), .Y(mai_mai_n690_));
  NO2        m0662(.A(mai_mai_n191_), .B(mai_mai_n187_), .Y(mai_mai_n691_));
  AOI220     m0663(.A0(mai_mai_n691_), .A1(mai_mai_n188_), .B0(mai_mai_n251_), .B1(mai_mai_n690_), .Y(mai_mai_n692_));
  INV        m0664(.A(mai_mai_n340_), .Y(mai_mai_n693_));
  NA2        m0665(.A(mai_mai_n693_), .B(mai_mai_n446_), .Y(mai_mai_n694_));
  NA2        m0666(.A(mai_mai_n694_), .B(mai_mai_n692_), .Y(mai_mai_n695_));
  NA2        m0667(.A(e), .B(d), .Y(mai_mai_n696_));
  NA3        m0668(.A(e), .B(mai_mai_n360_), .C(mai_mai_n403_), .Y(mai_mai_n697_));
  AOI210     m0669(.A0(mai_mai_n410_), .A1(mai_mai_n150_), .B0(mai_mai_n191_), .Y(mai_mai_n698_));
  AOI210     m0670(.A0(e), .A1(mai_mai_n281_), .B0(mai_mai_n698_), .Y(mai_mai_n699_));
  NA3        m0671(.A(mai_mai_n670_), .B(j), .C(mai_mai_n50_), .Y(mai_mai_n700_));
  NA3        m0672(.A(mai_mai_n139_), .B(b), .C(mai_mai_n33_), .Y(mai_mai_n701_));
  NA4        m0673(.A(mai_mai_n701_), .B(mai_mai_n700_), .C(mai_mai_n699_), .D(mai_mai_n697_), .Y(mai_mai_n702_));
  NO4        m0674(.A(mai_mai_n702_), .B(mai_mai_n695_), .C(mai_mai_n689_), .D(mai_mai_n688_), .Y(mai_mai_n703_));
  AO210      m0675(.A0(mai_mai_n275_), .A1(mai_mai_n1063_), .B0(mai_mai_n179_), .Y(mai_mai_n704_));
  AOI220     m0676(.A0(h), .A1(mai_mai_n674_), .B0(mai_mai_n482_), .B1(e), .Y(mai_mai_n705_));
  OAI210     m0677(.A0(mai_mai_n647_), .A1(d), .B0(mai_mai_n705_), .Y(mai_mai_n706_));
  OAI210     m0678(.A0(l), .A1(j), .B0(g), .Y(mai_mai_n707_));
  NO2        m0679(.A(mai_mai_n707_), .B(mai_mai_n478_), .Y(mai_mai_n708_));
  INV        m0680(.A(mai_mai_n667_), .Y(mai_mai_n709_));
  AO210      m0681(.A0(mai_mai_n210_), .A1(mai_mai_n651_), .B0(mai_mai_n709_), .Y(mai_mai_n710_));
  NOi31      m0682(.An(mai_mai_n436_), .B(mai_mai_n666_), .C(mai_mai_n242_), .Y(mai_mai_n711_));
  NO4        m0683(.A(mai_mai_n711_), .B(mai_mai_n710_), .C(mai_mai_n708_), .D(mai_mai_n706_), .Y(mai_mai_n712_));
  AO220      m0684(.A0(mai_mai_n360_), .A1(mai_mai_n585_), .B0(mai_mai_n145_), .B1(f), .Y(mai_mai_n713_));
  OAI210     m0685(.A0(mai_mai_n713_), .A1(mai_mai_n363_), .B0(e), .Y(mai_mai_n714_));
  NO2        m0686(.A(mai_mai_n347_), .B(mai_mai_n57_), .Y(mai_mai_n715_));
  OAI210     m0687(.A0(mai_mai_n654_), .A1(mai_mai_n715_), .B0(mai_mai_n1059_), .Y(mai_mai_n716_));
  AN4        m0688(.A(mai_mai_n716_), .B(mai_mai_n714_), .C(mai_mai_n712_), .D(mai_mai_n704_), .Y(mai_mai_n717_));
  NA4        m0689(.A(mai_mai_n717_), .B(mai_mai_n703_), .C(mai_mai_n685_), .D(mai_mai_n649_), .Y(mai12));
  NO4        m0690(.A(mai_mai_n352_), .B(mai_mai_n213_), .C(mai_mai_n463_), .D(mai_mai_n176_), .Y(mai_mai_n719_));
  NA2        m0691(.A(mai_mai_n719_), .B(d), .Y(mai_mai_n720_));
  NA2        m0692(.A(mai_mai_n436_), .B(mai_mai_n715_), .Y(mai_mai_n721_));
  NO2        m0693(.A(mai_mai_n657_), .B(mai_mai_n285_), .Y(mai_mai_n722_));
  NO2        m0694(.A(mai_mai_n512_), .B(mai_mai_n303_), .Y(mai_mai_n723_));
  AOI220     m0695(.A0(mai_mai_n723_), .A1(mai_mai_n1060_), .B0(mai_mai_n722_), .B1(d), .Y(mai_mai_n724_));
  NA4        m0696(.A(mai_mai_n724_), .B(mai_mai_n721_), .C(mai_mai_n720_), .D(mai_mai_n351_), .Y(mai_mai_n725_));
  AOI210     m0697(.A0(mai_mai_n193_), .A1(mai_mai_n274_), .B0(mai_mai_n166_), .Y(mai_mai_n726_));
  OR2        m0698(.A(mai_mai_n726_), .B(mai_mai_n719_), .Y(mai_mai_n727_));
  AOI210     m0699(.A0(mai_mai_n271_), .A1(mai_mai_n310_), .B0(mai_mai_n176_), .Y(mai_mai_n728_));
  OAI210     m0700(.A0(mai_mai_n728_), .A1(mai_mai_n727_), .B0(d), .Y(mai_mai_n729_));
  NO2        m0701(.A(mai_mai_n465_), .B(mai_mai_n650_), .Y(mai_mai_n730_));
  NA3        m0702(.A(mai_mai_n1062_), .B(mai_mai_n200_), .C(i), .Y(mai_mai_n731_));
  NA2        m0703(.A(mai_mai_n731_), .B(mai_mai_n729_), .Y(mai_mai_n732_));
  INV        m0704(.A(mai_mai_n286_), .Y(mai_mai_n733_));
  NO3        m0705(.A(mai_mai_n108_), .B(mai_mai_n128_), .C(mai_mai_n176_), .Y(mai_mai_n734_));
  NA2        m0706(.A(mai_mai_n734_), .B(mai_mai_n425_), .Y(mai_mai_n735_));
  NA4        m0707(.A(mai_mai_n353_), .B(d), .C(mai_mai_n151_), .D(g), .Y(mai_mai_n736_));
  NA3        m0708(.A(mai_mai_n736_), .B(mai_mai_n735_), .C(mai_mai_n733_), .Y(mai_mai_n737_));
  NO3        m0709(.A(mai_mai_n516_), .B(mai_mai_n75_), .C(mai_mai_n43_), .Y(mai_mai_n738_));
  NO4        m0710(.A(mai_mai_n738_), .B(mai_mai_n737_), .C(mai_mai_n732_), .D(mai_mai_n725_), .Y(mai_mai_n739_));
  NOi21      m0711(.An(mai_mai_n33_), .B(mai_mai_n506_), .Y(mai_mai_n740_));
  NA2        m0712(.A(mai_mai_n740_), .B(c), .Y(mai_mai_n741_));
  OAI210     m0713(.A0(mai_mai_n211_), .A1(mai_mai_n43_), .B0(mai_mai_n741_), .Y(mai_mai_n742_));
  NA2        m0714(.A(mai_mai_n345_), .B(mai_mai_n220_), .Y(mai_mai_n743_));
  NO2        m0715(.A(n), .B(mai_mai_n72_), .Y(mai_mai_n744_));
  NAi31      m0716(.An(mai_mai_n744_), .B(mai_mai_n743_), .C(mai_mai_n262_), .Y(mai_mai_n745_));
  NO2        m0717(.A(mai_mai_n399_), .B(mai_mai_n248_), .Y(mai_mai_n746_));
  NO2        m0718(.A(mai_mai_n173_), .B(f), .Y(mai_mai_n747_));
  OAI210     m0719(.A0(mai_mai_n573_), .A1(n), .B0(mai_mai_n295_), .Y(mai_mai_n748_));
  NO4        m0720(.A(mai_mai_n748_), .B(mai_mai_n747_), .C(mai_mai_n745_), .D(mai_mai_n742_), .Y(mai_mai_n749_));
  NA2        m0721(.A(mai_mai_n281_), .B(g), .Y(mai_mai_n750_));
  NA2        m0722(.A(h), .B(i), .Y(mai_mai_n751_));
  NA2        m0723(.A(mai_mai_n44_), .B(i), .Y(mai_mai_n752_));
  OAI220     m0724(.A0(mai_mai_n752_), .A1(mai_mai_n1051_), .B0(mai_mai_n751_), .B1(mai_mai_n75_), .Y(mai_mai_n753_));
  AOI210     m0725(.A0(m), .A1(mai_mai_n35_), .B0(mai_mai_n753_), .Y(mai_mai_n754_));
  OAI210     m0726(.A0(mai_mai_n754_), .A1(n), .B0(mai_mai_n750_), .Y(mai_mai_n755_));
  OAI220     m0727(.A0(g), .A1(h), .B0(mai_mai_n525_), .B1(mai_mai_n594_), .Y(mai_mai_n756_));
  NA2        m0728(.A(a), .B(mai_mai_n91_), .Y(mai_mai_n757_));
  NA3        m0729(.A(f), .B(mai_mai_n96_), .C(g), .Y(mai_mai_n758_));
  AOI210     m0730(.A0(mai_mai_n522_), .A1(mai_mai_n758_), .B0(m), .Y(mai_mai_n759_));
  OAI210     m0731(.A0(mai_mai_n759_), .A1(mai_mai_n722_), .B0(c), .Y(mai_mai_n760_));
  NA2        m0732(.A(mai_mai_n652_), .B(mai_mai_n348_), .Y(mai_mai_n761_));
  AOI220     m0733(.A0(h), .A1(mai_mai_n219_), .B0(mai_mai_n761_), .B1(mai_mai_n70_), .Y(mai_mai_n762_));
  NA3        m0734(.A(mai_mai_n762_), .B(mai_mai_n760_), .C(mai_mai_n756_), .Y(mai_mai_n763_));
  OAI210     m0735(.A0(m), .A1(m), .B0(mai_mai_n198_), .Y(mai_mai_n764_));
  NA2        m0736(.A(mai_mai_n515_), .B(m), .Y(mai_mai_n765_));
  NO2        m0737(.A(mai_mai_n366_), .B(mai_mai_n176_), .Y(mai_mai_n766_));
  AOI210     m0738(.A0(mai_mai_n766_), .A1(c), .B0(mai_mai_n180_), .Y(mai_mai_n767_));
  NA2        m0739(.A(mai_mai_n723_), .B(mai_mai_n1062_), .Y(mai_mai_n768_));
  NA4        m0740(.A(mai_mai_n768_), .B(mai_mai_n767_), .C(mai_mai_n765_), .D(mai_mai_n764_), .Y(mai_mai_n769_));
  OAI210     m0741(.A0(mai_mai_n761_), .A1(mai_mai_n730_), .B0(mai_mai_n1060_), .Y(mai_mai_n770_));
  AOI210     m0742(.A0(mai_mai_n332_), .A1(mai_mai_n326_), .B0(n), .Y(mai_mai_n771_));
  AOI210     m0743(.A0(mai_mai_n172_), .A1(mai_mai_n430_), .B0(mai_mai_n771_), .Y(mai_mai_n772_));
  NA2        m0744(.A(mai_mai_n759_), .B(d), .Y(mai_mai_n773_));
  NO2        m0745(.A(mai_mai_n46_), .B(mai_mai_n43_), .Y(mai_mai_n774_));
  AOI220     m0746(.A0(mai_mai_n774_), .A1(g), .B0(mai_mai_n500_), .B1(mai_mai_n425_), .Y(mai_mai_n775_));
  NA4        m0747(.A(mai_mai_n775_), .B(mai_mai_n773_), .C(mai_mai_n772_), .D(mai_mai_n770_), .Y(mai_mai_n776_));
  NO4        m0748(.A(mai_mai_n776_), .B(mai_mai_n769_), .C(mai_mai_n763_), .D(mai_mai_n755_), .Y(mai_mai_n777_));
  NAi31      m0749(.An(mai_mai_n118_), .B(mai_mai_n333_), .C(n), .Y(mai_mai_n778_));
  NO2        m0750(.A(m), .B(mai_mai_n778_), .Y(mai_mai_n779_));
  INV        m0751(.A(mai_mai_n224_), .Y(mai_mai_n780_));
  AOI210     m0752(.A0(mai_mai_n780_), .A1(mai_mai_n393_), .B0(mai_mai_n779_), .Y(mai_mai_n781_));
  NA2        m0753(.A(mai_mai_n386_), .B(i), .Y(mai_mai_n782_));
  NA2        m0754(.A(mai_mai_n782_), .B(mai_mai_n781_), .Y(mai_mai_n783_));
  NO3        m0755(.A(mai_mai_n254_), .B(mai_mai_n353_), .C(mai_mai_n145_), .Y(mai_mai_n784_));
  NOi31      m0756(.An(c), .B(mai_mai_n784_), .C(mai_mai_n176_), .Y(mai_mai_n785_));
  NAi21      m0757(.An(mai_mai_n444_), .B(mai_mai_n766_), .Y(mai_mai_n786_));
  NO3        m0758(.A(mai_mai_n347_), .B(k), .C(mai_mai_n61_), .Y(mai_mai_n787_));
  AOI220     m0759(.A0(mai_mai_n787_), .A1(mai_mai_n346_), .B0(mai_mai_n379_), .B1(g), .Y(mai_mai_n788_));
  NA2        m0760(.A(mai_mai_n788_), .B(mai_mai_n786_), .Y(mai_mai_n789_));
  NO2        m0761(.A(mai_mai_n778_), .B(mai_mai_n193_), .Y(mai_mai_n790_));
  NO2        m0762(.A(mai_mai_n513_), .B(mai_mai_n303_), .Y(mai_mai_n791_));
  NA2        m0763(.A(mai_mai_n726_), .B(d), .Y(mai_mai_n792_));
  OAI220     m0764(.A0(mai_mai_n723_), .A1(mai_mai_n730_), .B0(mai_mai_n436_), .B1(mai_mai_n339_), .Y(mai_mai_n793_));
  NA3        m0765(.A(mai_mai_n793_), .B(mai_mai_n792_), .C(mai_mai_n486_), .Y(mai_mai_n794_));
  OAI210     m0766(.A0(mai_mai_n726_), .A1(mai_mai_n719_), .B0(c), .Y(mai_mai_n795_));
  NA3        m0767(.A(c), .B(mai_mai_n382_), .C(mai_mai_n44_), .Y(mai_mai_n796_));
  INV        m0768(.A(mai_mai_n268_), .Y(mai_mai_n797_));
  NA4        m0769(.A(mai_mai_n797_), .B(mai_mai_n796_), .C(mai_mai_n795_), .D(mai_mai_n225_), .Y(mai_mai_n798_));
  OR4        m0770(.A(mai_mai_n798_), .B(mai_mai_n794_), .C(mai_mai_n791_), .D(mai_mai_n790_), .Y(mai_mai_n799_));
  NO4        m0771(.A(mai_mai_n799_), .B(mai_mai_n789_), .C(mai_mai_n785_), .D(mai_mai_n783_), .Y(mai_mai_n800_));
  NA4        m0772(.A(mai_mai_n800_), .B(mai_mai_n777_), .C(mai_mai_n749_), .D(mai_mai_n739_), .Y(mai13));
  NA3        m0773(.A(mai_mai_n210_), .B(b), .C(m), .Y(mai_mai_n802_));
  NA2        m0774(.A(d), .B(f), .Y(mai_mai_n803_));
  NO4        m0775(.A(mai_mai_n803_), .B(mai_mai_n802_), .C(j), .D(k), .Y(mai_mai_n804_));
  NO4        m0776(.A(mai_mai_n55_), .B(mai_mai_n803_), .C(mai_mai_n751_), .D(a), .Y(mai_mai_n805_));
  NAi32      m0777(.An(d), .Bn(c), .C(e), .Y(mai_mai_n806_));
  NA2        m0778(.A(mai_mai_n117_), .B(mai_mai_n43_), .Y(mai_mai_n807_));
  NO4        m0779(.A(mai_mai_n807_), .B(mai_mai_n806_), .C(mai_mai_n465_), .D(mai_mai_n253_), .Y(mai_mai_n808_));
  NA2        m0780(.A(mai_mai_n325_), .B(mai_mai_n175_), .Y(mai_mai_n809_));
  AN2        m0781(.A(d), .B(c), .Y(mai_mai_n810_));
  NA2        m0782(.A(mai_mai_n810_), .B(mai_mai_n94_), .Y(mai_mai_n811_));
  NO3        m0783(.A(mai_mai_n811_), .B(mai_mai_n809_), .C(mai_mai_n146_), .Y(mai_mai_n812_));
  NO3        m0784(.A(mai_mai_n807_), .B(h), .C(mai_mai_n253_), .Y(mai_mai_n813_));
  OR2        m0785(.A(mai_mai_n812_), .B(mai_mai_n813_), .Y(mai_mai_n814_));
  OR4        m0786(.A(mai_mai_n814_), .B(mai_mai_n808_), .C(mai_mai_n805_), .D(mai_mai_n804_), .Y(mai_mai_n815_));
  NAi32      m0787(.An(f), .Bn(e), .C(c), .Y(mai_mai_n816_));
  NO2        m0788(.A(mai_mai_n816_), .B(mai_mai_n123_), .Y(mai_mai_n817_));
  NA2        m0789(.A(mai_mai_n817_), .B(g), .Y(mai_mai_n818_));
  NO2        m0790(.A(mai_mai_n146_), .B(mai_mai_n818_), .Y(mai_mai_n819_));
  NO2        m0791(.A(e), .B(mai_mai_n253_), .Y(mai_mai_n820_));
  NOi21      m0792(.An(mai_mai_n820_), .B(f), .Y(mai_mai_n821_));
  NOi41      m0793(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n822_));
  NO2        m0794(.A(mai_mai_n1054_), .B(mai_mai_n818_), .Y(mai_mai_n823_));
  NA3        m0795(.A(k), .B(j), .C(i), .Y(mai_mai_n824_));
  NO2        m0796(.A(mai_mai_n824_), .B(mai_mai_n253_), .Y(mai_mai_n825_));
  OR4        m0797(.A(mai_mai_n825_), .B(mai_mai_n823_), .C(mai_mai_n821_), .D(mai_mai_n819_), .Y(mai_mai_n826_));
  NA3        m0798(.A(mai_mai_n372_), .B(mai_mai_n270_), .C(mai_mai_n50_), .Y(mai_mai_n827_));
  NO2        m0799(.A(mai_mai_n827_), .B(f), .Y(mai_mai_n828_));
  NO3        m0800(.A(mai_mai_n827_), .B(mai_mai_n356_), .C(mai_mai_n43_), .Y(mai_mai_n829_));
  NO2        m0801(.A(f), .B(c), .Y(mai_mai_n830_));
  NOi21      m0802(.An(mai_mai_n830_), .B(mai_mai_n352_), .Y(mai_mai_n831_));
  NA2        m0803(.A(mai_mai_n831_), .B(mai_mai_n51_), .Y(mai_mai_n832_));
  OR3        m0804(.A(mai_mai_n831_), .B(mai_mai_n826_), .C(mai_mai_n815_), .Y(mai02));
  OR2        m0805(.A(l), .B(k), .Y(mai_mai_n834_));
  OR3        m0806(.A(n), .B(m), .C(i), .Y(mai_mai_n835_));
  NO4        m0807(.A(mai_mai_n835_), .B(h), .C(mai_mai_n834_), .D(c), .Y(mai_mai_n836_));
  NO2        m0808(.A(mai_mai_n825_), .B(mai_mai_n808_), .Y(mai_mai_n837_));
  OR2        m0809(.A(mai_mai_n824_), .B(mai_mai_n253_), .Y(mai_mai_n838_));
  NO3        m0810(.A(mai_mai_n827_), .B(mai_mai_n807_), .C(h), .Y(mai_mai_n839_));
  NO2        m0811(.A(mai_mai_n839_), .B(mai_mai_n819_), .Y(mai_mai_n840_));
  NA3        m0812(.A(l), .B(k), .C(j), .Y(mai_mai_n841_));
  NA2        m0813(.A(i), .B(h), .Y(mai_mai_n842_));
  NO3        m0814(.A(mai_mai_n842_), .B(mai_mai_n841_), .C(mai_mai_n108_), .Y(mai_mai_n843_));
  NO3        m0815(.A(mai_mai_n119_), .B(mai_mai_n237_), .C(mai_mai_n176_), .Y(mai_mai_n844_));
  AOI210     m0816(.A0(mai_mai_n844_), .A1(mai_mai_n843_), .B0(mai_mai_n821_), .Y(mai_mai_n845_));
  NA3        m0817(.A(c), .B(b), .C(a), .Y(mai_mai_n846_));
  NO3        m0818(.A(mai_mai_n846_), .B(mai_mai_n696_), .C(mai_mai_n175_), .Y(mai_mai_n847_));
  AOI210     m0819(.A0(g), .A1(mai_mai_n847_), .B0(mai_mai_n828_), .Y(mai_mai_n848_));
  AN4        m0820(.A(mai_mai_n848_), .B(mai_mai_n845_), .C(mai_mai_n840_), .D(mai_mai_n838_), .Y(mai_mai_n849_));
  NO2        m0821(.A(mai_mai_n811_), .B(mai_mai_n809_), .Y(mai_mai_n850_));
  NA2        m0822(.A(mai_mai_n1054_), .B(mai_mai_n146_), .Y(mai_mai_n851_));
  AOI210     m0823(.A0(mai_mai_n851_), .A1(mai_mai_n850_), .B0(mai_mai_n804_), .Y(mai_mai_n852_));
  NAi41      m0824(.An(mai_mai_n836_), .B(mai_mai_n852_), .C(mai_mai_n849_), .D(mai_mai_n837_), .Y(mai03));
  NOi41      m0825(.An(mai_mai_n627_), .B(mai_mai_n660_), .C(mai_mai_n653_), .D(mai_mai_n552_), .Y(mai_mai_n854_));
  NO2        m0826(.A(mai_mai_n854_), .B(n), .Y(mai_mai_n855_));
  NA4        m0827(.A(i), .B(e), .C(mai_mai_n278_), .D(mai_mai_n270_), .Y(mai_mai_n856_));
  OAI210     m0828(.A0(n), .A1(mai_mai_n334_), .B0(mai_mai_n856_), .Y(mai_mai_n857_));
  NOi31      m0829(.An(m), .B(n), .C(f), .Y(mai_mai_n858_));
  NA2        m0830(.A(mai_mai_n858_), .B(mai_mai_n48_), .Y(mai_mai_n859_));
  OAI210     m0831(.A0(mai_mai_n683_), .A1(b), .B0(mai_mai_n859_), .Y(mai_mai_n860_));
  NOi21      m0832(.An(g), .B(mai_mai_n802_), .Y(mai_mai_n861_));
  NO4        m0833(.A(mai_mai_n861_), .B(mai_mai_n860_), .C(mai_mai_n857_), .D(mai_mai_n771_), .Y(mai_mai_n862_));
  INV        m0834(.A(mai_mai_n808_), .Y(mai_mai_n863_));
  NA3        m0835(.A(mai_mai_n832_), .B(mai_mai_n863_), .C(mai_mai_n862_), .Y(mai_mai_n864_));
  NO4        m0836(.A(mai_mai_n864_), .B(mai_mai_n855_), .C(mai_mai_n634_), .D(mai_mai_n450_), .Y(mai_mai_n865_));
  NA2        m0837(.A(c), .B(b), .Y(mai_mai_n866_));
  NA3        m0838(.A(mai_mai_n339_), .B(mai_mai_n445_), .C(f), .Y(mai_mai_n867_));
  OAI210     m0839(.A0(mai_mai_n439_), .A1(mai_mai_n37_), .B0(c), .Y(mai_mai_n868_));
  NA2        m0840(.A(mai_mai_n868_), .B(mai_mai_n867_), .Y(mai_mai_n869_));
  NAi21      m0841(.An(f), .B(d), .Y(mai_mai_n870_));
  NO2        m0842(.A(mai_mai_n870_), .B(mai_mai_n846_), .Y(mai_mai_n871_));
  AOI210     m0843(.A0(mai_mai_n871_), .A1(mai_mai_n91_), .B0(mai_mai_n869_), .Y(mai_mai_n872_));
  NO2        m0844(.A(mai_mai_n152_), .B(mai_mai_n197_), .Y(mai_mai_n873_));
  NA2        m0845(.A(mai_mai_n873_), .B(m), .Y(mai_mai_n874_));
  AOI210     m0846(.A0(mai_mai_n53_), .A1(mai_mai_n107_), .B0(mai_mai_n874_), .Y(mai_mai_n875_));
  NA2        m0847(.A(mai_mai_n446_), .B(mai_mai_n324_), .Y(mai_mai_n876_));
  NA2        m0848(.A(mai_mai_n91_), .B(mai_mai_n871_), .Y(mai_mai_n877_));
  NO2        m0849(.A(mai_mai_n297_), .B(d), .Y(mai_mai_n878_));
  AOI210     m0850(.A0(mai_mai_n873_), .A1(mai_mai_n341_), .B0(mai_mai_n744_), .Y(mai_mai_n879_));
  NAi41      m0851(.An(mai_mai_n878_), .B(mai_mai_n879_), .C(mai_mai_n877_), .D(mai_mai_n876_), .Y(mai_mai_n880_));
  NO2        m0852(.A(mai_mai_n880_), .B(mai_mai_n875_), .Y(mai_mai_n881_));
  NA3        m0853(.A(mai_mai_n881_), .B(mai_mai_n872_), .C(mai_mai_n865_), .Y(mai00));
  AOI210     m0854(.A0(mai_mai_n247_), .A1(mai_mai_n176_), .B0(mai_mai_n229_), .Y(mai_mai_n883_));
  NO2        m0855(.A(mai_mai_n883_), .B(mai_mai_n458_), .Y(mai_mai_n884_));
  INV        m0856(.A(mai_mai_n857_), .Y(mai_mai_n885_));
  NO3        m0857(.A(mai_mai_n839_), .B(mai_mai_n744_), .C(mai_mai_n549_), .Y(mai_mai_n886_));
  NA3        m0858(.A(mai_mai_n886_), .B(mai_mai_n885_), .C(mai_mai_n772_), .Y(mai_mai_n887_));
  NA2        m0859(.A(mai_mai_n405_), .B(f), .Y(mai_mai_n888_));
  OAI210     m0860(.A0(m), .A1(mai_mai_n38_), .B0(mai_mai_n501_), .Y(mai_mai_n889_));
  NA3        m0861(.A(mai_mai_n889_), .B(mai_mai_n218_), .C(n), .Y(mai_mai_n890_));
  AOI210     m0862(.A0(mai_mai_n890_), .A1(mai_mai_n888_), .B0(mai_mai_n811_), .Y(mai_mai_n891_));
  NO4        m0863(.A(mai_mai_n891_), .B(mai_mai_n887_), .C(mai_mai_n884_), .D(mai_mai_n826_), .Y(mai_mai_n892_));
  NA3        m0864(.A(mai_mai_n139_), .B(mai_mai_n44_), .C(mai_mai_n43_), .Y(mai_mai_n893_));
  NOi31      m0865(.An(n), .B(m), .C(i), .Y(mai_mai_n894_));
  NA3        m0866(.A(mai_mai_n894_), .B(d), .C(mai_mai_n48_), .Y(mai_mai_n895_));
  NA2        m0867(.A(mai_mai_n893_), .B(mai_mai_n895_), .Y(mai_mai_n896_));
  INV        m0868(.A(mai_mai_n457_), .Y(mai_mai_n897_));
  NO4        m0869(.A(mai_mai_n897_), .B(mai_mai_n896_), .C(mai_mai_n878_), .D(mai_mai_n711_), .Y(mai_mai_n898_));
  NO4        m0870(.A(mai_mai_n1055_), .B(mai_mai_n287_), .C(mai_mai_n866_), .D(mai_mai_n51_), .Y(mai_mai_n899_));
  NA3        m0871(.A(mai_mai_n304_), .B(mai_mai_n183_), .C(g), .Y(mai_mai_n900_));
  NO2        m0872(.A(h), .B(g), .Y(mai_mai_n901_));
  NA4        m0873(.A(mai_mai_n393_), .B(mai_mai_n372_), .C(mai_mai_n901_), .D(b), .Y(mai_mai_n902_));
  OAI210     m0874(.A0(mai_mai_n422_), .A1(mai_mai_n473_), .B0(mai_mai_n74_), .Y(mai_mai_n903_));
  AOI220     m0875(.A0(mai_mai_n903_), .A1(mai_mai_n430_), .B0(mai_mai_n734_), .B1(mai_mai_n456_), .Y(mai_mai_n904_));
  AOI220     m0876(.A0(mai_mai_n259_), .A1(mai_mai_n207_), .B0(mai_mai_n147_), .B1(mai_mai_n125_), .Y(mai_mai_n905_));
  NA4        m0877(.A(mai_mai_n905_), .B(mai_mai_n904_), .C(mai_mai_n902_), .D(mai_mai_n900_), .Y(mai_mai_n906_));
  NO3        m0878(.A(mai_mai_n906_), .B(mai_mai_n899_), .C(mai_mai_n219_), .Y(mai_mai_n907_));
  INV        m0879(.A(mai_mai_n263_), .Y(mai_mai_n908_));
  AOI210     m0880(.A0(mai_mai_n207_), .A1(mai_mai_n281_), .B0(mai_mai_n459_), .Y(mai_mai_n909_));
  NA3        m0881(.A(mai_mai_n909_), .B(mai_mai_n908_), .C(mai_mai_n130_), .Y(mai_mai_n910_));
  NO2        m0882(.A(mai_mai_n199_), .B(mai_mai_n151_), .Y(mai_mai_n911_));
  NA2        m0883(.A(mai_mai_n911_), .B(mai_mai_n339_), .Y(mai_mai_n912_));
  NA3        m0884(.A(mai_mai_n149_), .B(mai_mai_n90_), .C(g), .Y(mai_mai_n913_));
  NOi31      m0885(.An(j), .B(h), .C(mai_mai_n913_), .Y(mai_mai_n914_));
  NAi31      m0886(.An(mai_mai_n153_), .B(mai_mai_n664_), .C(mai_mai_n372_), .Y(mai_mai_n915_));
  NAi31      m0887(.An(mai_mai_n914_), .B(mai_mai_n915_), .C(mai_mai_n912_), .Y(mai_mai_n916_));
  NO2        m0888(.A(mai_mai_n228_), .B(mai_mai_n61_), .Y(mai_mai_n917_));
  NO2        m0889(.A(b), .B(n), .Y(mai_mai_n918_));
  AOI210     m0890(.A0(mai_mai_n918_), .A1(mai_mai_n917_), .B0(mai_mai_n836_), .Y(mai_mai_n919_));
  NAi31      m0891(.An(mai_mai_n813_), .B(mai_mai_n919_), .C(mai_mai_n60_), .Y(mai_mai_n920_));
  NO4        m0892(.A(mai_mai_n920_), .B(mai_mai_n916_), .C(mai_mai_n910_), .D(mai_mai_n414_), .Y(mai_mai_n921_));
  AN3        m0893(.A(mai_mai_n921_), .B(mai_mai_n907_), .C(mai_mai_n898_), .Y(mai_mai_n922_));
  NA2        m0894(.A(mai_mai_n430_), .B(mai_mai_n81_), .Y(mai_mai_n923_));
  NA3        m0895(.A(mai_mai_n858_), .B(a), .C(h), .Y(mai_mai_n924_));
  NA4        m0896(.A(mai_mai_n924_), .B(mai_mai_n447_), .C(mai_mai_n923_), .D(mai_mai_n201_), .Y(mai_mai_n925_));
  NA2        m0897(.A(g), .B(mai_mai_n430_), .Y(mai_mai_n926_));
  NA4        m0898(.A(d), .B(mai_mai_n170_), .C(mai_mai_n183_), .D(h), .Y(mai_mai_n927_));
  NA3        m0899(.A(mai_mai_n927_), .B(mai_mai_n926_), .C(mai_mai_n244_), .Y(mai_mai_n928_));
  OAI210     m0900(.A0(mai_mai_n371_), .A1(mai_mai_n97_), .B0(mai_mai_n667_), .Y(mai_mai_n929_));
  AOI210     m0901(.A0(mai_mai_n446_), .A1(mai_mai_n324_), .B0(mai_mai_n929_), .Y(mai_mai_n930_));
  OR3        m0902(.A(mai_mai_n224_), .B(mai_mai_n185_), .C(e), .Y(mai_mai_n931_));
  NO2        m0903(.A(mai_mai_n179_), .B(mai_mai_n176_), .Y(mai_mai_n932_));
  NA2        m0904(.A(n), .B(e), .Y(mai_mai_n933_));
  NO2        m0905(.A(mai_mai_n933_), .B(mai_mai_n123_), .Y(mai_mai_n934_));
  AOI220     m0906(.A0(mai_mai_n934_), .A1(mai_mai_n226_), .B0(mai_mai_n656_), .B1(mai_mai_n932_), .Y(mai_mai_n935_));
  OAI210     m0907(.A0(h), .A1(g), .B0(mai_mai_n355_), .Y(mai_mai_n936_));
  NA4        m0908(.A(mai_mai_n936_), .B(mai_mai_n935_), .C(mai_mai_n931_), .D(mai_mai_n930_), .Y(mai_mai_n937_));
  AOI210     m0909(.A0(mai_mai_n934_), .A1(mai_mai_n658_), .B0(mai_mai_n634_), .Y(mai_mai_n938_));
  AOI220     m0910(.A0(mai_mai_n740_), .A1(mai_mai_n456_), .B0(d), .B1(mai_mai_n204_), .Y(mai_mai_n939_));
  NO2        m0911(.A(mai_mai_n54_), .B(h), .Y(mai_mai_n940_));
  NO2        m0912(.A(mai_mai_n809_), .B(mai_mai_n566_), .Y(mai_mai_n941_));
  OAI210     m0913(.A0(mai_mai_n844_), .A1(mai_mai_n941_), .B0(mai_mai_n940_), .Y(mai_mai_n942_));
  NA4        m0914(.A(mai_mai_n942_), .B(mai_mai_n939_), .C(mai_mai_n938_), .D(mai_mai_n669_), .Y(mai_mai_n943_));
  NO4        m0915(.A(mai_mai_n943_), .B(mai_mai_n937_), .C(mai_mai_n928_), .D(mai_mai_n925_), .Y(mai_mai_n944_));
  NA2        m0916(.A(mai_mai_n646_), .B(mai_mai_n593_), .Y(mai_mai_n945_));
  NA4        m0917(.A(mai_mai_n945_), .B(mai_mai_n944_), .C(mai_mai_n922_), .D(mai_mai_n892_), .Y(mai01));
  NO3        m0918(.A(mai_mai_n624_), .B(mai_mai_n377_), .C(mai_mai_n235_), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n467_), .B(mai_mai_n240_), .Y(mai_mai_n948_));
  OAI210     m0920(.A0(mai_mai_n948_), .A1(mai_mai_n315_), .B0(i), .Y(mai_mai_n949_));
  NA3        m0921(.A(mai_mai_n949_), .B(mai_mai_n947_), .C(mai_mai_n792_), .Y(mai_mai_n950_));
  NA2        m0922(.A(mai_mai_n746_), .B(c), .Y(mai_mai_n951_));
  NA3        m0923(.A(mai_mai_n951_), .B(mai_mai_n705_), .C(mai_mai_n269_), .Y(mai_mai_n952_));
  INV        m0924(.A(mai_mai_n927_), .Y(mai_mai_n953_));
  AOI210     m0925(.A0(g), .A1(mai_mai_n493_), .B0(mai_mai_n953_), .Y(mai_mai_n954_));
  OA210      m0926(.A0(n), .A1(mai_mai_n296_), .B0(mai_mai_n464_), .Y(mai_mai_n955_));
  NAi41      m0927(.An(mai_mai_n135_), .B(mai_mai_n955_), .C(mai_mai_n954_), .D(mai_mai_n692_), .Y(mai_mai_n956_));
  NO2        m0928(.A(mai_mai_n524_), .B(mai_mai_n407_), .Y(mai_mai_n957_));
  NA4        m0929(.A(l), .B(g), .C(mai_mai_n43_), .D(mai_mai_n175_), .Y(mai_mai_n958_));
  OA210      m0930(.A0(mai_mai_n958_), .A1(mai_mai_n59_), .B0(mai_mai_n161_), .Y(mai_mai_n959_));
  NA3        m0931(.A(mai_mai_n959_), .B(mai_mai_n957_), .C(mai_mai_n114_), .Y(mai_mai_n960_));
  NO4        m0932(.A(mai_mai_n960_), .B(mai_mai_n956_), .C(mai_mai_n952_), .D(mai_mai_n950_), .Y(mai_mai_n961_));
  NO2        m0933(.A(n), .B(mai_mai_n168_), .Y(mai_mai_n962_));
  AOI210     m0934(.A0(mai_mai_n400_), .A1(c), .B0(mai_mai_n962_), .Y(mai_mai_n963_));
  NA3        m0935(.A(g), .B(k), .C(i), .Y(mai_mai_n964_));
  AOI210     m0936(.A0(mai_mai_n964_), .A1(mai_mai_n958_), .B0(mai_mai_n757_), .Y(mai_mai_n965_));
  INV        m0937(.A(mai_mai_n171_), .Y(mai_mai_n966_));
  NO3        m0938(.A(mai_mai_n966_), .B(mai_mai_n965_), .C(mai_mai_n896_), .Y(mai_mai_n967_));
  NA2        m0939(.A(mai_mai_n967_), .B(mai_mai_n963_), .Y(mai_mai_n968_));
  INV        m0940(.A(mai_mai_n751_), .Y(mai_mai_n969_));
  INV        m0941(.A(mai_mai_n752_), .Y(mai_mai_n970_));
  OAI210     m0942(.A0(mai_mai_n970_), .A1(mai_mai_n969_), .B0(mai_mai_n276_), .Y(mai_mai_n971_));
  NA2        m0943(.A(g), .B(mai_mai_n452_), .Y(mai_mai_n972_));
  NO3        m0944(.A(mai_mai_n65_), .B(mai_mai_n248_), .C(mai_mai_n43_), .Y(mai_mai_n973_));
  NA2        m0945(.A(mai_mai_n973_), .B(d), .Y(mai_mai_n974_));
  NA3        m0946(.A(mai_mai_n974_), .B(mai_mai_n972_), .C(mai_mai_n521_), .Y(mai_mai_n975_));
  BUFFER     m0947(.A(mai_mai_n900_), .Y(mai_mai_n976_));
  NO2        m0948(.A(mai_mai_n296_), .B(mai_mai_n59_), .Y(mai_mai_n977_));
  AOI210     m0949(.A0(g), .A1(mai_mai_n91_), .B0(mai_mai_n977_), .Y(mai_mai_n978_));
  NA2        m0950(.A(mai_mai_n973_), .B(c), .Y(mai_mai_n979_));
  NA4        m0951(.A(mai_mai_n979_), .B(mai_mai_n978_), .C(mai_mai_n976_), .D(mai_mai_n307_), .Y(mai_mai_n980_));
  NOi41      m0952(.An(mai_mai_n971_), .B(mai_mai_n980_), .C(mai_mai_n975_), .D(mai_mai_n968_), .Y(mai_mai_n981_));
  NO3        m0953(.A(mai_mai_n842_), .B(mai_mai_n146_), .C(mai_mai_n71_), .Y(mai_mai_n982_));
  NO3        m0954(.A(mai_mai_n842_), .B(mai_mai_n144_), .C(mai_mai_n71_), .Y(mai_mai_n983_));
  NO3        m0955(.A(mai_mai_n983_), .B(mai_mai_n982_), .C(mai_mai_n496_), .Y(mai_mai_n984_));
  NA3        m0956(.A(mai_mai_n984_), .B(mai_mai_n981_), .C(mai_mai_n961_), .Y(mai06));
  NO2        m0957(.A(mai_mai_n187_), .B(mai_mai_n83_), .Y(mai_mai_n986_));
  OAI210     m0958(.A0(mai_mai_n986_), .A1(mai_mai_n982_), .B0(c), .Y(mai_mai_n987_));
  NA3        m0959(.A(mai_mai_n683_), .B(mai_mai_n987_), .C(mai_mai_n971_), .Y(mai_mai_n988_));
  NO3        m0960(.A(mai_mai_n988_), .B(mai_mai_n975_), .C(mai_mai_n217_), .Y(mai_mai_n989_));
  AOI210     m0961(.A0(mai_mai_n43_), .A1(mai_mai_n43_), .B0(mai_mai_n274_), .Y(mai_mai_n990_));
  OAI210     m0962(.A0(mai_mai_n72_), .A1(mai_mai_n38_), .B0(mai_mai_n523_), .Y(mai_mai_n991_));
  NA2        m0963(.A(mai_mai_n991_), .B(mai_mai_n498_), .Y(mai_mai_n992_));
  INV        m0964(.A(mai_mai_n410_), .Y(mai_mai_n993_));
  INV        m0965(.A(mai_mai_n859_), .Y(mai_mai_n994_));
  NA2        m0966(.A(mai_mai_n208_), .B(mai_mai_n701_), .Y(mai_mai_n995_));
  NO4        m0967(.A(mai_mai_n995_), .B(mai_mai_n994_), .C(mai_mai_n113_), .D(mai_mai_n993_), .Y(mai_mai_n996_));
  OR2        m0968(.A(mai_mai_n475_), .B(mai_mai_n474_), .Y(mai_mai_n997_));
  INV        m0969(.A(mai_mai_n997_), .Y(mai_mai_n998_));
  NA3        m0970(.A(mai_mai_n998_), .B(mai_mai_n996_), .C(mai_mai_n992_), .Y(mai_mai_n999_));
  NOi21      m0971(.An(mai_mai_n172_), .B(mai_mai_n46_), .Y(mai_mai_n1000_));
  NO4        m0972(.A(mai_mai_n740_), .B(mai_mai_n1000_), .C(mai_mai_n999_), .D(mai_mai_n990_), .Y(mai_mai_n1001_));
  OAI220     m0973(.A0(mai_mai_n572_), .A1(mai_mai_n1058_), .B0(mai_mai_n187_), .B1(mai_mai_n483_), .Y(mai_mai_n1002_));
  INV        m0974(.A(mai_mai_n1002_), .Y(mai_mai_n1003_));
  NO3        m0975(.A(mai_mai_n203_), .B(mai_mai_n83_), .C(mai_mai_n237_), .Y(mai_mai_n1004_));
  OAI220     m0976(.A0(mai_mai_n1063_), .A1(mai_mai_n208_), .B0(c), .B1(mai_mai_n410_), .Y(mai_mai_n1005_));
  NOi21      m0977(.An(h), .B(mai_mai_n59_), .Y(mai_mai_n1006_));
  NO4        m0978(.A(mai_mai_n1006_), .B(mai_mai_n1005_), .C(mai_mai_n1004_), .D(mai_mai_n860_), .Y(mai_mai_n1007_));
  NAi31      m0979(.An(mai_mai_n586_), .B(mai_mai_n70_), .C(m), .Y(mai_mai_n1008_));
  NA4        m0980(.A(mai_mai_n1008_), .B(mai_mai_n1007_), .C(mai_mai_n1003_), .D(mai_mai_n939_), .Y(mai_mai_n1009_));
  OR3        m0981(.A(d), .B(mai_mai_n187_), .C(mai_mai_n483_), .Y(mai_mai_n1010_));
  AOI210     m0982(.A0(g), .A1(mai_mai_n355_), .B0(mai_mai_n298_), .Y(mai_mai_n1011_));
  NA2        m0983(.A(h), .B(mai_mai_n616_), .Y(mai_mai_n1012_));
  NA3        m0984(.A(mai_mai_n1012_), .B(mai_mai_n1011_), .C(mai_mai_n1010_), .Y(mai_mai_n1013_));
  AOI220     m0985(.A0(mai_mai_n172_), .A1(mai_mai_n593_), .B0(m), .B1(mai_mai_n198_), .Y(mai_mai_n1014_));
  NO4        m0986(.A(mai_mai_n719_), .B(mai_mai_n675_), .C(mai_mai_n396_), .D(mai_mai_n379_), .Y(mai_mai_n1015_));
  NA3        m0987(.A(mai_mai_n1015_), .B(mai_mai_n1014_), .C(mai_mai_n979_), .Y(mai_mai_n1016_));
  NAi21      m0988(.An(j), .B(i), .Y(mai_mai_n1017_));
  NO3        m0989(.A(mai_mai_n1017_), .B(mai_mai_n352_), .C(mai_mai_n195_), .Y(mai_mai_n1018_));
  NO4        m0990(.A(mai_mai_n1018_), .B(mai_mai_n1016_), .C(mai_mai_n1013_), .D(mai_mai_n1009_), .Y(mai_mai_n1019_));
  NA4        m0991(.A(mai_mai_n1019_), .B(mai_mai_n1001_), .C(mai_mai_n989_), .D(mai_mai_n984_), .Y(mai07));
  NOi31      m0992(.An(n), .B(m), .C(b), .Y(mai_mai_n1021_));
  NA3        m0993(.A(mai_mai_n539_), .B(mai_mai_n1056_), .C(mai_mai_n90_), .Y(mai_mai_n1022_));
  NO2        m0994(.A(mai_mai_n1022_), .B(mai_mai_n43_), .Y(mai_mai_n1023_));
  INV        m0995(.A(mai_mai_n1023_), .Y(mai_mai_n1024_));
  NA2        m0996(.A(mai_mai_n870_), .B(h), .Y(mai_mai_n1025_));
  NA2        m0997(.A(mai_mai_n115_), .B(mai_mai_n183_), .Y(mai_mai_n1026_));
  NO2        m0998(.A(mai_mai_n1026_), .B(mai_mai_n1025_), .Y(mai_mai_n1027_));
  INV        m0999(.A(mai_mai_n1027_), .Y(mai_mai_n1028_));
  OAI210     m1000(.A0(mai_mai_n152_), .A1(mai_mai_n421_), .B0(mai_mai_n822_), .Y(mai_mai_n1029_));
  AN2        m1001(.A(mai_mai_n1029_), .B(mai_mai_n1028_), .Y(mai_mai_n1030_));
  NO4        m1002(.A(mai_mai_n108_), .B(g), .C(f), .D(e), .Y(mai_mai_n1031_));
  NA2        m1003(.A(mai_mai_n1030_), .B(mai_mai_n1024_), .Y(mai_mai_n1032_));
  NO3        m1004(.A(mai_mai_n586_), .B(mai_mai_n144_), .C(mai_mai_n325_), .Y(mai_mai_n1033_));
  OR2        m1005(.A(n), .B(i), .Y(mai_mai_n1034_));
  OAI210     m1006(.A0(mai_mai_n1034_), .A1(mai_mai_n830_), .B0(mai_mai_n46_), .Y(mai_mai_n1035_));
  AOI220     m1007(.A0(mai_mai_n1035_), .A1(mai_mai_n901_), .B0(mai_mai_n637_), .B1(mai_mai_n160_), .Y(mai_mai_n1036_));
  NA2        m1008(.A(mai_mai_n1036_), .B(mai_mai_n1053_), .Y(mai_mai_n1037_));
  OAI210     m1009(.A0(mai_mai_n1031_), .A1(mai_mai_n1021_), .B0(mai_mai_n681_), .Y(mai_mai_n1038_));
  INV        m1010(.A(mai_mai_n1038_), .Y(mai_mai_n1039_));
  OR3        m1011(.A(mai_mai_n1039_), .B(mai_mai_n1037_), .C(mai_mai_n1032_), .Y(mai04));
  NOi31      m1012(.An(mai_mai_n1031_), .B(k), .C(mai_mai_n811_), .Y(mai_mai_n1041_));
  NO4        m1013(.A(mai_mai_n224_), .B(mai_mai_n802_), .C(mai_mai_n381_), .D(j), .Y(mai_mai_n1042_));
  OR3        m1014(.A(mai_mai_n1042_), .B(mai_mai_n1041_), .C(mai_mai_n823_), .Y(mai_mai_n1043_));
  INV        m1015(.A(mai_mai_n914_), .Y(mai_mai_n1044_));
  NA2        m1016(.A(mai_mai_n1044_), .B(mai_mai_n942_), .Y(mai_mai_n1045_));
  NO4        m1017(.A(mai_mai_n1045_), .B(mai_mai_n1043_), .C(mai_mai_n829_), .D(mai_mai_n815_), .Y(mai_mai_n1046_));
  NA4        m1018(.A(mai_mai_n1046_), .B(mai_mai_n832_), .C(mai_mai_n856_), .D(mai_mai_n849_), .Y(mai05));
  INV        m1019(.A(m), .Y(mai_mai_n1050_));
  INV        m1020(.A(m), .Y(mai_mai_n1051_));
  INV        m1021(.A(mai_mai_n539_), .Y(mai_mai_n1052_));
  INV        m1022(.A(mai_mai_n1033_), .Y(mai_mai_n1053_));
  INV        m1023(.A(mai_mai_n822_), .Y(mai_mai_n1054_));
  INV        m1024(.A(mai_mai_n183_), .Y(mai_mai_n1055_));
  INV        m1025(.A(m), .Y(mai_mai_n1056_));
  INV        m1026(.A(m), .Y(mai_mai_n1057_));
  INV        m1027(.A(g), .Y(mai_mai_n1058_));
  INV        m1028(.A(n), .Y(mai_mai_n1059_));
  INV        m1029(.A(n), .Y(mai_mai_n1060_));
  INV        m1030(.A(n), .Y(mai_mai_n1061_));
  INV        m1031(.A(n), .Y(mai_mai_n1062_));
  INV        m1032(.A(e), .Y(mai_mai_n1063_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(g), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(g), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(g), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(g), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(g), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(g), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NO2        u0066(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u0067(.A(m), .B(l), .Y(men_men_n96_));
  NAi31      u0068(.An(k), .B(j), .C(g), .Y(men_men_n97_));
  NO3        u0069(.A(men_men_n97_), .B(men_men_n96_), .C(f), .Y(men_men_n98_));
  AN2        u0070(.A(j), .B(g), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(l), .C(i), .Y(men_men_n100_));
  NOi21      u0072(.An(g), .B(i), .Y(men_men_n101_));
  NOi32      u0073(.An(m), .Bn(j), .C(k), .Y(men_men_n102_));
  AOI220     u0074(.A0(men_men_n102_), .A1(men_men_n101_), .B0(men_men_n100_), .B1(men_men_n99_), .Y(men_men_n103_));
  NO2        u0075(.A(men_men_n103_), .B(f), .Y(men_men_n104_));
  NO4        u0076(.A(men_men_n104_), .B(men_men_n98_), .C(men_men_n95_), .D(men_men_n92_), .Y(men_men_n105_));
  NAi41      u0077(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n106_));
  AN2        u0078(.A(e), .B(b), .Y(men_men_n107_));
  NOi31      u0079(.An(c), .B(h), .C(f), .Y(men_men_n108_));
  NA2        u0080(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NO3        u0081(.A(men_men_n109_), .B(men_men_n106_), .C(g), .Y(men_men_n110_));
  NOi21      u0082(.An(g), .B(f), .Y(men_men_n111_));
  NOi21      u0083(.An(i), .B(h), .Y(men_men_n112_));
  NA3        u0084(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n36_), .Y(men_men_n113_));
  INV        u0085(.A(a), .Y(men_men_n114_));
  NA2        u0086(.A(men_men_n107_), .B(men_men_n114_), .Y(men_men_n115_));
  INV        u0087(.A(l), .Y(men_men_n116_));
  NOi21      u0088(.An(m), .B(n), .Y(men_men_n117_));
  AN2        u0089(.A(k), .B(h), .Y(men_men_n118_));
  NO2        u0090(.A(men_men_n113_), .B(men_men_n88_), .Y(men_men_n119_));
  INV        u0091(.A(b), .Y(men_men_n120_));
  NA2        u0092(.A(l), .B(j), .Y(men_men_n121_));
  AN2        u0093(.A(k), .B(i), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n121_), .Y(men_men_n123_));
  NA2        u0095(.A(g), .B(e), .Y(men_men_n124_));
  NOi32      u0096(.An(c), .Bn(a), .C(d), .Y(men_men_n125_));
  NA2        u0097(.A(men_men_n125_), .B(men_men_n117_), .Y(men_men_n126_));
  NO4        u0098(.A(men_men_n126_), .B(men_men_n124_), .C(men_men_n123_), .D(men_men_n120_), .Y(men_men_n127_));
  NO3        u0099(.A(men_men_n127_), .B(men_men_n119_), .C(men_men_n110_), .Y(men_men_n128_));
  OAI210     u0100(.A0(men_men_n105_), .A1(men_men_n88_), .B0(men_men_n128_), .Y(men_men_n129_));
  NOi31      u0101(.An(k), .B(m), .C(j), .Y(men_men_n130_));
  NA3        u0102(.A(men_men_n130_), .B(men_men_n79_), .C(men_men_n78_), .Y(men_men_n131_));
  NOi31      u0103(.An(k), .B(m), .C(i), .Y(men_men_n132_));
  NA3        u0104(.A(men_men_n132_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n133_));
  NA2        u0105(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n134_));
  NOi32      u0106(.An(f), .Bn(b), .C(e), .Y(men_men_n135_));
  NAi21      u0107(.An(g), .B(h), .Y(men_men_n136_));
  NAi21      u0108(.An(m), .B(n), .Y(men_men_n137_));
  NAi21      u0109(.An(j), .B(k), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n136_), .Y(men_men_n139_));
  NAi41      u0111(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n140_));
  NAi31      u0112(.An(j), .B(k), .C(h), .Y(men_men_n141_));
  NO3        u0113(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n137_), .Y(men_men_n142_));
  AOI210     u0114(.A0(men_men_n139_), .A1(men_men_n135_), .B0(men_men_n142_), .Y(men_men_n143_));
  NO2        u0115(.A(k), .B(j), .Y(men_men_n144_));
  NO2        u0116(.A(men_men_n144_), .B(men_men_n137_), .Y(men_men_n145_));
  AN2        u0117(.A(k), .B(j), .Y(men_men_n146_));
  NAi21      u0118(.An(c), .B(b), .Y(men_men_n147_));
  NA2        u0119(.A(f), .B(d), .Y(men_men_n148_));
  NO4        u0120(.A(men_men_n148_), .B(men_men_n147_), .C(men_men_n146_), .D(men_men_n136_), .Y(men_men_n149_));
  NA2        u0121(.A(h), .B(c), .Y(men_men_n150_));
  NAi31      u0122(.An(f), .B(e), .C(b), .Y(men_men_n151_));
  NA2        u0123(.A(men_men_n149_), .B(men_men_n145_), .Y(men_men_n152_));
  NA2        u0124(.A(d), .B(b), .Y(men_men_n153_));
  NAi21      u0125(.An(e), .B(f), .Y(men_men_n154_));
  NO2        u0126(.A(men_men_n154_), .B(men_men_n153_), .Y(men_men_n155_));
  NA2        u0127(.A(b), .B(a), .Y(men_men_n156_));
  NAi21      u0128(.An(e), .B(g), .Y(men_men_n157_));
  NAi21      u0129(.An(c), .B(d), .Y(men_men_n158_));
  NAi31      u0130(.An(l), .B(k), .C(h), .Y(men_men_n159_));
  NO2        u0131(.A(men_men_n137_), .B(men_men_n159_), .Y(men_men_n160_));
  NA2        u0132(.A(men_men_n160_), .B(men_men_n155_), .Y(men_men_n161_));
  NAi41      u0133(.An(men_men_n134_), .B(men_men_n161_), .C(men_men_n152_), .D(men_men_n143_), .Y(men_men_n162_));
  NAi31      u0134(.An(e), .B(f), .C(b), .Y(men_men_n163_));
  NOi21      u0135(.An(g), .B(d), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  NOi21      u0137(.An(h), .B(i), .Y(men_men_n166_));
  NOi21      u0138(.An(k), .B(m), .Y(men_men_n167_));
  NA3        u0139(.A(men_men_n167_), .B(men_men_n166_), .C(n), .Y(men_men_n168_));
  NOi21      u0140(.An(men_men_n165_), .B(men_men_n168_), .Y(men_men_n169_));
  NOi21      u0141(.An(h), .B(g), .Y(men_men_n170_));
  NO2        u0142(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n171_));
  NA2        u0143(.A(men_men_n171_), .B(men_men_n170_), .Y(men_men_n172_));
  NAi31      u0144(.An(l), .B(j), .C(h), .Y(men_men_n173_));
  NO2        u0145(.A(men_men_n173_), .B(men_men_n49_), .Y(men_men_n174_));
  NA2        u0146(.A(men_men_n174_), .B(men_men_n67_), .Y(men_men_n175_));
  NOi32      u0147(.An(n), .Bn(k), .C(m), .Y(men_men_n176_));
  NA2        u0148(.A(l), .B(i), .Y(men_men_n177_));
  NA2        u0149(.A(men_men_n177_), .B(men_men_n176_), .Y(men_men_n178_));
  OAI210     u0150(.A0(men_men_n178_), .A1(men_men_n172_), .B0(men_men_n175_), .Y(men_men_n179_));
  NAi31      u0151(.An(d), .B(f), .C(c), .Y(men_men_n180_));
  NAi31      u0152(.An(e), .B(f), .C(c), .Y(men_men_n181_));
  NA2        u0153(.A(men_men_n181_), .B(men_men_n180_), .Y(men_men_n182_));
  NA2        u0154(.A(j), .B(h), .Y(men_men_n183_));
  OR3        u0155(.A(n), .B(m), .C(k), .Y(men_men_n184_));
  NO2        u0156(.A(men_men_n184_), .B(men_men_n183_), .Y(men_men_n185_));
  NAi32      u0157(.An(m), .Bn(k), .C(n), .Y(men_men_n186_));
  NO2        u0158(.A(men_men_n186_), .B(men_men_n183_), .Y(men_men_n187_));
  AOI220     u0159(.A0(men_men_n187_), .A1(men_men_n165_), .B0(men_men_n185_), .B1(men_men_n182_), .Y(men_men_n188_));
  NO2        u0160(.A(n), .B(m), .Y(men_men_n189_));
  NA2        u0161(.A(men_men_n189_), .B(men_men_n50_), .Y(men_men_n190_));
  NAi21      u0162(.An(f), .B(e), .Y(men_men_n191_));
  NA2        u0163(.A(d), .B(c), .Y(men_men_n192_));
  NO2        u0164(.A(men_men_n192_), .B(men_men_n191_), .Y(men_men_n193_));
  NOi21      u0165(.An(men_men_n193_), .B(men_men_n190_), .Y(men_men_n194_));
  NAi21      u0166(.An(d), .B(c), .Y(men_men_n195_));
  NAi31      u0167(.An(m), .B(n), .C(b), .Y(men_men_n196_));
  NA2        u0168(.A(k), .B(i), .Y(men_men_n197_));
  NAi21      u0169(.An(h), .B(f), .Y(men_men_n198_));
  INV        u0170(.A(men_men_n198_), .Y(men_men_n199_));
  NO2        u0171(.A(men_men_n196_), .B(men_men_n158_), .Y(men_men_n200_));
  NA2        u0172(.A(men_men_n200_), .B(men_men_n199_), .Y(men_men_n201_));
  NOi32      u0173(.An(f), .Bn(c), .C(d), .Y(men_men_n202_));
  NOi32      u0174(.An(f), .Bn(c), .C(e), .Y(men_men_n203_));
  NO2        u0175(.A(men_men_n203_), .B(men_men_n202_), .Y(men_men_n204_));
  NO3        u0176(.A(n), .B(m), .C(j), .Y(men_men_n205_));
  NA2        u0177(.A(men_men_n205_), .B(men_men_n118_), .Y(men_men_n206_));
  AO210      u0178(.A0(men_men_n206_), .A1(men_men_n190_), .B0(men_men_n204_), .Y(men_men_n207_));
  NAi41      u0179(.An(men_men_n194_), .B(men_men_n207_), .C(men_men_n201_), .D(men_men_n188_), .Y(men_men_n208_));
  OR4        u0180(.A(men_men_n208_), .B(men_men_n179_), .C(men_men_n169_), .D(men_men_n162_), .Y(men_men_n209_));
  NO4        u0181(.A(men_men_n209_), .B(men_men_n129_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n210_));
  NA3        u0182(.A(m), .B(men_men_n116_), .C(j), .Y(men_men_n211_));
  NAi31      u0183(.An(n), .B(h), .C(g), .Y(men_men_n212_));
  NO2        u0184(.A(men_men_n212_), .B(men_men_n211_), .Y(men_men_n213_));
  NOi32      u0185(.An(m), .Bn(k), .C(l), .Y(men_men_n214_));
  NA3        u0186(.A(men_men_n214_), .B(men_men_n89_), .C(g), .Y(men_men_n215_));
  NO2        u0187(.A(men_men_n215_), .B(n), .Y(men_men_n216_));
  NOi21      u0188(.An(k), .B(j), .Y(men_men_n217_));
  NA4        u0189(.A(men_men_n217_), .B(men_men_n117_), .C(i), .D(g), .Y(men_men_n218_));
  AN2        u0190(.A(i), .B(g), .Y(men_men_n219_));
  NA3        u0191(.A(men_men_n76_), .B(men_men_n219_), .C(men_men_n117_), .Y(men_men_n220_));
  NA2        u0192(.A(men_men_n220_), .B(men_men_n218_), .Y(men_men_n221_));
  NO3        u0193(.A(men_men_n221_), .B(men_men_n216_), .C(men_men_n213_), .Y(men_men_n222_));
  NAi41      u0194(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n223_));
  INV        u0195(.A(men_men_n223_), .Y(men_men_n224_));
  INV        u0196(.A(f), .Y(men_men_n225_));
  INV        u0197(.A(g), .Y(men_men_n226_));
  NOi31      u0198(.An(i), .B(j), .C(h), .Y(men_men_n227_));
  NOi21      u0199(.An(l), .B(m), .Y(men_men_n228_));
  NA2        u0200(.A(men_men_n228_), .B(men_men_n227_), .Y(men_men_n229_));
  NO3        u0201(.A(men_men_n229_), .B(men_men_n226_), .C(men_men_n225_), .Y(men_men_n230_));
  NA2        u0202(.A(men_men_n230_), .B(men_men_n224_), .Y(men_men_n231_));
  OAI210     u0203(.A0(men_men_n222_), .A1(men_men_n32_), .B0(men_men_n231_), .Y(men_men_n232_));
  NOi21      u0204(.An(n), .B(m), .Y(men_men_n233_));
  NOi32      u0205(.An(l), .Bn(i), .C(j), .Y(men_men_n234_));
  NA2        u0206(.A(men_men_n234_), .B(men_men_n233_), .Y(men_men_n235_));
  OA220      u0207(.A0(men_men_n235_), .A1(men_men_n109_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n236_));
  NAi21      u0208(.An(j), .B(h), .Y(men_men_n237_));
  XN2        u0209(.A(i), .B(h), .Y(men_men_n238_));
  NA2        u0210(.A(men_men_n238_), .B(men_men_n237_), .Y(men_men_n239_));
  NOi31      u0211(.An(k), .B(n), .C(m), .Y(men_men_n240_));
  NOi31      u0212(.An(men_men_n240_), .B(men_men_n192_), .C(men_men_n191_), .Y(men_men_n241_));
  NA2        u0213(.A(men_men_n241_), .B(men_men_n239_), .Y(men_men_n242_));
  NAi31      u0214(.An(f), .B(e), .C(c), .Y(men_men_n243_));
  NO4        u0215(.A(men_men_n243_), .B(men_men_n184_), .C(men_men_n183_), .D(men_men_n59_), .Y(men_men_n244_));
  NA4        u0216(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n245_));
  NAi32      u0217(.An(m), .Bn(i), .C(k), .Y(men_men_n246_));
  NO3        u0218(.A(men_men_n246_), .B(men_men_n93_), .C(men_men_n245_), .Y(men_men_n247_));
  NA2        u0219(.A(k), .B(h), .Y(men_men_n248_));
  NO2        u0220(.A(men_men_n247_), .B(men_men_n244_), .Y(men_men_n249_));
  NAi21      u0221(.An(n), .B(a), .Y(men_men_n250_));
  NO2        u0222(.A(men_men_n250_), .B(men_men_n153_), .Y(men_men_n251_));
  NAi41      u0223(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n252_));
  NO2        u0224(.A(men_men_n252_), .B(e), .Y(men_men_n253_));
  NO3        u0225(.A(men_men_n154_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n254_));
  OAI210     u0226(.A0(men_men_n254_), .A1(men_men_n253_), .B0(men_men_n251_), .Y(men_men_n255_));
  AN4        u0227(.A(men_men_n255_), .B(men_men_n249_), .C(men_men_n242_), .D(men_men_n236_), .Y(men_men_n256_));
  OR2        u0228(.A(h), .B(g), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n257_), .B(men_men_n106_), .Y(men_men_n258_));
  NA2        u0230(.A(men_men_n258_), .B(men_men_n135_), .Y(men_men_n259_));
  NAi41      u0231(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n260_));
  NO2        u0232(.A(men_men_n260_), .B(men_men_n225_), .Y(men_men_n261_));
  NA2        u0233(.A(men_men_n167_), .B(men_men_n112_), .Y(men_men_n262_));
  NAi21      u0234(.An(men_men_n262_), .B(men_men_n261_), .Y(men_men_n263_));
  NO2        u0235(.A(n), .B(a), .Y(men_men_n264_));
  NAi31      u0236(.An(men_men_n252_), .B(men_men_n264_), .C(men_men_n107_), .Y(men_men_n265_));
  AN2        u0237(.A(men_men_n265_), .B(men_men_n263_), .Y(men_men_n266_));
  NAi21      u0238(.An(h), .B(i), .Y(men_men_n267_));
  NA2        u0239(.A(men_men_n189_), .B(k), .Y(men_men_n268_));
  NO2        u0240(.A(men_men_n268_), .B(men_men_n267_), .Y(men_men_n269_));
  NA2        u0241(.A(men_men_n269_), .B(men_men_n202_), .Y(men_men_n270_));
  NA3        u0242(.A(men_men_n270_), .B(men_men_n266_), .C(men_men_n259_), .Y(men_men_n271_));
  NOi21      u0243(.An(g), .B(e), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n273_));
  NA2        u0245(.A(men_men_n273_), .B(men_men_n272_), .Y(men_men_n274_));
  NOi32      u0246(.An(l), .Bn(j), .C(i), .Y(men_men_n275_));
  AOI210     u0247(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n275_), .Y(men_men_n276_));
  NO2        u0248(.A(men_men_n267_), .B(men_men_n44_), .Y(men_men_n277_));
  NAi21      u0249(.An(f), .B(g), .Y(men_men_n278_));
  NO2        u0250(.A(men_men_n278_), .B(men_men_n65_), .Y(men_men_n279_));
  NO2        u0251(.A(men_men_n69_), .B(men_men_n121_), .Y(men_men_n280_));
  AOI220     u0252(.A0(men_men_n280_), .A1(men_men_n279_), .B0(men_men_n277_), .B1(men_men_n67_), .Y(men_men_n281_));
  OAI210     u0253(.A0(men_men_n276_), .A1(men_men_n274_), .B0(men_men_n281_), .Y(men_men_n282_));
  NO3        u0254(.A(men_men_n138_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n283_));
  NOi41      u0255(.An(men_men_n256_), .B(men_men_n282_), .C(men_men_n271_), .D(men_men_n232_), .Y(men_men_n284_));
  NO4        u0256(.A(men_men_n213_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n285_));
  NO2        u0257(.A(men_men_n285_), .B(men_men_n115_), .Y(men_men_n286_));
  NA3        u0258(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n287_));
  NAi21      u0259(.An(h), .B(g), .Y(men_men_n288_));
  OR4        u0260(.A(men_men_n288_), .B(men_men_n287_), .C(men_men_n235_), .D(e), .Y(men_men_n289_));
  NO2        u0261(.A(men_men_n262_), .B(men_men_n278_), .Y(men_men_n290_));
  NA2        u0262(.A(men_men_n290_), .B(men_men_n78_), .Y(men_men_n291_));
  NAi31      u0263(.An(g), .B(k), .C(h), .Y(men_men_n292_));
  NO3        u0264(.A(men_men_n137_), .B(men_men_n292_), .C(l), .Y(men_men_n293_));
  NAi31      u0265(.An(e), .B(d), .C(a), .Y(men_men_n294_));
  NA2        u0266(.A(men_men_n293_), .B(men_men_n135_), .Y(men_men_n295_));
  NA3        u0267(.A(men_men_n295_), .B(men_men_n291_), .C(men_men_n289_), .Y(men_men_n296_));
  NA4        u0268(.A(men_men_n167_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n121_), .Y(men_men_n297_));
  NA3        u0269(.A(men_men_n167_), .B(men_men_n166_), .C(men_men_n86_), .Y(men_men_n298_));
  NO2        u0270(.A(men_men_n298_), .B(men_men_n204_), .Y(men_men_n299_));
  NOi21      u0271(.An(men_men_n297_), .B(men_men_n299_), .Y(men_men_n300_));
  NA3        u0272(.A(e), .B(c), .C(b), .Y(men_men_n301_));
  NO2        u0273(.A(men_men_n60_), .B(men_men_n301_), .Y(men_men_n302_));
  NAi32      u0274(.An(k), .Bn(i), .C(j), .Y(men_men_n303_));
  NAi31      u0275(.An(h), .B(l), .C(i), .Y(men_men_n304_));
  NA3        u0276(.A(men_men_n304_), .B(men_men_n303_), .C(men_men_n173_), .Y(men_men_n305_));
  NOi21      u0277(.An(men_men_n305_), .B(men_men_n49_), .Y(men_men_n306_));
  OAI210     u0278(.A0(men_men_n279_), .A1(men_men_n302_), .B0(men_men_n306_), .Y(men_men_n307_));
  NAi21      u0279(.An(l), .B(k), .Y(men_men_n308_));
  NO2        u0280(.A(men_men_n308_), .B(men_men_n49_), .Y(men_men_n309_));
  NOi21      u0281(.An(l), .B(j), .Y(men_men_n310_));
  NA2        u0282(.A(men_men_n170_), .B(men_men_n310_), .Y(men_men_n311_));
  NA3        u0283(.A(men_men_n122_), .B(men_men_n121_), .C(g), .Y(men_men_n312_));
  OR3        u0284(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n313_));
  AOI210     u0285(.A0(men_men_n312_), .A1(men_men_n311_), .B0(men_men_n313_), .Y(men_men_n314_));
  INV        u0286(.A(men_men_n314_), .Y(men_men_n315_));
  NAi32      u0287(.An(j), .Bn(h), .C(i), .Y(men_men_n316_));
  NAi21      u0288(.An(m), .B(l), .Y(men_men_n317_));
  NO3        u0289(.A(men_men_n317_), .B(men_men_n316_), .C(men_men_n86_), .Y(men_men_n318_));
  NA2        u0290(.A(h), .B(g), .Y(men_men_n319_));
  NA2        u0291(.A(men_men_n176_), .B(men_men_n45_), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n320_), .B(men_men_n319_), .Y(men_men_n321_));
  OAI210     u0293(.A0(men_men_n321_), .A1(men_men_n318_), .B0(men_men_n171_), .Y(men_men_n322_));
  NA4        u0294(.A(men_men_n322_), .B(men_men_n315_), .C(men_men_n307_), .D(men_men_n300_), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n151_), .B(d), .Y(men_men_n324_));
  NA2        u0296(.A(men_men_n324_), .B(men_men_n53_), .Y(men_men_n325_));
  NO2        u0297(.A(men_men_n109_), .B(men_men_n106_), .Y(men_men_n326_));
  NAi32      u0298(.An(n), .Bn(m), .C(l), .Y(men_men_n327_));
  NO2        u0299(.A(men_men_n327_), .B(men_men_n316_), .Y(men_men_n328_));
  AOI220     u0300(.A0(men_men_n328_), .A1(men_men_n193_), .B0(men_men_n326_), .B1(men_men_n59_), .Y(men_men_n329_));
  NO2        u0301(.A(men_men_n126_), .B(men_men_n120_), .Y(men_men_n330_));
  NAi31      u0302(.An(k), .B(l), .C(j), .Y(men_men_n331_));
  OAI210     u0303(.A0(men_men_n308_), .A1(j), .B0(men_men_n331_), .Y(men_men_n332_));
  NOi21      u0304(.An(men_men_n332_), .B(men_men_n124_), .Y(men_men_n333_));
  NA2        u0305(.A(men_men_n333_), .B(men_men_n330_), .Y(men_men_n334_));
  NA3        u0306(.A(men_men_n334_), .B(men_men_n329_), .C(men_men_n325_), .Y(men_men_n335_));
  NO4        u0307(.A(men_men_n335_), .B(men_men_n323_), .C(men_men_n296_), .D(men_men_n286_), .Y(men_men_n336_));
  NA2        u0308(.A(men_men_n269_), .B(men_men_n203_), .Y(men_men_n337_));
  NAi21      u0309(.An(m), .B(k), .Y(men_men_n338_));
  NO2        u0310(.A(men_men_n238_), .B(men_men_n338_), .Y(men_men_n339_));
  NAi41      u0311(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n340_));
  NO2        u0312(.A(men_men_n340_), .B(men_men_n157_), .Y(men_men_n341_));
  NA2        u0313(.A(men_men_n341_), .B(men_men_n339_), .Y(men_men_n342_));
  NAi31      u0314(.An(i), .B(l), .C(h), .Y(men_men_n343_));
  NO4        u0315(.A(men_men_n343_), .B(men_men_n157_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n344_));
  NA2        u0316(.A(e), .B(c), .Y(men_men_n345_));
  NO3        u0317(.A(men_men_n345_), .B(n), .C(d), .Y(men_men_n346_));
  NOi21      u0318(.An(f), .B(h), .Y(men_men_n347_));
  NA2        u0319(.A(men_men_n347_), .B(men_men_n122_), .Y(men_men_n348_));
  NO2        u0320(.A(men_men_n348_), .B(men_men_n226_), .Y(men_men_n349_));
  NAi31      u0321(.An(d), .B(e), .C(b), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n137_), .B(men_men_n350_), .Y(men_men_n351_));
  NA2        u0323(.A(men_men_n351_), .B(men_men_n349_), .Y(men_men_n352_));
  NAi41      u0324(.An(men_men_n344_), .B(men_men_n352_), .C(men_men_n342_), .D(men_men_n337_), .Y(men_men_n353_));
  NO4        u0325(.A(men_men_n340_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n226_), .Y(men_men_n354_));
  NA2        u0326(.A(men_men_n264_), .B(men_men_n107_), .Y(men_men_n355_));
  OR2        u0327(.A(men_men_n355_), .B(men_men_n215_), .Y(men_men_n356_));
  NOi31      u0328(.An(l), .B(n), .C(m), .Y(men_men_n357_));
  NA2        u0329(.A(men_men_n357_), .B(men_men_n227_), .Y(men_men_n358_));
  NO2        u0330(.A(men_men_n358_), .B(men_men_n204_), .Y(men_men_n359_));
  NAi32      u0331(.An(men_men_n359_), .Bn(men_men_n354_), .C(men_men_n356_), .Y(men_men_n360_));
  NAi32      u0332(.An(m), .Bn(j), .C(k), .Y(men_men_n361_));
  NAi41      u0333(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n362_));
  OAI210     u0334(.A0(men_men_n223_), .A1(men_men_n361_), .B0(men_men_n362_), .Y(men_men_n363_));
  NOi31      u0335(.An(j), .B(m), .C(k), .Y(men_men_n364_));
  NO2        u0336(.A(men_men_n130_), .B(men_men_n364_), .Y(men_men_n365_));
  AN3        u0337(.A(h), .B(g), .C(f), .Y(men_men_n366_));
  NAi31      u0338(.An(men_men_n365_), .B(men_men_n366_), .C(men_men_n363_), .Y(men_men_n367_));
  NOi32      u0339(.An(m), .Bn(j), .C(l), .Y(men_men_n368_));
  NO2        u0340(.A(men_men_n368_), .B(men_men_n100_), .Y(men_men_n369_));
  NAi32      u0341(.An(men_men_n369_), .Bn(men_men_n212_), .C(men_men_n324_), .Y(men_men_n370_));
  NO2        u0342(.A(men_men_n317_), .B(men_men_n316_), .Y(men_men_n371_));
  NO2        u0343(.A(men_men_n229_), .B(g), .Y(men_men_n372_));
  NO2        u0344(.A(men_men_n163_), .B(men_men_n86_), .Y(men_men_n373_));
  AOI220     u0345(.A0(men_men_n373_), .A1(men_men_n372_), .B0(men_men_n261_), .B1(men_men_n371_), .Y(men_men_n374_));
  NA2        u0346(.A(men_men_n246_), .B(men_men_n81_), .Y(men_men_n375_));
  NA3        u0347(.A(men_men_n375_), .B(men_men_n366_), .C(men_men_n224_), .Y(men_men_n376_));
  NA4        u0348(.A(men_men_n376_), .B(men_men_n374_), .C(men_men_n370_), .D(men_men_n367_), .Y(men_men_n377_));
  NA3        u0349(.A(h), .B(g), .C(f), .Y(men_men_n378_));
  NO2        u0350(.A(men_men_n378_), .B(men_men_n77_), .Y(men_men_n379_));
  NA2        u0351(.A(men_men_n362_), .B(men_men_n223_), .Y(men_men_n380_));
  NA2        u0352(.A(men_men_n170_), .B(e), .Y(men_men_n381_));
  NO2        u0353(.A(men_men_n381_), .B(men_men_n41_), .Y(men_men_n382_));
  AOI220     u0354(.A0(men_men_n382_), .A1(men_men_n330_), .B0(men_men_n380_), .B1(men_men_n379_), .Y(men_men_n383_));
  NOi32      u0355(.An(j), .Bn(g), .C(i), .Y(men_men_n384_));
  NA3        u0356(.A(men_men_n384_), .B(men_men_n308_), .C(men_men_n117_), .Y(men_men_n385_));
  AO210      u0357(.A0(men_men_n115_), .A1(men_men_n32_), .B0(men_men_n385_), .Y(men_men_n386_));
  NOi32      u0358(.An(e), .Bn(b), .C(a), .Y(men_men_n387_));
  AN2        u0359(.A(l), .B(j), .Y(men_men_n388_));
  NO2        u0360(.A(men_men_n338_), .B(men_men_n388_), .Y(men_men_n389_));
  NO3        u0361(.A(men_men_n340_), .B(men_men_n72_), .C(men_men_n226_), .Y(men_men_n390_));
  NA3        u0362(.A(men_men_n220_), .B(men_men_n218_), .C(men_men_n35_), .Y(men_men_n391_));
  AOI220     u0363(.A0(men_men_n391_), .A1(men_men_n387_), .B0(men_men_n390_), .B1(men_men_n389_), .Y(men_men_n392_));
  NO2        u0364(.A(men_men_n350_), .B(n), .Y(men_men_n393_));
  NA2        u0365(.A(men_men_n219_), .B(k), .Y(men_men_n394_));
  NA3        u0366(.A(m), .B(men_men_n116_), .C(men_men_n225_), .Y(men_men_n395_));
  NA4        u0367(.A(men_men_n214_), .B(men_men_n89_), .C(g), .D(men_men_n225_), .Y(men_men_n396_));
  OAI210     u0368(.A0(men_men_n395_), .A1(men_men_n394_), .B0(men_men_n396_), .Y(men_men_n397_));
  NAi41      u0369(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n398_));
  NA2        u0370(.A(men_men_n51_), .B(men_men_n117_), .Y(men_men_n399_));
  NO2        u0371(.A(men_men_n399_), .B(men_men_n398_), .Y(men_men_n400_));
  AOI220     u0372(.A0(men_men_n400_), .A1(b), .B0(men_men_n397_), .B1(men_men_n393_), .Y(men_men_n401_));
  NA4        u0373(.A(men_men_n401_), .B(men_men_n392_), .C(men_men_n386_), .D(men_men_n383_), .Y(men_men_n402_));
  NO4        u0374(.A(men_men_n402_), .B(men_men_n377_), .C(men_men_n360_), .D(men_men_n353_), .Y(men_men_n403_));
  NA4        u0375(.A(men_men_n403_), .B(men_men_n336_), .C(men_men_n284_), .D(men_men_n210_), .Y(men10));
  NA3        u0376(.A(m), .B(k), .C(i), .Y(men_men_n405_));
  NO3        u0377(.A(men_men_n405_), .B(j), .C(men_men_n226_), .Y(men_men_n406_));
  NOi21      u0378(.An(e), .B(f), .Y(men_men_n407_));
  NO4        u0379(.A(men_men_n158_), .B(men_men_n407_), .C(n), .D(men_men_n114_), .Y(men_men_n408_));
  NAi31      u0380(.An(b), .B(f), .C(c), .Y(men_men_n409_));
  INV        u0381(.A(men_men_n409_), .Y(men_men_n410_));
  NOi32      u0382(.An(k), .Bn(h), .C(j), .Y(men_men_n411_));
  NA2        u0383(.A(men_men_n411_), .B(men_men_n233_), .Y(men_men_n412_));
  NA2        u0384(.A(men_men_n168_), .B(men_men_n412_), .Y(men_men_n413_));
  AOI220     u0385(.A0(men_men_n413_), .A1(men_men_n410_), .B0(men_men_n408_), .B1(men_men_n406_), .Y(men_men_n414_));
  AN2        u0386(.A(j), .B(h), .Y(men_men_n415_));
  NO3        u0387(.A(n), .B(m), .C(k), .Y(men_men_n416_));
  NA2        u0388(.A(men_men_n416_), .B(men_men_n415_), .Y(men_men_n417_));
  NO3        u0389(.A(men_men_n417_), .B(men_men_n158_), .C(men_men_n225_), .Y(men_men_n418_));
  OR2        u0390(.A(m), .B(k), .Y(men_men_n419_));
  NO2        u0391(.A(men_men_n183_), .B(men_men_n419_), .Y(men_men_n420_));
  NA4        u0392(.A(n), .B(f), .C(c), .D(men_men_n120_), .Y(men_men_n421_));
  NOi21      u0393(.An(men_men_n420_), .B(men_men_n421_), .Y(men_men_n422_));
  NOi32      u0394(.An(d), .Bn(a), .C(c), .Y(men_men_n423_));
  NA2        u0395(.A(men_men_n423_), .B(men_men_n191_), .Y(men_men_n424_));
  NAi21      u0396(.An(i), .B(g), .Y(men_men_n425_));
  NAi31      u0397(.An(k), .B(m), .C(j), .Y(men_men_n426_));
  NO3        u0398(.A(men_men_n426_), .B(men_men_n425_), .C(n), .Y(men_men_n427_));
  NOi21      u0399(.An(men_men_n427_), .B(men_men_n424_), .Y(men_men_n428_));
  NO3        u0400(.A(men_men_n428_), .B(men_men_n422_), .C(men_men_n418_), .Y(men_men_n429_));
  NO2        u0401(.A(men_men_n421_), .B(men_men_n317_), .Y(men_men_n430_));
  NOi32      u0402(.An(f), .Bn(d), .C(c), .Y(men_men_n431_));
  AOI220     u0403(.A0(men_men_n431_), .A1(men_men_n328_), .B0(men_men_n430_), .B1(men_men_n227_), .Y(men_men_n432_));
  NA3        u0404(.A(men_men_n432_), .B(men_men_n429_), .C(men_men_n414_), .Y(men_men_n433_));
  NO2        u0405(.A(men_men_n59_), .B(men_men_n120_), .Y(men_men_n434_));
  NA2        u0406(.A(men_men_n264_), .B(men_men_n434_), .Y(men_men_n435_));
  INV        u0407(.A(e), .Y(men_men_n436_));
  NA2        u0408(.A(men_men_n46_), .B(e), .Y(men_men_n437_));
  OAI220     u0409(.A0(men_men_n437_), .A1(men_men_n211_), .B0(men_men_n215_), .B1(men_men_n436_), .Y(men_men_n438_));
  AN2        u0410(.A(g), .B(e), .Y(men_men_n439_));
  NA3        u0411(.A(men_men_n439_), .B(men_men_n214_), .C(i), .Y(men_men_n440_));
  OAI210     u0412(.A0(men_men_n91_), .A1(men_men_n436_), .B0(men_men_n440_), .Y(men_men_n441_));
  NO2        u0413(.A(men_men_n103_), .B(men_men_n436_), .Y(men_men_n442_));
  NO3        u0414(.A(men_men_n442_), .B(men_men_n441_), .C(men_men_n438_), .Y(men_men_n443_));
  NOi32      u0415(.An(h), .Bn(e), .C(g), .Y(men_men_n444_));
  NA3        u0416(.A(men_men_n444_), .B(men_men_n310_), .C(m), .Y(men_men_n445_));
  NOi21      u0417(.An(g), .B(h), .Y(men_men_n446_));
  AN3        u0418(.A(m), .B(l), .C(i), .Y(men_men_n447_));
  NA3        u0419(.A(men_men_n447_), .B(men_men_n446_), .C(e), .Y(men_men_n448_));
  AN3        u0420(.A(h), .B(g), .C(e), .Y(men_men_n449_));
  NA2        u0421(.A(men_men_n449_), .B(men_men_n100_), .Y(men_men_n450_));
  AN3        u0422(.A(men_men_n450_), .B(men_men_n448_), .C(men_men_n445_), .Y(men_men_n451_));
  AOI210     u0423(.A0(men_men_n451_), .A1(men_men_n443_), .B0(men_men_n435_), .Y(men_men_n452_));
  NA3        u0424(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n453_));
  NO2        u0425(.A(men_men_n453_), .B(men_men_n435_), .Y(men_men_n454_));
  NA3        u0426(.A(men_men_n423_), .B(men_men_n191_), .C(men_men_n86_), .Y(men_men_n455_));
  NAi31      u0427(.An(b), .B(c), .C(a), .Y(men_men_n456_));
  NO2        u0428(.A(men_men_n456_), .B(n), .Y(men_men_n457_));
  OAI210     u0429(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n458_));
  NO2        u0430(.A(men_men_n458_), .B(men_men_n154_), .Y(men_men_n459_));
  NA2        u0431(.A(men_men_n459_), .B(men_men_n457_), .Y(men_men_n460_));
  INV        u0432(.A(men_men_n460_), .Y(men_men_n461_));
  NO4        u0433(.A(men_men_n461_), .B(men_men_n454_), .C(men_men_n452_), .D(men_men_n433_), .Y(men_men_n462_));
  NA2        u0434(.A(i), .B(g), .Y(men_men_n463_));
  NO3        u0435(.A(men_men_n294_), .B(men_men_n463_), .C(c), .Y(men_men_n464_));
  NOi21      u0436(.An(a), .B(n), .Y(men_men_n465_));
  NOi21      u0437(.An(d), .B(c), .Y(men_men_n466_));
  NA2        u0438(.A(men_men_n466_), .B(men_men_n465_), .Y(men_men_n467_));
  NA3        u0439(.A(i), .B(g), .C(f), .Y(men_men_n468_));
  OR2        u0440(.A(men_men_n468_), .B(men_men_n71_), .Y(men_men_n469_));
  NA3        u0441(.A(men_men_n447_), .B(men_men_n446_), .C(men_men_n191_), .Y(men_men_n470_));
  AOI210     u0442(.A0(men_men_n470_), .A1(men_men_n469_), .B0(men_men_n467_), .Y(men_men_n471_));
  AOI210     u0443(.A0(men_men_n464_), .A1(men_men_n309_), .B0(men_men_n471_), .Y(men_men_n472_));
  OR2        u0444(.A(n), .B(m), .Y(men_men_n473_));
  NO2        u0445(.A(men_men_n473_), .B(men_men_n159_), .Y(men_men_n474_));
  NO2        u0446(.A(men_men_n192_), .B(men_men_n154_), .Y(men_men_n475_));
  OAI210     u0447(.A0(men_men_n474_), .A1(men_men_n185_), .B0(men_men_n475_), .Y(men_men_n476_));
  INV        u0448(.A(men_men_n399_), .Y(men_men_n477_));
  NA3        u0449(.A(men_men_n477_), .B(men_men_n387_), .C(d), .Y(men_men_n478_));
  NO2        u0450(.A(men_men_n456_), .B(men_men_n49_), .Y(men_men_n479_));
  NO3        u0451(.A(men_men_n66_), .B(men_men_n116_), .C(e), .Y(men_men_n480_));
  NAi21      u0452(.An(k), .B(j), .Y(men_men_n481_));
  NA2        u0453(.A(men_men_n267_), .B(men_men_n481_), .Y(men_men_n482_));
  NA3        u0454(.A(men_men_n482_), .B(men_men_n480_), .C(men_men_n479_), .Y(men_men_n483_));
  NAi21      u0455(.An(e), .B(d), .Y(men_men_n484_));
  NO2        u0456(.A(men_men_n484_), .B(men_men_n56_), .Y(men_men_n485_));
  NO2        u0457(.A(men_men_n268_), .B(men_men_n225_), .Y(men_men_n486_));
  NA3        u0458(.A(men_men_n486_), .B(men_men_n485_), .C(men_men_n239_), .Y(men_men_n487_));
  NA4        u0459(.A(men_men_n487_), .B(men_men_n483_), .C(men_men_n478_), .D(men_men_n476_), .Y(men_men_n488_));
  NO2        u0460(.A(men_men_n358_), .B(men_men_n225_), .Y(men_men_n489_));
  NA2        u0461(.A(men_men_n489_), .B(men_men_n485_), .Y(men_men_n490_));
  NOi31      u0462(.An(n), .B(m), .C(k), .Y(men_men_n491_));
  AOI220     u0463(.A0(men_men_n491_), .A1(men_men_n415_), .B0(men_men_n233_), .B1(men_men_n50_), .Y(men_men_n492_));
  NAi31      u0464(.An(g), .B(f), .C(c), .Y(men_men_n493_));
  OR3        u0465(.A(men_men_n493_), .B(men_men_n492_), .C(e), .Y(men_men_n494_));
  NA3        u0466(.A(men_men_n494_), .B(men_men_n490_), .C(men_men_n329_), .Y(men_men_n495_));
  NOi41      u0467(.An(men_men_n472_), .B(men_men_n495_), .C(men_men_n488_), .D(men_men_n282_), .Y(men_men_n496_));
  NOi32      u0468(.An(c), .Bn(a), .C(b), .Y(men_men_n497_));
  NA2        u0469(.A(men_men_n497_), .B(men_men_n117_), .Y(men_men_n498_));
  NA2        u0470(.A(men_men_n292_), .B(men_men_n159_), .Y(men_men_n499_));
  AN2        u0471(.A(e), .B(d), .Y(men_men_n500_));
  NA2        u0472(.A(men_men_n500_), .B(men_men_n499_), .Y(men_men_n501_));
  INV        u0473(.A(men_men_n154_), .Y(men_men_n502_));
  NO2        u0474(.A(men_men_n136_), .B(men_men_n41_), .Y(men_men_n503_));
  NO2        u0475(.A(men_men_n66_), .B(e), .Y(men_men_n504_));
  NOi31      u0476(.An(j), .B(k), .C(i), .Y(men_men_n505_));
  NOi21      u0477(.An(men_men_n173_), .B(men_men_n505_), .Y(men_men_n506_));
  NA4        u0478(.A(men_men_n343_), .B(men_men_n506_), .C(men_men_n276_), .D(men_men_n123_), .Y(men_men_n507_));
  AOI220     u0479(.A0(men_men_n507_), .A1(men_men_n504_), .B0(men_men_n503_), .B1(men_men_n502_), .Y(men_men_n508_));
  AOI210     u0480(.A0(men_men_n508_), .A1(men_men_n501_), .B0(men_men_n498_), .Y(men_men_n509_));
  NO2        u0481(.A(men_men_n221_), .B(men_men_n216_), .Y(men_men_n510_));
  NOi21      u0482(.An(a), .B(b), .Y(men_men_n511_));
  NA3        u0483(.A(e), .B(d), .C(c), .Y(men_men_n512_));
  NAi21      u0484(.An(men_men_n512_), .B(men_men_n511_), .Y(men_men_n513_));
  NO2        u0485(.A(men_men_n455_), .B(men_men_n215_), .Y(men_men_n514_));
  NOi21      u0486(.An(men_men_n513_), .B(men_men_n514_), .Y(men_men_n515_));
  AOI210     u0487(.A0(men_men_n285_), .A1(men_men_n510_), .B0(men_men_n515_), .Y(men_men_n516_));
  NO4        u0488(.A(men_men_n198_), .B(men_men_n106_), .C(men_men_n56_), .D(b), .Y(men_men_n517_));
  NA2        u0489(.A(men_men_n410_), .B(men_men_n160_), .Y(men_men_n518_));
  OR2        u0490(.A(k), .B(j), .Y(men_men_n519_));
  NA2        u0491(.A(l), .B(k), .Y(men_men_n520_));
  NA3        u0492(.A(men_men_n520_), .B(men_men_n519_), .C(men_men_n233_), .Y(men_men_n521_));
  AOI210     u0493(.A0(men_men_n246_), .A1(men_men_n361_), .B0(men_men_n86_), .Y(men_men_n522_));
  NOi21      u0494(.An(men_men_n521_), .B(men_men_n522_), .Y(men_men_n523_));
  OR3        u0495(.A(men_men_n523_), .B(men_men_n150_), .C(men_men_n140_), .Y(men_men_n524_));
  NA3        u0496(.A(men_men_n297_), .B(men_men_n133_), .C(men_men_n131_), .Y(men_men_n525_));
  NA2        u0497(.A(men_men_n423_), .B(men_men_n117_), .Y(men_men_n526_));
  NO4        u0498(.A(men_men_n526_), .B(men_men_n97_), .C(men_men_n116_), .D(e), .Y(men_men_n527_));
  NO3        u0499(.A(men_men_n455_), .B(men_men_n94_), .C(men_men_n136_), .Y(men_men_n528_));
  NO4        u0500(.A(men_men_n528_), .B(men_men_n527_), .C(men_men_n525_), .D(men_men_n344_), .Y(men_men_n529_));
  NA3        u0501(.A(men_men_n529_), .B(men_men_n524_), .C(men_men_n518_), .Y(men_men_n530_));
  NO4        u0502(.A(men_men_n530_), .B(men_men_n517_), .C(men_men_n516_), .D(men_men_n509_), .Y(men_men_n531_));
  NA2        u0503(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n532_));
  NOi21      u0504(.An(d), .B(e), .Y(men_men_n533_));
  NO2        u0505(.A(men_men_n198_), .B(men_men_n56_), .Y(men_men_n534_));
  NAi31      u0506(.An(j), .B(l), .C(i), .Y(men_men_n535_));
  NA4        u0507(.A(n), .B(men_men_n534_), .C(men_men_n533_), .D(b), .Y(men_men_n536_));
  NO3        u0508(.A(men_men_n424_), .B(men_men_n369_), .C(men_men_n212_), .Y(men_men_n537_));
  NO2        u0509(.A(men_men_n424_), .B(men_men_n399_), .Y(men_men_n538_));
  NO4        u0510(.A(men_men_n538_), .B(men_men_n537_), .C(men_men_n194_), .D(men_men_n326_), .Y(men_men_n539_));
  NA4        u0511(.A(men_men_n539_), .B(men_men_n536_), .C(men_men_n532_), .D(men_men_n256_), .Y(men_men_n540_));
  OAI210     u0512(.A0(men_men_n132_), .A1(men_men_n130_), .B0(n), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n541_), .B(men_men_n136_), .Y(men_men_n542_));
  AO210      u0514(.A0(men_men_n318_), .A1(men_men_n226_), .B0(men_men_n258_), .Y(men_men_n543_));
  OA210      u0515(.A0(men_men_n543_), .A1(men_men_n542_), .B0(men_men_n203_), .Y(men_men_n544_));
  XO2        u0516(.A(i), .B(h), .Y(men_men_n545_));
  NA3        u0517(.A(men_men_n545_), .B(men_men_n167_), .C(n), .Y(men_men_n546_));
  NAi41      u0518(.An(men_men_n318_), .B(men_men_n546_), .C(men_men_n492_), .D(men_men_n412_), .Y(men_men_n547_));
  NOi32      u0519(.An(men_men_n547_), .Bn(men_men_n504_), .C(men_men_n287_), .Y(men_men_n548_));
  NAi31      u0520(.An(c), .B(f), .C(d), .Y(men_men_n549_));
  AOI210     u0521(.A0(men_men_n298_), .A1(men_men_n206_), .B0(men_men_n549_), .Y(men_men_n550_));
  NOi21      u0522(.An(men_men_n84_), .B(men_men_n550_), .Y(men_men_n551_));
  NA3        u0523(.A(men_men_n408_), .B(men_men_n100_), .C(men_men_n99_), .Y(men_men_n552_));
  NA2        u0524(.A(men_men_n240_), .B(men_men_n112_), .Y(men_men_n553_));
  AOI210     u0525(.A0(men_men_n553_), .A1(men_men_n190_), .B0(men_men_n549_), .Y(men_men_n554_));
  AOI210     u0526(.A0(men_men_n385_), .A1(men_men_n35_), .B0(men_men_n513_), .Y(men_men_n555_));
  NOi31      u0527(.An(men_men_n552_), .B(men_men_n555_), .C(men_men_n554_), .Y(men_men_n556_));
  AO220      u0528(.A0(men_men_n306_), .A1(men_men_n279_), .B0(men_men_n174_), .B1(men_men_n67_), .Y(men_men_n557_));
  NA3        u0529(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n558_));
  NO2        u0530(.A(men_men_n558_), .B(men_men_n467_), .Y(men_men_n559_));
  NO2        u0531(.A(men_men_n559_), .B(men_men_n314_), .Y(men_men_n560_));
  NAi41      u0532(.An(men_men_n557_), .B(men_men_n560_), .C(men_men_n556_), .D(men_men_n551_), .Y(men_men_n561_));
  NO4        u0533(.A(men_men_n561_), .B(men_men_n548_), .C(men_men_n544_), .D(men_men_n540_), .Y(men_men_n562_));
  NA4        u0534(.A(men_men_n562_), .B(men_men_n531_), .C(men_men_n496_), .D(men_men_n462_), .Y(men11));
  NO2        u0535(.A(men_men_n73_), .B(f), .Y(men_men_n564_));
  NA2        u0536(.A(j), .B(g), .Y(men_men_n565_));
  NAi31      u0537(.An(i), .B(m), .C(l), .Y(men_men_n566_));
  NA3        u0538(.A(m), .B(k), .C(j), .Y(men_men_n567_));
  OAI220     u0539(.A0(men_men_n567_), .A1(men_men_n136_), .B0(men_men_n566_), .B1(men_men_n565_), .Y(men_men_n568_));
  NA2        u0540(.A(men_men_n568_), .B(men_men_n564_), .Y(men_men_n569_));
  NOi32      u0541(.An(e), .Bn(b), .C(f), .Y(men_men_n570_));
  NA2        u0542(.A(men_men_n275_), .B(men_men_n117_), .Y(men_men_n571_));
  NA2        u0543(.A(men_men_n46_), .B(j), .Y(men_men_n572_));
  OAI220     u0544(.A0(men_men_n572_), .A1(men_men_n320_), .B0(men_men_n571_), .B1(men_men_n226_), .Y(men_men_n573_));
  NAi31      u0545(.An(d), .B(e), .C(a), .Y(men_men_n574_));
  NO2        u0546(.A(men_men_n574_), .B(n), .Y(men_men_n575_));
  AOI220     u0547(.A0(men_men_n575_), .A1(men_men_n104_), .B0(men_men_n573_), .B1(men_men_n570_), .Y(men_men_n576_));
  NAi41      u0548(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n577_));
  AN2        u0549(.A(men_men_n577_), .B(men_men_n398_), .Y(men_men_n578_));
  AOI210     u0550(.A0(men_men_n578_), .A1(men_men_n424_), .B0(men_men_n288_), .Y(men_men_n579_));
  NA2        u0551(.A(j), .B(i), .Y(men_men_n580_));
  NAi31      u0552(.An(n), .B(m), .C(k), .Y(men_men_n581_));
  NO3        u0553(.A(men_men_n581_), .B(men_men_n580_), .C(men_men_n116_), .Y(men_men_n582_));
  NO4        u0554(.A(n), .B(d), .C(men_men_n120_), .D(a), .Y(men_men_n583_));
  NO2        u0555(.A(c), .B(men_men_n156_), .Y(men_men_n584_));
  NO2        u0556(.A(men_men_n584_), .B(men_men_n583_), .Y(men_men_n585_));
  NOi32      u0557(.An(g), .Bn(f), .C(i), .Y(men_men_n586_));
  AOI220     u0558(.A0(men_men_n586_), .A1(men_men_n102_), .B0(men_men_n568_), .B1(f), .Y(men_men_n587_));
  NO2        u0559(.A(men_men_n292_), .B(men_men_n49_), .Y(men_men_n588_));
  NO2        u0560(.A(men_men_n587_), .B(men_men_n585_), .Y(men_men_n589_));
  AOI210     u0561(.A0(men_men_n582_), .A1(men_men_n579_), .B0(men_men_n589_), .Y(men_men_n590_));
  NA2        u0562(.A(men_men_n146_), .B(men_men_n34_), .Y(men_men_n591_));
  OAI220     u0563(.A0(men_men_n591_), .A1(m), .B0(men_men_n572_), .B1(men_men_n246_), .Y(men_men_n592_));
  NOi41      u0564(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n593_));
  NAi32      u0565(.An(e), .Bn(b), .C(c), .Y(men_men_n594_));
  OR2        u0566(.A(men_men_n594_), .B(men_men_n86_), .Y(men_men_n595_));
  AN2        u0567(.A(men_men_n362_), .B(men_men_n340_), .Y(men_men_n596_));
  NA2        u0568(.A(men_men_n596_), .B(men_men_n595_), .Y(men_men_n597_));
  OA210      u0569(.A0(men_men_n597_), .A1(men_men_n593_), .B0(men_men_n592_), .Y(men_men_n598_));
  OAI220     u0570(.A0(men_men_n426_), .A1(men_men_n425_), .B0(men_men_n566_), .B1(men_men_n565_), .Y(men_men_n599_));
  NAi31      u0571(.An(d), .B(c), .C(a), .Y(men_men_n600_));
  NO2        u0572(.A(men_men_n600_), .B(n), .Y(men_men_n601_));
  NA3        u0573(.A(men_men_n601_), .B(men_men_n599_), .C(e), .Y(men_men_n602_));
  NO3        u0574(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n226_), .Y(men_men_n603_));
  NO2        u0575(.A(men_men_n243_), .B(men_men_n114_), .Y(men_men_n604_));
  OAI210     u0576(.A0(men_men_n603_), .A1(men_men_n427_), .B0(men_men_n604_), .Y(men_men_n605_));
  NA2        u0577(.A(men_men_n605_), .B(men_men_n602_), .Y(men_men_n606_));
  NO2        u0578(.A(men_men_n294_), .B(n), .Y(men_men_n607_));
  NO2        u0579(.A(men_men_n457_), .B(men_men_n607_), .Y(men_men_n608_));
  NA2        u0580(.A(men_men_n599_), .B(f), .Y(men_men_n609_));
  NAi32      u0581(.An(d), .Bn(a), .C(b), .Y(men_men_n610_));
  NO2        u0582(.A(men_men_n610_), .B(men_men_n49_), .Y(men_men_n611_));
  NA2        u0583(.A(h), .B(f), .Y(men_men_n612_));
  NO2        u0584(.A(men_men_n612_), .B(men_men_n97_), .Y(men_men_n613_));
  NO3        u0585(.A(men_men_n186_), .B(men_men_n183_), .C(g), .Y(men_men_n614_));
  AOI220     u0586(.A0(men_men_n614_), .A1(men_men_n58_), .B0(men_men_n613_), .B1(men_men_n611_), .Y(men_men_n615_));
  OAI210     u0587(.A0(men_men_n609_), .A1(men_men_n608_), .B0(men_men_n615_), .Y(men_men_n616_));
  AN3        u0588(.A(j), .B(h), .C(g), .Y(men_men_n617_));
  NO2        u0589(.A(men_men_n153_), .B(c), .Y(men_men_n618_));
  NA3        u0590(.A(men_men_n618_), .B(men_men_n617_), .C(men_men_n491_), .Y(men_men_n619_));
  NA3        u0591(.A(f), .B(d), .C(b), .Y(men_men_n620_));
  NO4        u0592(.A(men_men_n620_), .B(men_men_n186_), .C(men_men_n183_), .D(g), .Y(men_men_n621_));
  NAi21      u0593(.An(men_men_n621_), .B(men_men_n619_), .Y(men_men_n622_));
  NO4        u0594(.A(men_men_n622_), .B(men_men_n616_), .C(men_men_n606_), .D(men_men_n598_), .Y(men_men_n623_));
  AN4        u0595(.A(men_men_n623_), .B(men_men_n590_), .C(men_men_n576_), .D(men_men_n569_), .Y(men_men_n624_));
  INV        u0596(.A(k), .Y(men_men_n625_));
  NA3        u0597(.A(l), .B(men_men_n625_), .C(i), .Y(men_men_n626_));
  INV        u0598(.A(men_men_n626_), .Y(men_men_n627_));
  NA4        u0599(.A(men_men_n423_), .B(men_men_n446_), .C(men_men_n191_), .D(men_men_n117_), .Y(men_men_n628_));
  NAi32      u0600(.An(h), .Bn(f), .C(g), .Y(men_men_n629_));
  NAi41      u0601(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n630_));
  OAI210     u0602(.A0(men_men_n574_), .A1(n), .B0(men_men_n630_), .Y(men_men_n631_));
  NA2        u0603(.A(men_men_n631_), .B(m), .Y(men_men_n632_));
  NAi31      u0604(.An(h), .B(g), .C(f), .Y(men_men_n633_));
  OR3        u0605(.A(men_men_n633_), .B(men_men_n294_), .C(men_men_n49_), .Y(men_men_n634_));
  NA4        u0606(.A(men_men_n446_), .B(men_men_n125_), .C(men_men_n117_), .D(e), .Y(men_men_n635_));
  AN2        u0607(.A(men_men_n635_), .B(men_men_n634_), .Y(men_men_n636_));
  OA210      u0608(.A0(men_men_n632_), .A1(men_men_n629_), .B0(men_men_n636_), .Y(men_men_n637_));
  NO3        u0609(.A(men_men_n629_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n638_));
  NO4        u0610(.A(men_men_n633_), .B(c), .C(men_men_n156_), .D(men_men_n75_), .Y(men_men_n639_));
  OR2        u0611(.A(men_men_n639_), .B(men_men_n638_), .Y(men_men_n640_));
  NAi31      u0612(.An(men_men_n640_), .B(men_men_n637_), .C(men_men_n628_), .Y(men_men_n641_));
  NAi31      u0613(.An(f), .B(h), .C(g), .Y(men_men_n642_));
  NO4        u0614(.A(men_men_n331_), .B(men_men_n642_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n643_));
  NOi32      u0615(.An(b), .Bn(a), .C(c), .Y(men_men_n644_));
  NOi41      u0616(.An(men_men_n644_), .B(men_men_n378_), .C(men_men_n69_), .D(men_men_n121_), .Y(men_men_n645_));
  OR2        u0617(.A(men_men_n645_), .B(men_men_n643_), .Y(men_men_n646_));
  NOi32      u0618(.An(d), .Bn(a), .C(e), .Y(men_men_n647_));
  NA2        u0619(.A(men_men_n647_), .B(men_men_n117_), .Y(men_men_n648_));
  NO2        u0620(.A(n), .B(c), .Y(men_men_n649_));
  NA3        u0621(.A(men_men_n649_), .B(men_men_n29_), .C(m), .Y(men_men_n650_));
  NAi32      u0622(.An(n), .Bn(f), .C(m), .Y(men_men_n651_));
  NA3        u0623(.A(men_men_n651_), .B(men_men_n650_), .C(men_men_n648_), .Y(men_men_n652_));
  NOi32      u0624(.An(e), .Bn(a), .C(d), .Y(men_men_n653_));
  AOI210     u0625(.A0(men_men_n29_), .A1(d), .B0(men_men_n653_), .Y(men_men_n654_));
  AOI210     u0626(.A0(men_men_n654_), .A1(men_men_n225_), .B0(men_men_n591_), .Y(men_men_n655_));
  AOI210     u0627(.A0(men_men_n655_), .A1(men_men_n652_), .B0(men_men_n646_), .Y(men_men_n656_));
  OAI210     u0628(.A0(men_men_n263_), .A1(men_men_n89_), .B0(men_men_n656_), .Y(men_men_n657_));
  AOI210     u0629(.A0(men_men_n641_), .A1(men_men_n627_), .B0(men_men_n657_), .Y(men_men_n658_));
  NO3        u0630(.A(men_men_n338_), .B(men_men_n61_), .C(n), .Y(men_men_n659_));
  NA3        u0631(.A(men_men_n549_), .B(men_men_n181_), .C(men_men_n180_), .Y(men_men_n660_));
  NA2        u0632(.A(men_men_n493_), .B(men_men_n243_), .Y(men_men_n661_));
  OR2        u0633(.A(men_men_n661_), .B(men_men_n660_), .Y(men_men_n662_));
  NA2        u0634(.A(men_men_n76_), .B(men_men_n117_), .Y(men_men_n663_));
  NO2        u0635(.A(men_men_n663_), .B(men_men_n45_), .Y(men_men_n664_));
  AOI220     u0636(.A0(men_men_n664_), .A1(men_men_n579_), .B0(men_men_n662_), .B1(men_men_n659_), .Y(men_men_n665_));
  NO2        u0637(.A(men_men_n665_), .B(men_men_n89_), .Y(men_men_n666_));
  NA3        u0638(.A(men_men_n593_), .B(men_men_n364_), .C(men_men_n46_), .Y(men_men_n667_));
  NOi32      u0639(.An(e), .Bn(c), .C(f), .Y(men_men_n668_));
  NOi21      u0640(.An(f), .B(g), .Y(men_men_n669_));
  NO2        u0641(.A(men_men_n669_), .B(men_men_n223_), .Y(men_men_n670_));
  AOI220     u0642(.A0(men_men_n670_), .A1(men_men_n420_), .B0(men_men_n668_), .B1(men_men_n185_), .Y(men_men_n671_));
  NA3        u0643(.A(men_men_n671_), .B(men_men_n667_), .C(men_men_n188_), .Y(men_men_n672_));
  AOI210     u0644(.A0(men_men_n578_), .A1(men_men_n424_), .B0(men_men_n319_), .Y(men_men_n673_));
  NA2        u0645(.A(men_men_n673_), .B(men_men_n280_), .Y(men_men_n674_));
  NOi21      u0646(.An(j), .B(l), .Y(men_men_n675_));
  NAi21      u0647(.An(k), .B(h), .Y(men_men_n676_));
  NO2        u0648(.A(men_men_n676_), .B(men_men_n278_), .Y(men_men_n677_));
  NA2        u0649(.A(men_men_n677_), .B(men_men_n675_), .Y(men_men_n678_));
  OR2        u0650(.A(men_men_n678_), .B(men_men_n632_), .Y(men_men_n679_));
  NOi31      u0651(.An(m), .B(n), .C(k), .Y(men_men_n680_));
  NA2        u0652(.A(men_men_n675_), .B(men_men_n680_), .Y(men_men_n681_));
  AOI210     u0653(.A0(men_men_n424_), .A1(men_men_n398_), .B0(men_men_n319_), .Y(men_men_n682_));
  NAi21      u0654(.An(men_men_n681_), .B(men_men_n682_), .Y(men_men_n683_));
  NO2        u0655(.A(men_men_n294_), .B(men_men_n49_), .Y(men_men_n684_));
  NO2        u0656(.A(men_men_n331_), .B(men_men_n642_), .Y(men_men_n685_));
  NO2        u0657(.A(men_men_n574_), .B(men_men_n49_), .Y(men_men_n686_));
  AOI220     u0658(.A0(men_men_n686_), .A1(men_men_n685_), .B0(men_men_n684_), .B1(men_men_n613_), .Y(men_men_n687_));
  NA4        u0659(.A(men_men_n687_), .B(men_men_n683_), .C(men_men_n679_), .D(men_men_n674_), .Y(men_men_n688_));
  NA2        u0660(.A(men_men_n112_), .B(men_men_n36_), .Y(men_men_n689_));
  NO2        u0661(.A(k), .B(men_men_n226_), .Y(men_men_n690_));
  NO2        u0662(.A(men_men_n570_), .B(men_men_n387_), .Y(men_men_n691_));
  NAi31      u0663(.An(men_men_n689_), .B(men_men_n387_), .C(men_men_n690_), .Y(men_men_n692_));
  NO2        u0664(.A(men_men_n572_), .B(men_men_n186_), .Y(men_men_n693_));
  NA3        u0665(.A(men_men_n594_), .B(men_men_n287_), .C(men_men_n151_), .Y(men_men_n694_));
  NA2        u0666(.A(men_men_n545_), .B(men_men_n167_), .Y(men_men_n695_));
  NO2        u0667(.A(men_men_n421_), .B(men_men_n89_), .Y(men_men_n696_));
  AOI210     u0668(.A0(men_men_n694_), .A1(men_men_n693_), .B0(men_men_n696_), .Y(men_men_n697_));
  AN3        u0669(.A(f), .B(d), .C(b), .Y(men_men_n698_));
  OAI210     u0670(.A0(men_men_n698_), .A1(men_men_n135_), .B0(n), .Y(men_men_n699_));
  NA3        u0671(.A(men_men_n545_), .B(men_men_n167_), .C(men_men_n226_), .Y(men_men_n700_));
  AOI210     u0672(.A0(men_men_n699_), .A1(men_men_n245_), .B0(men_men_n700_), .Y(men_men_n701_));
  NAi31      u0673(.An(m), .B(n), .C(k), .Y(men_men_n702_));
  OR2        u0674(.A(men_men_n140_), .B(men_men_n61_), .Y(men_men_n703_));
  OAI210     u0675(.A0(men_men_n703_), .A1(men_men_n702_), .B0(men_men_n265_), .Y(men_men_n704_));
  OAI210     u0676(.A0(men_men_n704_), .A1(men_men_n701_), .B0(j), .Y(men_men_n705_));
  NA3        u0677(.A(men_men_n705_), .B(men_men_n697_), .C(men_men_n692_), .Y(men_men_n706_));
  NO4        u0678(.A(men_men_n706_), .B(men_men_n688_), .C(men_men_n672_), .D(men_men_n666_), .Y(men_men_n707_));
  NA2        u0679(.A(men_men_n408_), .B(men_men_n170_), .Y(men_men_n708_));
  NAi31      u0680(.An(g), .B(h), .C(f), .Y(men_men_n709_));
  OR3        u0681(.A(men_men_n709_), .B(men_men_n294_), .C(n), .Y(men_men_n710_));
  OA210      u0682(.A0(men_men_n574_), .A1(n), .B0(men_men_n630_), .Y(men_men_n711_));
  NA3        u0683(.A(men_men_n444_), .B(men_men_n125_), .C(men_men_n86_), .Y(men_men_n712_));
  OAI210     u0684(.A0(men_men_n711_), .A1(men_men_n93_), .B0(men_men_n712_), .Y(men_men_n713_));
  NOi21      u0685(.An(men_men_n710_), .B(men_men_n713_), .Y(men_men_n714_));
  AOI210     u0686(.A0(men_men_n714_), .A1(men_men_n708_), .B0(men_men_n567_), .Y(men_men_n715_));
  NO3        u0687(.A(g), .B(men_men_n225_), .C(men_men_n56_), .Y(men_men_n716_));
  NAi21      u0688(.An(h), .B(j), .Y(men_men_n717_));
  OAI210     u0689(.A0(men_men_n240_), .A1(men_men_n420_), .B0(men_men_n716_), .Y(men_men_n718_));
  OR2        u0690(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n719_));
  NA2        u0691(.A(men_men_n644_), .B(men_men_n366_), .Y(men_men_n720_));
  OA220      u0692(.A0(men_men_n681_), .A1(men_men_n720_), .B0(men_men_n678_), .B1(men_men_n719_), .Y(men_men_n721_));
  NA3        u0693(.A(men_men_n564_), .B(men_men_n102_), .C(men_men_n101_), .Y(men_men_n722_));
  AN2        u0694(.A(h), .B(f), .Y(men_men_n723_));
  NA2        u0695(.A(men_men_n723_), .B(men_men_n37_), .Y(men_men_n724_));
  NA2        u0696(.A(men_men_n102_), .B(men_men_n46_), .Y(men_men_n725_));
  OAI220     u0697(.A0(men_men_n725_), .A1(men_men_n355_), .B0(men_men_n724_), .B1(men_men_n498_), .Y(men_men_n726_));
  AOI210     u0698(.A0(men_men_n610_), .A1(men_men_n456_), .B0(men_men_n49_), .Y(men_men_n727_));
  OAI220     u0699(.A0(men_men_n633_), .A1(men_men_n626_), .B0(men_men_n348_), .B1(men_men_n565_), .Y(men_men_n728_));
  AOI210     u0700(.A0(men_men_n728_), .A1(men_men_n727_), .B0(men_men_n726_), .Y(men_men_n729_));
  NA4        u0701(.A(men_men_n729_), .B(men_men_n722_), .C(men_men_n721_), .D(men_men_n718_), .Y(men_men_n730_));
  NO2        u0702(.A(men_men_n267_), .B(f), .Y(men_men_n731_));
  NO2        u0703(.A(men_men_n669_), .B(men_men_n61_), .Y(men_men_n732_));
  NO3        u0704(.A(men_men_n732_), .B(men_men_n731_), .C(men_men_n34_), .Y(men_men_n733_));
  NA2        u0705(.A(men_men_n351_), .B(men_men_n146_), .Y(men_men_n734_));
  NA2        u0706(.A(men_men_n137_), .B(men_men_n49_), .Y(men_men_n735_));
  AOI220     u0707(.A0(men_men_n735_), .A1(men_men_n570_), .B0(men_men_n387_), .B1(men_men_n117_), .Y(men_men_n736_));
  OA220      u0708(.A0(men_men_n736_), .A1(men_men_n591_), .B0(men_men_n385_), .B1(men_men_n115_), .Y(men_men_n737_));
  OAI210     u0709(.A0(men_men_n734_), .A1(men_men_n733_), .B0(men_men_n737_), .Y(men_men_n738_));
  NO3        u0710(.A(men_men_n431_), .B(men_men_n203_), .C(men_men_n202_), .Y(men_men_n739_));
  NA2        u0711(.A(men_men_n739_), .B(men_men_n243_), .Y(men_men_n740_));
  NA3        u0712(.A(men_men_n740_), .B(men_men_n269_), .C(j), .Y(men_men_n741_));
  NO3        u0713(.A(men_men_n493_), .B(men_men_n183_), .C(i), .Y(men_men_n742_));
  NA2        u0714(.A(men_men_n497_), .B(men_men_n86_), .Y(men_men_n743_));
  NO4        u0715(.A(men_men_n567_), .B(men_men_n743_), .C(men_men_n136_), .D(men_men_n225_), .Y(men_men_n744_));
  AOI210     u0716(.A0(men_men_n742_), .A1(men_men_n176_), .B0(men_men_n744_), .Y(men_men_n745_));
  NA4        u0717(.A(men_men_n745_), .B(men_men_n741_), .C(men_men_n552_), .D(men_men_n429_), .Y(men_men_n746_));
  NO4        u0718(.A(men_men_n746_), .B(men_men_n738_), .C(men_men_n730_), .D(men_men_n715_), .Y(men_men_n747_));
  NA4        u0719(.A(men_men_n747_), .B(men_men_n707_), .C(men_men_n658_), .D(men_men_n624_), .Y(men08));
  NO2        u0720(.A(k), .B(h), .Y(men_men_n749_));
  AO210      u0721(.A0(men_men_n267_), .A1(men_men_n481_), .B0(men_men_n749_), .Y(men_men_n750_));
  NO2        u0722(.A(men_men_n750_), .B(men_men_n317_), .Y(men_men_n751_));
  NA2        u0723(.A(men_men_n668_), .B(men_men_n86_), .Y(men_men_n752_));
  NA2        u0724(.A(men_men_n752_), .B(men_men_n493_), .Y(men_men_n753_));
  AOI210     u0725(.A0(men_men_n753_), .A1(men_men_n751_), .B0(men_men_n528_), .Y(men_men_n754_));
  NO2        u0726(.A(a), .B(men_men_n57_), .Y(men_men_n755_));
  NO4        u0727(.A(men_men_n405_), .B(men_men_n116_), .C(j), .D(men_men_n226_), .Y(men_men_n756_));
  OAI210     u0728(.A0(men_men_n620_), .A1(men_men_n86_), .B0(men_men_n245_), .Y(men_men_n757_));
  AOI220     u0729(.A0(men_men_n757_), .A1(men_men_n372_), .B0(men_men_n756_), .B1(men_men_n755_), .Y(men_men_n758_));
  AOI210     u0730(.A0(men_men_n620_), .A1(men_men_n163_), .B0(men_men_n86_), .Y(men_men_n759_));
  NA4        u0731(.A(men_men_n228_), .B(men_men_n146_), .C(men_men_n45_), .D(h), .Y(men_men_n760_));
  AN2        u0732(.A(l), .B(k), .Y(men_men_n761_));
  NA4        u0733(.A(men_men_n761_), .B(men_men_n112_), .C(men_men_n75_), .D(men_men_n226_), .Y(men_men_n762_));
  OAI210     u0734(.A0(men_men_n760_), .A1(g), .B0(men_men_n762_), .Y(men_men_n763_));
  NA2        u0735(.A(men_men_n763_), .B(men_men_n759_), .Y(men_men_n764_));
  NA4        u0736(.A(men_men_n764_), .B(men_men_n758_), .C(men_men_n754_), .D(men_men_n374_), .Y(men_men_n765_));
  AN2        u0737(.A(men_men_n575_), .B(men_men_n98_), .Y(men_men_n766_));
  NO4        u0738(.A(men_men_n183_), .B(men_men_n419_), .C(men_men_n116_), .D(g), .Y(men_men_n767_));
  AOI210     u0739(.A0(men_men_n767_), .A1(men_men_n757_), .B0(men_men_n559_), .Y(men_men_n768_));
  NO2        u0740(.A(men_men_n38_), .B(men_men_n225_), .Y(men_men_n769_));
  AOI220     u0741(.A0(men_men_n670_), .A1(men_men_n371_), .B0(men_men_n769_), .B1(men_men_n607_), .Y(men_men_n770_));
  NAi31      u0742(.An(men_men_n766_), .B(men_men_n770_), .C(men_men_n768_), .Y(men_men_n771_));
  NO2        u0743(.A(men_men_n578_), .B(men_men_n35_), .Y(men_men_n772_));
  OAI210     u0744(.A0(men_men_n594_), .A1(men_men_n47_), .B0(men_men_n703_), .Y(men_men_n773_));
  AOI210     u0745(.A0(n), .A1(men_men_n773_), .B0(men_men_n772_), .Y(men_men_n774_));
  NO3        u0746(.A(men_men_n338_), .B(men_men_n136_), .C(men_men_n41_), .Y(men_men_n775_));
  NAi21      u0747(.An(men_men_n775_), .B(men_men_n762_), .Y(men_men_n776_));
  NA2        u0748(.A(men_men_n750_), .B(men_men_n141_), .Y(men_men_n777_));
  AOI220     u0749(.A0(men_men_n777_), .A1(men_men_n430_), .B0(men_men_n776_), .B1(men_men_n78_), .Y(men_men_n778_));
  OAI210     u0750(.A0(men_men_n774_), .A1(men_men_n89_), .B0(men_men_n778_), .Y(men_men_n779_));
  NA2        u0751(.A(men_men_n387_), .B(men_men_n43_), .Y(men_men_n780_));
  NA3        u0752(.A(men_men_n740_), .B(men_men_n357_), .C(men_men_n411_), .Y(men_men_n781_));
  NA2        u0753(.A(men_men_n761_), .B(men_men_n233_), .Y(men_men_n782_));
  NO2        u0754(.A(men_men_n782_), .B(men_men_n350_), .Y(men_men_n783_));
  AOI210     u0755(.A0(men_men_n783_), .A1(men_men_n731_), .B0(men_men_n527_), .Y(men_men_n784_));
  NA3        u0756(.A(m), .B(l), .C(k), .Y(men_men_n785_));
  AOI210     u0757(.A0(men_men_n712_), .A1(men_men_n710_), .B0(men_men_n785_), .Y(men_men_n786_));
  NO2        u0758(.A(men_men_n577_), .B(men_men_n288_), .Y(men_men_n787_));
  NOi21      u0759(.An(men_men_n787_), .B(men_men_n571_), .Y(men_men_n788_));
  NA4        u0760(.A(men_men_n117_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n789_));
  NA3        u0761(.A(men_men_n125_), .B(men_men_n439_), .C(i), .Y(men_men_n790_));
  NO2        u0762(.A(men_men_n790_), .B(men_men_n789_), .Y(men_men_n791_));
  NO3        u0763(.A(men_men_n791_), .B(men_men_n788_), .C(men_men_n786_), .Y(men_men_n792_));
  NA4        u0764(.A(men_men_n792_), .B(men_men_n784_), .C(men_men_n781_), .D(men_men_n780_), .Y(men_men_n793_));
  NO4        u0765(.A(men_men_n793_), .B(men_men_n779_), .C(men_men_n771_), .D(men_men_n765_), .Y(men_men_n794_));
  NA2        u0766(.A(men_men_n670_), .B(men_men_n420_), .Y(men_men_n795_));
  NOi31      u0767(.An(g), .B(h), .C(f), .Y(men_men_n796_));
  NA2        u0768(.A(men_men_n686_), .B(men_men_n796_), .Y(men_men_n797_));
  AO210      u0769(.A0(men_men_n797_), .A1(men_men_n634_), .B0(men_men_n580_), .Y(men_men_n798_));
  NO3        u0770(.A(men_men_n424_), .B(men_men_n565_), .C(h), .Y(men_men_n799_));
  AOI210     u0771(.A0(men_men_n799_), .A1(men_men_n117_), .B0(men_men_n538_), .Y(men_men_n800_));
  NA4        u0772(.A(men_men_n800_), .B(men_men_n798_), .C(men_men_n795_), .D(men_men_n266_), .Y(men_men_n801_));
  NA2        u0773(.A(men_men_n761_), .B(men_men_n75_), .Y(men_men_n802_));
  NO4        u0774(.A(men_men_n739_), .B(men_men_n183_), .C(n), .D(i), .Y(men_men_n803_));
  NOi21      u0775(.An(h), .B(j), .Y(men_men_n804_));
  NA2        u0776(.A(men_men_n804_), .B(f), .Y(men_men_n805_));
  NO2        u0777(.A(men_men_n805_), .B(men_men_n260_), .Y(men_men_n806_));
  NO3        u0778(.A(men_men_n806_), .B(men_men_n803_), .C(men_men_n742_), .Y(men_men_n807_));
  OAI220     u0779(.A0(men_men_n807_), .A1(men_men_n802_), .B0(men_men_n636_), .B1(men_men_n62_), .Y(men_men_n808_));
  AOI210     u0780(.A0(men_men_n801_), .A1(l), .B0(men_men_n808_), .Y(men_men_n809_));
  NO2        u0781(.A(j), .B(i), .Y(men_men_n810_));
  NA3        u0782(.A(men_men_n810_), .B(men_men_n82_), .C(l), .Y(men_men_n811_));
  NA2        u0783(.A(men_men_n810_), .B(men_men_n33_), .Y(men_men_n812_));
  NA2        u0784(.A(men_men_n449_), .B(men_men_n125_), .Y(men_men_n813_));
  OA220      u0785(.A0(men_men_n813_), .A1(men_men_n812_), .B0(men_men_n811_), .B1(men_men_n632_), .Y(men_men_n814_));
  NO3        u0786(.A(men_men_n158_), .B(men_men_n49_), .C(men_men_n114_), .Y(men_men_n815_));
  NO3        u0787(.A(c), .B(men_men_n156_), .C(men_men_n75_), .Y(men_men_n816_));
  NO3        u0788(.A(men_men_n520_), .B(men_men_n468_), .C(j), .Y(men_men_n817_));
  OAI210     u0789(.A0(men_men_n816_), .A1(men_men_n815_), .B0(men_men_n817_), .Y(men_men_n818_));
  OAI210     u0790(.A0(men_men_n797_), .A1(men_men_n62_), .B0(men_men_n818_), .Y(men_men_n819_));
  NA2        u0791(.A(k), .B(j), .Y(men_men_n820_));
  NO3        u0792(.A(men_men_n317_), .B(men_men_n820_), .C(men_men_n40_), .Y(men_men_n821_));
  AOI210     u0793(.A0(men_men_n570_), .A1(n), .B0(men_men_n593_), .Y(men_men_n822_));
  NA2        u0794(.A(men_men_n822_), .B(men_men_n596_), .Y(men_men_n823_));
  AN3        u0795(.A(men_men_n823_), .B(men_men_n821_), .C(men_men_n101_), .Y(men_men_n824_));
  NO3        u0796(.A(men_men_n183_), .B(men_men_n419_), .C(men_men_n116_), .Y(men_men_n825_));
  AOI220     u0797(.A0(men_men_n825_), .A1(men_men_n261_), .B0(men_men_n661_), .B1(men_men_n328_), .Y(men_men_n826_));
  NAi31      u0798(.An(men_men_n654_), .B(men_men_n95_), .C(men_men_n86_), .Y(men_men_n827_));
  NA2        u0799(.A(men_men_n827_), .B(men_men_n826_), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n317_), .B(men_men_n141_), .Y(men_men_n829_));
  AOI220     u0801(.A0(men_men_n829_), .A1(men_men_n670_), .B0(men_men_n775_), .B1(men_men_n759_), .Y(men_men_n830_));
  NO2        u0802(.A(men_men_n785_), .B(men_men_n93_), .Y(men_men_n831_));
  NA2        u0803(.A(men_men_n831_), .B(men_men_n631_), .Y(men_men_n832_));
  NO2        u0804(.A(men_men_n633_), .B(men_men_n121_), .Y(men_men_n833_));
  OAI210     u0805(.A0(men_men_n833_), .A1(men_men_n817_), .B0(men_men_n727_), .Y(men_men_n834_));
  NA3        u0806(.A(men_men_n834_), .B(men_men_n832_), .C(men_men_n830_), .Y(men_men_n835_));
  OR4        u0807(.A(men_men_n835_), .B(men_men_n828_), .C(men_men_n824_), .D(men_men_n819_), .Y(men_men_n836_));
  NA3        u0808(.A(men_men_n822_), .B(men_men_n596_), .C(men_men_n595_), .Y(men_men_n837_));
  NA4        u0809(.A(men_men_n837_), .B(men_men_n228_), .C(men_men_n481_), .D(men_men_n34_), .Y(men_men_n838_));
  NO4        u0810(.A(men_men_n520_), .B(men_men_n463_), .C(j), .D(f), .Y(men_men_n839_));
  OAI220     u0811(.A0(men_men_n760_), .A1(men_men_n752_), .B0(men_men_n355_), .B1(men_men_n38_), .Y(men_men_n840_));
  AOI210     u0812(.A0(men_men_n839_), .A1(men_men_n273_), .B0(men_men_n840_), .Y(men_men_n841_));
  NA3        u0813(.A(men_men_n586_), .B(men_men_n310_), .C(h), .Y(men_men_n842_));
  NOi21      u0814(.An(men_men_n727_), .B(men_men_n842_), .Y(men_men_n843_));
  NO2        u0815(.A(men_men_n94_), .B(men_men_n47_), .Y(men_men_n844_));
  OAI220     u0816(.A0(men_men_n842_), .A1(men_men_n650_), .B0(men_men_n811_), .B1(men_men_n719_), .Y(men_men_n845_));
  AOI210     u0817(.A0(men_men_n844_), .A1(men_men_n387_), .B0(men_men_n845_), .Y(men_men_n846_));
  NAi41      u0818(.An(men_men_n843_), .B(men_men_n846_), .C(men_men_n841_), .D(men_men_n838_), .Y(men_men_n847_));
  OR2        u0819(.A(men_men_n831_), .B(men_men_n98_), .Y(men_men_n848_));
  AOI220     u0820(.A0(men_men_n848_), .A1(men_men_n251_), .B0(men_men_n817_), .B1(men_men_n684_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n711_), .B(men_men_n75_), .Y(men_men_n850_));
  AOI210     u0822(.A0(men_men_n839_), .A1(men_men_n850_), .B0(men_men_n359_), .Y(men_men_n851_));
  OAI210     u0823(.A0(men_men_n785_), .A1(men_men_n709_), .B0(men_men_n558_), .Y(men_men_n852_));
  NA3        u0824(.A(men_men_n264_), .B(men_men_n59_), .C(b), .Y(men_men_n853_));
  AOI220     u0825(.A0(men_men_n649_), .A1(men_men_n29_), .B0(men_men_n497_), .B1(men_men_n86_), .Y(men_men_n854_));
  NA2        u0826(.A(men_men_n854_), .B(men_men_n853_), .Y(men_men_n855_));
  NO2        u0827(.A(men_men_n842_), .B(men_men_n526_), .Y(men_men_n856_));
  AOI210     u0828(.A0(men_men_n855_), .A1(men_men_n852_), .B0(men_men_n856_), .Y(men_men_n857_));
  NA3        u0829(.A(men_men_n857_), .B(men_men_n851_), .C(men_men_n849_), .Y(men_men_n858_));
  NOi41      u0830(.An(men_men_n814_), .B(men_men_n858_), .C(men_men_n847_), .D(men_men_n836_), .Y(men_men_n859_));
  OR3        u0831(.A(men_men_n760_), .B(men_men_n245_), .C(g), .Y(men_men_n860_));
  NO3        u0832(.A(men_men_n365_), .B(men_men_n319_), .C(men_men_n116_), .Y(men_men_n861_));
  NA2        u0833(.A(men_men_n861_), .B(men_men_n823_), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n863_));
  NO3        u0835(.A(men_men_n863_), .B(men_men_n812_), .C(men_men_n294_), .Y(men_men_n864_));
  NO3        u0836(.A(men_men_n565_), .B(men_men_n96_), .C(h), .Y(men_men_n865_));
  AOI210     u0837(.A0(men_men_n865_), .A1(men_men_n755_), .B0(men_men_n864_), .Y(men_men_n866_));
  NA4        u0838(.A(men_men_n866_), .B(men_men_n862_), .C(men_men_n860_), .D(men_men_n432_), .Y(men_men_n867_));
  OR2        u0839(.A(men_men_n709_), .B(men_men_n94_), .Y(men_men_n868_));
  NOi31      u0840(.An(b), .B(d), .C(a), .Y(men_men_n869_));
  NO2        u0841(.A(men_men_n869_), .B(men_men_n647_), .Y(men_men_n870_));
  NO2        u0842(.A(men_men_n870_), .B(n), .Y(men_men_n871_));
  NOi21      u0843(.An(men_men_n854_), .B(men_men_n871_), .Y(men_men_n872_));
  OAI220     u0844(.A0(men_men_n872_), .A1(men_men_n868_), .B0(men_men_n842_), .B1(men_men_n648_), .Y(men_men_n873_));
  NO2        u0845(.A(men_men_n594_), .B(men_men_n86_), .Y(men_men_n874_));
  NO3        u0846(.A(men_men_n669_), .B(men_men_n350_), .C(men_men_n121_), .Y(men_men_n875_));
  NOi21      u0847(.An(men_men_n875_), .B(men_men_n168_), .Y(men_men_n876_));
  AOI210     u0848(.A0(men_men_n861_), .A1(men_men_n874_), .B0(men_men_n876_), .Y(men_men_n877_));
  OAI210     u0849(.A0(men_men_n760_), .A1(men_men_n421_), .B0(men_men_n877_), .Y(men_men_n878_));
  NO2        u0850(.A(men_men_n739_), .B(n), .Y(men_men_n879_));
  AOI220     u0851(.A0(men_men_n829_), .A1(men_men_n716_), .B0(men_men_n879_), .B1(men_men_n751_), .Y(men_men_n880_));
  NO2        u0852(.A(men_men_n345_), .B(men_men_n250_), .Y(men_men_n881_));
  OAI210     u0853(.A0(men_men_n98_), .A1(men_men_n95_), .B0(men_men_n881_), .Y(men_men_n882_));
  NA2        u0854(.A(men_men_n125_), .B(men_men_n86_), .Y(men_men_n883_));
  AOI210     u0855(.A0(men_men_n453_), .A1(men_men_n445_), .B0(men_men_n883_), .Y(men_men_n884_));
  NAi21      u0856(.An(men_men_n884_), .B(men_men_n882_), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n783_), .B(men_men_n34_), .Y(men_men_n886_));
  NAi21      u0858(.An(men_men_n789_), .B(men_men_n464_), .Y(men_men_n887_));
  NO2        u0859(.A(men_men_n288_), .B(i), .Y(men_men_n888_));
  NA2        u0860(.A(men_men_n767_), .B(men_men_n373_), .Y(men_men_n889_));
  OAI210     u0861(.A0(men_men_n639_), .A1(men_men_n638_), .B0(men_men_n388_), .Y(men_men_n890_));
  AN3        u0862(.A(men_men_n890_), .B(men_men_n889_), .C(men_men_n887_), .Y(men_men_n891_));
  NAi41      u0863(.An(men_men_n885_), .B(men_men_n891_), .C(men_men_n886_), .D(men_men_n880_), .Y(men_men_n892_));
  NO4        u0864(.A(men_men_n892_), .B(men_men_n878_), .C(men_men_n873_), .D(men_men_n867_), .Y(men_men_n893_));
  NA4        u0865(.A(men_men_n893_), .B(men_men_n859_), .C(men_men_n809_), .D(men_men_n794_), .Y(men09));
  INV        u0866(.A(men_men_n126_), .Y(men_men_n895_));
  NA2        u0867(.A(f), .B(e), .Y(men_men_n896_));
  NO2        u0868(.A(men_men_n238_), .B(men_men_n116_), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n897_), .B(g), .Y(men_men_n898_));
  NA4        u0870(.A(men_men_n331_), .B(men_men_n506_), .C(men_men_n276_), .D(men_men_n123_), .Y(men_men_n899_));
  AOI210     u0871(.A0(men_men_n899_), .A1(g), .B0(men_men_n503_), .Y(men_men_n900_));
  AOI210     u0872(.A0(men_men_n900_), .A1(men_men_n898_), .B0(men_men_n896_), .Y(men_men_n901_));
  NO2        u0873(.A(men_men_n473_), .B(men_men_n549_), .Y(men_men_n902_));
  AOI210     u0874(.A0(men_men_n901_), .A1(men_men_n895_), .B0(men_men_n902_), .Y(men_men_n903_));
  NO2        u0875(.A(men_men_n215_), .B(men_men_n225_), .Y(men_men_n904_));
  NA3        u0876(.A(m), .B(l), .C(i), .Y(men_men_n905_));
  OAI220     u0877(.A0(men_men_n633_), .A1(men_men_n905_), .B0(men_men_n378_), .B1(men_men_n566_), .Y(men_men_n906_));
  NA4        u0878(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(f), .Y(men_men_n907_));
  NAi31      u0879(.An(men_men_n906_), .B(men_men_n907_), .C(men_men_n469_), .Y(men_men_n908_));
  OA210      u0880(.A0(men_men_n908_), .A1(men_men_n904_), .B0(men_men_n607_), .Y(men_men_n909_));
  NA3        u0881(.A(men_men_n868_), .B(men_men_n609_), .C(men_men_n558_), .Y(men_men_n910_));
  OA210      u0882(.A0(men_men_n910_), .A1(men_men_n909_), .B0(men_men_n871_), .Y(men_men_n911_));
  INV        u0883(.A(men_men_n362_), .Y(men_men_n912_));
  NO2        u0884(.A(men_men_n132_), .B(men_men_n130_), .Y(men_men_n913_));
  NOi31      u0885(.An(k), .B(m), .C(l), .Y(men_men_n914_));
  NO2        u0886(.A(men_men_n364_), .B(men_men_n914_), .Y(men_men_n915_));
  AOI210     u0887(.A0(men_men_n915_), .A1(men_men_n913_), .B0(men_men_n642_), .Y(men_men_n916_));
  NA2        u0888(.A(men_men_n853_), .B(men_men_n355_), .Y(men_men_n917_));
  NA2        u0889(.A(men_men_n366_), .B(men_men_n368_), .Y(men_men_n918_));
  OAI210     u0890(.A0(men_men_n215_), .A1(men_men_n225_), .B0(men_men_n918_), .Y(men_men_n919_));
  AOI220     u0891(.A0(men_men_n919_), .A1(men_men_n917_), .B0(men_men_n916_), .B1(men_men_n912_), .Y(men_men_n920_));
  NA2        u0892(.A(men_men_n177_), .B(men_men_n118_), .Y(men_men_n921_));
  NA3        u0893(.A(men_men_n921_), .B(men_men_n750_), .C(men_men_n141_), .Y(men_men_n922_));
  NA3        u0894(.A(men_men_n922_), .B(men_men_n200_), .C(men_men_n31_), .Y(men_men_n923_));
  NA4        u0895(.A(men_men_n923_), .B(men_men_n920_), .C(men_men_n671_), .D(men_men_n84_), .Y(men_men_n924_));
  NO2        u0896(.A(men_men_n629_), .B(men_men_n535_), .Y(men_men_n925_));
  NA2        u0897(.A(men_men_n925_), .B(men_men_n200_), .Y(men_men_n926_));
  NOi21      u0898(.An(f), .B(d), .Y(men_men_n927_));
  NA2        u0899(.A(men_men_n927_), .B(m), .Y(men_men_n928_));
  NO2        u0900(.A(men_men_n928_), .B(men_men_n52_), .Y(men_men_n929_));
  NOi32      u0901(.An(g), .Bn(f), .C(d), .Y(men_men_n930_));
  NA4        u0902(.A(men_men_n930_), .B(men_men_n649_), .C(men_men_n29_), .D(m), .Y(men_men_n931_));
  NOi21      u0903(.An(men_men_n332_), .B(men_men_n931_), .Y(men_men_n932_));
  AOI210     u0904(.A0(men_men_n929_), .A1(men_men_n584_), .B0(men_men_n932_), .Y(men_men_n933_));
  NA3        u0905(.A(men_men_n331_), .B(men_men_n276_), .C(men_men_n123_), .Y(men_men_n934_));
  AN2        u0906(.A(f), .B(d), .Y(men_men_n935_));
  NA3        u0907(.A(men_men_n511_), .B(men_men_n935_), .C(men_men_n86_), .Y(men_men_n936_));
  NO3        u0908(.A(men_men_n936_), .B(men_men_n75_), .C(men_men_n226_), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n303_), .B(men_men_n56_), .Y(men_men_n938_));
  OAI210     u0910(.A0(men_men_n938_), .A1(men_men_n934_), .B0(men_men_n937_), .Y(men_men_n939_));
  NAi41      u0911(.An(men_men_n525_), .B(men_men_n939_), .C(men_men_n933_), .D(men_men_n926_), .Y(men_men_n940_));
  NO4        u0912(.A(men_men_n669_), .B(men_men_n137_), .C(men_men_n350_), .D(men_men_n159_), .Y(men_men_n941_));
  NO2        u0913(.A(men_men_n702_), .B(men_men_n350_), .Y(men_men_n942_));
  AN2        u0914(.A(men_men_n942_), .B(men_men_n731_), .Y(men_men_n943_));
  NO3        u0915(.A(men_men_n943_), .B(men_men_n941_), .C(men_men_n247_), .Y(men_men_n944_));
  NA2        u0916(.A(men_men_n647_), .B(men_men_n86_), .Y(men_men_n945_));
  OAI220     u0917(.A0(men_men_n918_), .A1(men_men_n945_), .B0(men_men_n853_), .B1(men_men_n469_), .Y(men_men_n946_));
  NA3        u0918(.A(men_men_n167_), .B(men_men_n112_), .C(men_men_n111_), .Y(men_men_n947_));
  OAI220     u0919(.A0(men_men_n936_), .A1(men_men_n458_), .B0(men_men_n362_), .B1(men_men_n947_), .Y(men_men_n948_));
  NOi41      u0920(.An(men_men_n236_), .B(men_men_n948_), .C(men_men_n946_), .D(men_men_n326_), .Y(men_men_n949_));
  NA2        u0921(.A(c), .B(men_men_n120_), .Y(men_men_n950_));
  NO2        u0922(.A(men_men_n950_), .B(men_men_n436_), .Y(men_men_n951_));
  NA3        u0923(.A(men_men_n951_), .B(men_men_n547_), .C(f), .Y(men_men_n952_));
  OR2        u0924(.A(men_men_n709_), .B(men_men_n581_), .Y(men_men_n953_));
  OAI210     u0925(.A0(men_men_n612_), .A1(men_men_n663_), .B0(men_men_n953_), .Y(men_men_n954_));
  NA2        u0926(.A(men_men_n870_), .B(men_men_n115_), .Y(men_men_n955_));
  NA2        u0927(.A(men_men_n955_), .B(men_men_n954_), .Y(men_men_n956_));
  NA4        u0928(.A(men_men_n956_), .B(men_men_n952_), .C(men_men_n949_), .D(men_men_n944_), .Y(men_men_n957_));
  NO4        u0929(.A(men_men_n957_), .B(men_men_n940_), .C(men_men_n924_), .D(men_men_n911_), .Y(men_men_n958_));
  OR2        u0930(.A(men_men_n936_), .B(men_men_n75_), .Y(men_men_n959_));
  NA2        u0931(.A(men_men_n116_), .B(j), .Y(men_men_n960_));
  NO2        u0932(.A(men_men_n960_), .B(men_men_n150_), .Y(men_men_n961_));
  OAI210     u0933(.A0(men_men_n961_), .A1(men_men_n897_), .B0(g), .Y(men_men_n962_));
  AOI210     u0934(.A0(men_men_n962_), .A1(men_men_n311_), .B0(men_men_n959_), .Y(men_men_n963_));
  AOI210     u0935(.A0(men_men_n853_), .A1(men_men_n355_), .B0(men_men_n907_), .Y(men_men_n964_));
  NO2        u0936(.A(men_men_n141_), .B(men_men_n137_), .Y(men_men_n965_));
  NO2        u0937(.A(men_men_n243_), .B(men_men_n237_), .Y(men_men_n966_));
  AOI220     u0938(.A0(men_men_n966_), .A1(men_men_n240_), .B0(men_men_n324_), .B1(men_men_n965_), .Y(men_men_n967_));
  NO2        u0939(.A(men_men_n458_), .B(men_men_n896_), .Y(men_men_n968_));
  NA2        u0940(.A(men_men_n968_), .B(men_men_n601_), .Y(men_men_n969_));
  NA2        u0941(.A(men_men_n969_), .B(men_men_n967_), .Y(men_men_n970_));
  NA2        u0942(.A(e), .B(d), .Y(men_men_n971_));
  OAI220     u0943(.A0(men_men_n971_), .A1(c), .B0(men_men_n345_), .B1(d), .Y(men_men_n972_));
  NA3        u0944(.A(men_men_n972_), .B(men_men_n486_), .C(men_men_n545_), .Y(men_men_n973_));
  AOI210     u0945(.A0(men_men_n553_), .A1(men_men_n190_), .B0(men_men_n243_), .Y(men_men_n974_));
  AOI210     u0946(.A0(men_men_n670_), .A1(men_men_n371_), .B0(men_men_n974_), .Y(men_men_n975_));
  NA2        u0947(.A(men_men_n303_), .B(men_men_n173_), .Y(men_men_n976_));
  NA3        u0948(.A(men_men_n937_), .B(men_men_n976_), .C(men_men_n56_), .Y(men_men_n977_));
  NA3        u0949(.A(men_men_n176_), .B(men_men_n87_), .C(men_men_n34_), .Y(men_men_n978_));
  NA4        u0950(.A(men_men_n978_), .B(men_men_n977_), .C(men_men_n975_), .D(men_men_n973_), .Y(men_men_n979_));
  NO4        u0951(.A(men_men_n979_), .B(men_men_n970_), .C(men_men_n964_), .D(men_men_n963_), .Y(men_men_n980_));
  NA2        u0952(.A(men_men_n912_), .B(men_men_n31_), .Y(men_men_n981_));
  AO210      u0953(.A0(men_men_n981_), .A1(men_men_n752_), .B0(men_men_n229_), .Y(men_men_n982_));
  OAI220     u0954(.A0(men_men_n669_), .A1(men_men_n61_), .B0(men_men_n319_), .B1(j), .Y(men_men_n983_));
  AOI220     u0955(.A0(men_men_n983_), .A1(men_men_n942_), .B0(men_men_n659_), .B1(men_men_n668_), .Y(men_men_n984_));
  OAI210     u0956(.A0(men_men_n473_), .A1(men_men_n180_), .B0(men_men_n984_), .Y(men_men_n985_));
  OAI210     u0957(.A0(men_men_n897_), .A1(men_men_n976_), .B0(men_men_n930_), .Y(men_men_n986_));
  NO2        u0958(.A(men_men_n986_), .B(men_men_n650_), .Y(men_men_n987_));
  AOI210     u0959(.A0(men_men_n122_), .A1(men_men_n121_), .B0(men_men_n275_), .Y(men_men_n988_));
  NO2        u0960(.A(men_men_n988_), .B(men_men_n931_), .Y(men_men_n989_));
  AO210      u0961(.A0(men_men_n917_), .A1(men_men_n906_), .B0(men_men_n989_), .Y(men_men_n990_));
  NOi31      u0962(.An(men_men_n584_), .B(men_men_n928_), .C(men_men_n311_), .Y(men_men_n991_));
  NO4        u0963(.A(men_men_n991_), .B(men_men_n990_), .C(men_men_n987_), .D(men_men_n985_), .Y(men_men_n992_));
  AO220      u0964(.A0(men_men_n486_), .A1(men_men_n804_), .B0(men_men_n185_), .B1(f), .Y(men_men_n993_));
  OAI210     u0965(.A0(men_men_n993_), .A1(men_men_n489_), .B0(men_men_n972_), .Y(men_men_n994_));
  NO2        u0966(.A(men_men_n468_), .B(men_men_n71_), .Y(men_men_n995_));
  OAI210     u0967(.A0(men_men_n910_), .A1(men_men_n995_), .B0(men_men_n755_), .Y(men_men_n996_));
  AN4        u0968(.A(men_men_n996_), .B(men_men_n994_), .C(men_men_n992_), .D(men_men_n982_), .Y(men_men_n997_));
  NA4        u0969(.A(men_men_n997_), .B(men_men_n980_), .C(men_men_n958_), .D(men_men_n903_), .Y(men12));
  NO2        u0970(.A(men_men_n484_), .B(c), .Y(men_men_n999_));
  NO4        u0971(.A(men_men_n473_), .B(men_men_n267_), .C(men_men_n625_), .D(men_men_n226_), .Y(men_men_n1000_));
  NA2        u0972(.A(men_men_n1000_), .B(men_men_n999_), .Y(men_men_n1001_));
  NA2        u0973(.A(men_men_n584_), .B(men_men_n995_), .Y(men_men_n1002_));
  NO3        u0974(.A(men_men_n484_), .B(men_men_n86_), .C(men_men_n120_), .Y(men_men_n1003_));
  NO2        u0975(.A(men_men_n913_), .B(men_men_n378_), .Y(men_men_n1004_));
  NO2        u0976(.A(men_men_n709_), .B(men_men_n405_), .Y(men_men_n1005_));
  AOI220     u0977(.A0(men_men_n1005_), .A1(men_men_n583_), .B0(men_men_n1004_), .B1(men_men_n1003_), .Y(men_men_n1006_));
  NA4        u0978(.A(men_men_n1006_), .B(men_men_n1002_), .C(men_men_n1001_), .D(men_men_n472_), .Y(men_men_n1007_));
  AOI210     u0979(.A0(men_men_n246_), .A1(men_men_n361_), .B0(men_men_n212_), .Y(men_men_n1008_));
  OR2        u0980(.A(men_men_n1008_), .B(men_men_n1000_), .Y(men_men_n1009_));
  OAI210     u0981(.A0(men_men_n416_), .A1(men_men_n1009_), .B0(men_men_n431_), .Y(men_men_n1010_));
  NO2        u0982(.A(men_men_n689_), .B(men_men_n278_), .Y(men_men_n1011_));
  NO2        u0983(.A(men_men_n633_), .B(men_men_n905_), .Y(men_men_n1012_));
  AOI220     u0984(.A0(men_men_n1012_), .A1(men_men_n607_), .B0(men_men_n881_), .B1(men_men_n1011_), .Y(men_men_n1013_));
  NO2        u0985(.A(men_men_n158_), .B(men_men_n250_), .Y(men_men_n1014_));
  NA3        u0986(.A(men_men_n1014_), .B(men_men_n253_), .C(i), .Y(men_men_n1015_));
  NA3        u0987(.A(men_men_n1015_), .B(men_men_n1013_), .C(men_men_n1010_), .Y(men_men_n1016_));
  OR2        u0988(.A(men_men_n346_), .B(men_men_n1003_), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n1017_), .B(men_men_n379_), .Y(men_men_n1018_));
  NO3        u0990(.A(men_men_n137_), .B(men_men_n159_), .C(men_men_n226_), .Y(men_men_n1019_));
  NA2        u0991(.A(men_men_n1019_), .B(men_men_n570_), .Y(men_men_n1020_));
  NA4        u0992(.A(men_men_n474_), .B(men_men_n466_), .C(men_men_n191_), .D(g), .Y(men_men_n1021_));
  NA3        u0993(.A(men_men_n1021_), .B(men_men_n1020_), .C(men_men_n1018_), .Y(men_men_n1022_));
  NO3        u0994(.A(men_men_n714_), .B(men_men_n94_), .C(men_men_n45_), .Y(men_men_n1023_));
  NO4        u0995(.A(men_men_n1023_), .B(men_men_n1022_), .C(men_men_n1016_), .D(men_men_n1007_), .Y(men_men_n1024_));
  NO2        u0996(.A(men_men_n395_), .B(men_men_n394_), .Y(men_men_n1025_));
  NA2        u0997(.A(men_men_n630_), .B(men_men_n73_), .Y(men_men_n1026_));
  NA2        u0998(.A(men_men_n594_), .B(men_men_n151_), .Y(men_men_n1027_));
  NOi21      u0999(.An(men_men_n34_), .B(men_men_n702_), .Y(men_men_n1028_));
  AOI220     u1000(.A0(men_men_n1028_), .A1(men_men_n1027_), .B0(men_men_n1026_), .B1(men_men_n1025_), .Y(men_men_n1029_));
  OAI210     u1001(.A0(men_men_n265_), .A1(men_men_n45_), .B0(men_men_n1029_), .Y(men_men_n1030_));
  NA2        u1002(.A(men_men_n464_), .B(men_men_n280_), .Y(men_men_n1031_));
  NO3        u1003(.A(men_men_n883_), .B(men_men_n91_), .C(men_men_n436_), .Y(men_men_n1032_));
  NAi31      u1004(.An(men_men_n1032_), .B(men_men_n1031_), .C(men_men_n342_), .Y(men_men_n1033_));
  NO2        u1005(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n1034_));
  NO2        u1006(.A(men_men_n541_), .B(men_men_n319_), .Y(men_men_n1035_));
  NO2        u1007(.A(men_men_n541_), .B(men_men_n151_), .Y(men_men_n1036_));
  NA2        u1008(.A(men_men_n680_), .B(men_men_n388_), .Y(men_men_n1037_));
  OAI210     u1009(.A0(men_men_n790_), .A1(men_men_n1037_), .B0(men_men_n392_), .Y(men_men_n1038_));
  NO4        u1010(.A(men_men_n1038_), .B(men_men_n1036_), .C(men_men_n1033_), .D(men_men_n1030_), .Y(men_men_n1039_));
  NA2        u1011(.A(men_men_n371_), .B(g), .Y(men_men_n1040_));
  NA2        u1012(.A(men_men_n170_), .B(i), .Y(men_men_n1041_));
  NA2        u1013(.A(men_men_n46_), .B(i), .Y(men_men_n1042_));
  OAI220     u1014(.A0(men_men_n1042_), .A1(men_men_n211_), .B0(men_men_n1041_), .B1(men_men_n94_), .Y(men_men_n1043_));
  AOI210     u1015(.A0(men_men_n447_), .A1(men_men_n37_), .B0(men_men_n1043_), .Y(men_men_n1044_));
  NO2        u1016(.A(men_men_n151_), .B(men_men_n86_), .Y(men_men_n1045_));
  OR2        u1017(.A(men_men_n1045_), .B(men_men_n593_), .Y(men_men_n1046_));
  NA2        u1018(.A(men_men_n594_), .B(men_men_n409_), .Y(men_men_n1047_));
  AOI210     u1019(.A0(men_men_n1047_), .A1(n), .B0(men_men_n1046_), .Y(men_men_n1048_));
  OAI220     u1020(.A0(men_men_n1048_), .A1(men_men_n1040_), .B0(men_men_n1044_), .B1(men_men_n355_), .Y(men_men_n1049_));
  NO2        u1021(.A(men_men_n709_), .B(men_men_n535_), .Y(men_men_n1050_));
  NA3        u1022(.A(men_men_n366_), .B(men_men_n675_), .C(i), .Y(men_men_n1051_));
  OAI210     u1023(.A0(men_men_n468_), .A1(men_men_n331_), .B0(men_men_n1051_), .Y(men_men_n1052_));
  OAI220     u1024(.A0(men_men_n1052_), .A1(men_men_n1050_), .B0(men_men_n727_), .B1(men_men_n816_), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n653_), .B(men_men_n117_), .Y(men_men_n1054_));
  OR3        u1026(.A(men_men_n331_), .B(men_men_n463_), .C(f), .Y(men_men_n1055_));
  NA3        u1027(.A(men_men_n675_), .B(men_men_n82_), .C(i), .Y(men_men_n1056_));
  OA220      u1028(.A0(men_men_n1056_), .A1(men_men_n1054_), .B0(men_men_n1055_), .B1(men_men_n632_), .Y(men_men_n1057_));
  NA3        u1029(.A(men_men_n347_), .B(men_men_n122_), .C(g), .Y(men_men_n1058_));
  AOI210     u1030(.A0(men_men_n724_), .A1(men_men_n1058_), .B0(m), .Y(men_men_n1059_));
  OAI210     u1031(.A0(men_men_n1059_), .A1(men_men_n1004_), .B0(men_men_n346_), .Y(men_men_n1060_));
  NA2        u1032(.A(men_men_n743_), .B(men_men_n945_), .Y(men_men_n1061_));
  NA2        u1033(.A(men_men_n907_), .B(men_men_n469_), .Y(men_men_n1062_));
  NA2        u1034(.A(men_men_n234_), .B(men_men_n79_), .Y(men_men_n1063_));
  NA3        u1035(.A(men_men_n1063_), .B(men_men_n1056_), .C(men_men_n1055_), .Y(men_men_n1064_));
  AOI220     u1036(.A0(men_men_n1064_), .A1(men_men_n273_), .B0(men_men_n1062_), .B1(men_men_n1061_), .Y(men_men_n1065_));
  NA4        u1037(.A(men_men_n1065_), .B(men_men_n1060_), .C(men_men_n1057_), .D(men_men_n1053_), .Y(men_men_n1066_));
  NO2        u1038(.A(men_men_n405_), .B(men_men_n93_), .Y(men_men_n1067_));
  OAI210     u1039(.A0(men_men_n1067_), .A1(men_men_n1011_), .B0(men_men_n251_), .Y(men_men_n1068_));
  NA2        u1040(.A(men_men_n713_), .B(men_men_n90_), .Y(men_men_n1069_));
  NO2        u1041(.A(men_men_n492_), .B(men_men_n226_), .Y(men_men_n1070_));
  AOI220     u1042(.A0(men_men_n1070_), .A1(men_men_n410_), .B0(men_men_n1017_), .B1(men_men_n230_), .Y(men_men_n1071_));
  AOI220     u1043(.A0(men_men_n1005_), .A1(men_men_n1014_), .B0(men_men_n631_), .B1(men_men_n92_), .Y(men_men_n1072_));
  NA4        u1044(.A(men_men_n1072_), .B(men_men_n1071_), .C(men_men_n1069_), .D(men_men_n1068_), .Y(men_men_n1073_));
  OAI210     u1045(.A0(men_men_n1062_), .A1(men_men_n1012_), .B0(men_men_n583_), .Y(men_men_n1074_));
  AOI210     u1046(.A0(men_men_n448_), .A1(men_men_n440_), .B0(men_men_n883_), .Y(men_men_n1075_));
  OAI210     u1047(.A0(men_men_n395_), .A1(men_men_n394_), .B0(men_men_n113_), .Y(men_men_n1076_));
  AOI210     u1048(.A0(men_men_n1076_), .A1(men_men_n575_), .B0(men_men_n1075_), .Y(men_men_n1077_));
  NA2        u1049(.A(men_men_n1059_), .B(men_men_n1003_), .Y(men_men_n1078_));
  NO3        u1050(.A(men_men_n960_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1079_));
  AOI220     u1051(.A0(men_men_n1079_), .A1(men_men_n673_), .B0(men_men_n693_), .B1(men_men_n570_), .Y(men_men_n1080_));
  NA4        u1052(.A(men_men_n1080_), .B(men_men_n1078_), .C(men_men_n1077_), .D(men_men_n1074_), .Y(men_men_n1081_));
  NO4        u1053(.A(men_men_n1081_), .B(men_men_n1073_), .C(men_men_n1066_), .D(men_men_n1049_), .Y(men_men_n1082_));
  NAi31      u1054(.An(men_men_n147_), .B(men_men_n449_), .C(n), .Y(men_men_n1083_));
  NO3        u1055(.A(men_men_n130_), .B(men_men_n364_), .C(men_men_n914_), .Y(men_men_n1084_));
  NO2        u1056(.A(men_men_n1084_), .B(men_men_n1083_), .Y(men_men_n1085_));
  NO3        u1057(.A(men_men_n288_), .B(men_men_n147_), .C(men_men_n436_), .Y(men_men_n1086_));
  AOI210     u1058(.A0(men_men_n1086_), .A1(n), .B0(men_men_n1085_), .Y(men_men_n1087_));
  NA2        u1059(.A(men_men_n528_), .B(i), .Y(men_men_n1088_));
  NA2        u1060(.A(men_men_n1088_), .B(men_men_n1087_), .Y(men_men_n1089_));
  NA2        u1061(.A(men_men_n243_), .B(men_men_n181_), .Y(men_men_n1090_));
  NO3        u1062(.A(men_men_n328_), .B(men_men_n474_), .C(men_men_n185_), .Y(men_men_n1091_));
  NOi31      u1063(.An(men_men_n1090_), .B(men_men_n1091_), .C(men_men_n226_), .Y(men_men_n1092_));
  NAi21      u1064(.An(men_men_n594_), .B(men_men_n1070_), .Y(men_men_n1093_));
  NA2        u1065(.A(men_men_n467_), .B(men_men_n945_), .Y(men_men_n1094_));
  NO3        u1066(.A(men_men_n468_), .B(men_men_n331_), .C(men_men_n75_), .Y(men_men_n1095_));
  AOI220     u1067(.A0(men_men_n1095_), .A1(men_men_n1094_), .B0(men_men_n517_), .B1(g), .Y(men_men_n1096_));
  NA2        u1068(.A(men_men_n1096_), .B(men_men_n1093_), .Y(men_men_n1097_));
  OAI220     u1069(.A0(men_men_n1083_), .A1(men_men_n246_), .B0(men_men_n1051_), .B1(men_men_n648_), .Y(men_men_n1098_));
  NO2        u1070(.A(men_men_n710_), .B(men_men_n405_), .Y(men_men_n1099_));
  NA2        u1071(.A(men_men_n1008_), .B(men_men_n999_), .Y(men_men_n1100_));
  NO3        u1072(.A(c), .B(men_men_n156_), .C(men_men_n225_), .Y(men_men_n1101_));
  OAI210     u1073(.A0(men_men_n1101_), .A1(men_men_n564_), .B0(men_men_n406_), .Y(men_men_n1102_));
  OAI220     u1074(.A0(men_men_n1005_), .A1(men_men_n1012_), .B0(men_men_n584_), .B1(men_men_n457_), .Y(men_men_n1103_));
  NA4        u1075(.A(men_men_n1103_), .B(men_men_n1102_), .C(men_men_n1100_), .D(men_men_n667_), .Y(men_men_n1104_));
  OAI210     u1076(.A0(men_men_n1008_), .A1(men_men_n1000_), .B0(men_men_n1090_), .Y(men_men_n1105_));
  NA3        u1077(.A(men_men_n1047_), .B(men_men_n522_), .C(men_men_n46_), .Y(men_men_n1106_));
  AOI210     u1078(.A0(men_men_n408_), .A1(men_men_n406_), .B0(men_men_n354_), .Y(men_men_n1107_));
  NA4        u1079(.A(men_men_n1107_), .B(men_men_n1106_), .C(men_men_n1105_), .D(men_men_n289_), .Y(men_men_n1108_));
  OR4        u1080(.A(men_men_n1108_), .B(men_men_n1104_), .C(men_men_n1099_), .D(men_men_n1098_), .Y(men_men_n1109_));
  NO4        u1081(.A(men_men_n1109_), .B(men_men_n1097_), .C(men_men_n1092_), .D(men_men_n1089_), .Y(men_men_n1110_));
  NA4        u1082(.A(men_men_n1110_), .B(men_men_n1082_), .C(men_men_n1039_), .D(men_men_n1024_), .Y(men13));
  NA2        u1083(.A(men_men_n46_), .B(men_men_n89_), .Y(men_men_n1112_));
  AN2        u1084(.A(c), .B(b), .Y(men_men_n1113_));
  NA3        u1085(.A(men_men_n264_), .B(men_men_n1113_), .C(m), .Y(men_men_n1114_));
  NO4        u1086(.A(e), .B(men_men_n1114_), .C(men_men_n1112_), .D(men_men_n626_), .Y(men_men_n1115_));
  NA2        u1087(.A(men_men_n280_), .B(men_men_n1113_), .Y(men_men_n1116_));
  NO4        u1088(.A(men_men_n1116_), .B(e), .C(men_men_n1041_), .D(a), .Y(men_men_n1117_));
  NAi32      u1089(.An(d), .Bn(c), .C(e), .Y(men_men_n1118_));
  NA2        u1090(.A(men_men_n146_), .B(men_men_n45_), .Y(men_men_n1119_));
  NO4        u1091(.A(men_men_n1119_), .B(men_men_n1118_), .C(men_men_n633_), .D(men_men_n327_), .Y(men_men_n1120_));
  NA2        u1092(.A(men_men_n717_), .B(men_men_n237_), .Y(men_men_n1121_));
  NA2        u1093(.A(men_men_n439_), .B(men_men_n225_), .Y(men_men_n1122_));
  AN2        u1094(.A(d), .B(c), .Y(men_men_n1123_));
  NA2        u1095(.A(men_men_n1123_), .B(men_men_n120_), .Y(men_men_n1124_));
  NO4        u1096(.A(men_men_n1124_), .B(men_men_n1122_), .C(men_men_n186_), .D(men_men_n177_), .Y(men_men_n1125_));
  NA2        u1097(.A(men_men_n533_), .B(c), .Y(men_men_n1126_));
  NO4        u1098(.A(men_men_n1119_), .B(men_men_n629_), .C(men_men_n1126_), .D(men_men_n327_), .Y(men_men_n1127_));
  AO210      u1099(.A0(men_men_n1125_), .A1(men_men_n1121_), .B0(men_men_n1127_), .Y(men_men_n1128_));
  OR4        u1100(.A(men_men_n1128_), .B(men_men_n1120_), .C(men_men_n1117_), .D(men_men_n1115_), .Y(men_men_n1129_));
  NAi32      u1101(.An(f), .Bn(e), .C(c), .Y(men_men_n1130_));
  NO2        u1102(.A(men_men_n1130_), .B(men_men_n153_), .Y(men_men_n1131_));
  NA2        u1103(.A(men_men_n1131_), .B(g), .Y(men_men_n1132_));
  OR3        u1104(.A(men_men_n237_), .B(men_men_n186_), .C(men_men_n177_), .Y(men_men_n1133_));
  NO2        u1105(.A(men_men_n1133_), .B(men_men_n1132_), .Y(men_men_n1134_));
  NO2        u1106(.A(men_men_n1126_), .B(men_men_n327_), .Y(men_men_n1135_));
  NO2        u1107(.A(j), .B(men_men_n45_), .Y(men_men_n1136_));
  NA2        u1108(.A(men_men_n677_), .B(men_men_n1136_), .Y(men_men_n1137_));
  NOi21      u1109(.An(men_men_n1135_), .B(men_men_n1137_), .Y(men_men_n1138_));
  NO2        u1110(.A(men_men_n820_), .B(men_men_n116_), .Y(men_men_n1139_));
  NOi41      u1111(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1140_));
  NA2        u1112(.A(men_men_n1140_), .B(men_men_n1139_), .Y(men_men_n1141_));
  NO2        u1113(.A(men_men_n1141_), .B(men_men_n1132_), .Y(men_men_n1142_));
  OR3        u1114(.A(e), .B(d), .C(c), .Y(men_men_n1143_));
  NA3        u1115(.A(k), .B(j), .C(i), .Y(men_men_n1144_));
  NO3        u1116(.A(men_men_n1144_), .B(men_men_n327_), .C(men_men_n93_), .Y(men_men_n1145_));
  NOi21      u1117(.An(men_men_n1145_), .B(men_men_n1143_), .Y(men_men_n1146_));
  OR4        u1118(.A(men_men_n1146_), .B(men_men_n1142_), .C(men_men_n1138_), .D(men_men_n1134_), .Y(men_men_n1147_));
  NA3        u1119(.A(men_men_n500_), .B(men_men_n357_), .C(men_men_n56_), .Y(men_men_n1148_));
  NO2        u1120(.A(men_men_n1148_), .B(men_men_n1137_), .Y(men_men_n1149_));
  NO4        u1121(.A(men_men_n1148_), .B(men_men_n629_), .C(men_men_n481_), .D(men_men_n45_), .Y(men_men_n1150_));
  NO2        u1122(.A(f), .B(c), .Y(men_men_n1151_));
  NOi21      u1123(.An(men_men_n1151_), .B(men_men_n473_), .Y(men_men_n1152_));
  NA2        u1124(.A(men_men_n1152_), .B(men_men_n59_), .Y(men_men_n1153_));
  OR2        u1125(.A(k), .B(i), .Y(men_men_n1154_));
  NO3        u1126(.A(men_men_n1154_), .B(men_men_n257_), .C(l), .Y(men_men_n1155_));
  NOi31      u1127(.An(men_men_n1155_), .B(men_men_n1153_), .C(j), .Y(men_men_n1156_));
  OR3        u1128(.A(men_men_n1156_), .B(men_men_n1150_), .C(men_men_n1149_), .Y(men_men_n1157_));
  OR3        u1129(.A(men_men_n1157_), .B(men_men_n1147_), .C(men_men_n1129_), .Y(men02));
  OR2        u1130(.A(l), .B(k), .Y(men_men_n1159_));
  OR3        u1131(.A(h), .B(g), .C(f), .Y(men_men_n1160_));
  OR3        u1132(.A(n), .B(m), .C(i), .Y(men_men_n1161_));
  NO4        u1133(.A(men_men_n1161_), .B(men_men_n1160_), .C(men_men_n1159_), .D(men_men_n1143_), .Y(men_men_n1162_));
  NOi31      u1134(.An(e), .B(d), .C(c), .Y(men_men_n1163_));
  AOI210     u1135(.A0(men_men_n1145_), .A1(men_men_n1163_), .B0(men_men_n1120_), .Y(men_men_n1164_));
  AN3        u1136(.A(g), .B(f), .C(c), .Y(men_men_n1165_));
  NA3        u1137(.A(men_men_n1165_), .B(men_men_n500_), .C(h), .Y(men_men_n1166_));
  OR2        u1138(.A(men_men_n1144_), .B(men_men_n327_), .Y(men_men_n1167_));
  OR2        u1139(.A(men_men_n1167_), .B(men_men_n1166_), .Y(men_men_n1168_));
  NO3        u1140(.A(men_men_n1148_), .B(men_men_n1119_), .C(men_men_n629_), .Y(men_men_n1169_));
  NO2        u1141(.A(men_men_n1169_), .B(men_men_n1134_), .Y(men_men_n1170_));
  NA3        u1142(.A(l), .B(k), .C(j), .Y(men_men_n1171_));
  NA2        u1143(.A(i), .B(h), .Y(men_men_n1172_));
  NO3        u1144(.A(men_men_n1172_), .B(men_men_n1171_), .C(men_men_n137_), .Y(men_men_n1173_));
  NO3        u1145(.A(men_men_n148_), .B(men_men_n301_), .C(men_men_n226_), .Y(men_men_n1174_));
  AOI210     u1146(.A0(men_men_n1174_), .A1(men_men_n1173_), .B0(men_men_n1138_), .Y(men_men_n1175_));
  NA3        u1147(.A(c), .B(b), .C(a), .Y(men_men_n1176_));
  NO3        u1148(.A(men_men_n1176_), .B(men_men_n971_), .C(men_men_n225_), .Y(men_men_n1177_));
  NO4        u1149(.A(men_men_n1144_), .B(men_men_n319_), .C(men_men_n49_), .D(men_men_n116_), .Y(men_men_n1178_));
  AOI210     u1150(.A0(men_men_n1178_), .A1(men_men_n1177_), .B0(men_men_n1149_), .Y(men_men_n1179_));
  AN4        u1151(.A(men_men_n1179_), .B(men_men_n1175_), .C(men_men_n1170_), .D(men_men_n1168_), .Y(men_men_n1180_));
  NA2        u1152(.A(men_men_n1141_), .B(men_men_n1133_), .Y(men_men_n1181_));
  AOI210     u1153(.A0(men_men_n1181_), .A1(men_men_n225_), .B0(men_men_n1115_), .Y(men_men_n1182_));
  NAi41      u1154(.An(men_men_n1162_), .B(men_men_n1182_), .C(men_men_n1180_), .D(men_men_n1164_), .Y(men03));
  NO2        u1155(.A(men_men_n566_), .B(men_men_n642_), .Y(men_men_n1184_));
  NA4        u1156(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(men_men_n225_), .Y(men_men_n1185_));
  NA4        u1157(.A(men_men_n617_), .B(m), .C(men_men_n116_), .D(men_men_n225_), .Y(men_men_n1186_));
  NA3        u1158(.A(men_men_n1186_), .B(men_men_n396_), .C(men_men_n1185_), .Y(men_men_n1187_));
  NO3        u1159(.A(men_men_n1187_), .B(men_men_n1184_), .C(men_men_n1076_), .Y(men_men_n1188_));
  NOi41      u1160(.An(men_men_n868_), .B(men_men_n919_), .C(men_men_n908_), .D(men_men_n769_), .Y(men_men_n1189_));
  OAI220     u1161(.A0(men_men_n1189_), .A1(men_men_n743_), .B0(men_men_n1188_), .B1(men_men_n630_), .Y(men_men_n1190_));
  NOi31      u1162(.An(i), .B(k), .C(j), .Y(men_men_n1191_));
  NA4        u1163(.A(men_men_n1191_), .B(men_men_n1163_), .C(men_men_n366_), .D(men_men_n357_), .Y(men_men_n1192_));
  OAI210     u1164(.A0(men_men_n883_), .A1(men_men_n450_), .B0(men_men_n1192_), .Y(men_men_n1193_));
  NOi31      u1165(.An(m), .B(n), .C(f), .Y(men_men_n1194_));
  NA2        u1166(.A(men_men_n1194_), .B(men_men_n51_), .Y(men_men_n1195_));
  AN2        u1167(.A(e), .B(c), .Y(men_men_n1196_));
  NA2        u1168(.A(men_men_n1196_), .B(a), .Y(men_men_n1197_));
  OAI220     u1169(.A0(men_men_n1197_), .A1(men_men_n1195_), .B0(men_men_n953_), .B1(men_men_n456_), .Y(men_men_n1198_));
  NA2        u1170(.A(men_men_n545_), .B(l), .Y(men_men_n1199_));
  NOi31      u1171(.An(men_men_n930_), .B(men_men_n1114_), .C(men_men_n1199_), .Y(men_men_n1200_));
  NO4        u1172(.A(men_men_n1200_), .B(men_men_n1198_), .C(men_men_n1193_), .D(men_men_n1075_), .Y(men_men_n1201_));
  NO2        u1173(.A(men_men_n301_), .B(a), .Y(men_men_n1202_));
  INV        u1174(.A(men_men_n1120_), .Y(men_men_n1203_));
  NO2        u1175(.A(men_men_n1172_), .B(men_men_n520_), .Y(men_men_n1204_));
  NO2        u1176(.A(men_men_n89_), .B(g), .Y(men_men_n1205_));
  AOI210     u1177(.A0(men_men_n1205_), .A1(men_men_n1204_), .B0(men_men_n1155_), .Y(men_men_n1206_));
  OR2        u1178(.A(men_men_n1206_), .B(men_men_n1153_), .Y(men_men_n1207_));
  NA3        u1179(.A(men_men_n1207_), .B(men_men_n1203_), .C(men_men_n1201_), .Y(men_men_n1208_));
  NO4        u1180(.A(men_men_n1208_), .B(men_men_n1190_), .C(men_men_n885_), .D(men_men_n606_), .Y(men_men_n1209_));
  NA2        u1181(.A(c), .B(b), .Y(men_men_n1210_));
  NO2        u1182(.A(a), .B(men_men_n1210_), .Y(men_men_n1211_));
  OAI210     u1183(.A0(men_men_n928_), .A1(men_men_n900_), .B0(men_men_n443_), .Y(men_men_n1212_));
  OAI210     u1184(.A0(men_men_n1212_), .A1(men_men_n929_), .B0(men_men_n1211_), .Y(men_men_n1213_));
  NAi21      u1185(.An(men_men_n451_), .B(men_men_n1211_), .Y(men_men_n1214_));
  NA3        u1186(.A(men_men_n457_), .B(men_men_n599_), .C(f), .Y(men_men_n1215_));
  OAI210     u1187(.A0(men_men_n588_), .A1(men_men_n39_), .B0(men_men_n1202_), .Y(men_men_n1216_));
  NA3        u1188(.A(men_men_n1216_), .B(men_men_n1215_), .C(men_men_n1214_), .Y(men_men_n1217_));
  NA2        u1189(.A(men_men_n276_), .B(men_men_n123_), .Y(men_men_n1218_));
  OAI210     u1190(.A0(men_men_n1218_), .A1(men_men_n305_), .B0(g), .Y(men_men_n1219_));
  NAi21      u1191(.An(f), .B(d), .Y(men_men_n1220_));
  NO2        u1192(.A(men_men_n1220_), .B(men_men_n1176_), .Y(men_men_n1221_));
  INV        u1193(.A(men_men_n1221_), .Y(men_men_n1222_));
  AOI210     u1194(.A0(men_men_n1219_), .A1(men_men_n311_), .B0(men_men_n1222_), .Y(men_men_n1223_));
  AOI210     u1195(.A0(men_men_n1223_), .A1(men_men_n117_), .B0(men_men_n1217_), .Y(men_men_n1224_));
  NA2        u1196(.A(men_men_n503_), .B(men_men_n502_), .Y(men_men_n1225_));
  NO2        u1197(.A(men_men_n192_), .B(men_men_n250_), .Y(men_men_n1226_));
  NA2        u1198(.A(men_men_n1226_), .B(m), .Y(men_men_n1227_));
  NA3        u1199(.A(men_men_n988_), .B(men_men_n1199_), .C(men_men_n506_), .Y(men_men_n1228_));
  OAI210     u1200(.A0(men_men_n1228_), .A1(men_men_n332_), .B0(men_men_n504_), .Y(men_men_n1229_));
  AOI210     u1201(.A0(men_men_n1229_), .A1(men_men_n1225_), .B0(men_men_n1227_), .Y(men_men_n1230_));
  NA2        u1202(.A(men_men_n601_), .B(men_men_n438_), .Y(men_men_n1231_));
  NA2        u1203(.A(men_men_n166_), .B(men_men_n33_), .Y(men_men_n1232_));
  AOI210     u1204(.A0(men_men_n1037_), .A1(men_men_n1232_), .B0(men_men_n226_), .Y(men_men_n1233_));
  OAI210     u1205(.A0(men_men_n1233_), .A1(men_men_n477_), .B0(men_men_n1221_), .Y(men_men_n1234_));
  NO2        u1206(.A(men_men_n399_), .B(men_men_n398_), .Y(men_men_n1235_));
  AOI210     u1207(.A0(men_men_n1226_), .A1(men_men_n459_), .B0(men_men_n1032_), .Y(men_men_n1236_));
  NAi41      u1208(.An(men_men_n1235_), .B(men_men_n1236_), .C(men_men_n1234_), .D(men_men_n1231_), .Y(men_men_n1237_));
  NO2        u1209(.A(men_men_n1237_), .B(men_men_n1230_), .Y(men_men_n1238_));
  NA4        u1210(.A(men_men_n1238_), .B(men_men_n1224_), .C(men_men_n1213_), .D(men_men_n1209_), .Y(men00));
  AOI210     u1211(.A0(men_men_n318_), .A1(men_men_n226_), .B0(men_men_n293_), .Y(men_men_n1240_));
  NO2        u1212(.A(men_men_n1240_), .B(men_men_n620_), .Y(men_men_n1241_));
  AOI210     u1213(.A0(men_men_n968_), .A1(men_men_n1014_), .B0(men_men_n1193_), .Y(men_men_n1242_));
  NO3        u1214(.A(men_men_n1169_), .B(men_men_n1032_), .C(men_men_n766_), .Y(men_men_n1243_));
  NA3        u1215(.A(men_men_n1243_), .B(men_men_n1242_), .C(men_men_n1077_), .Y(men_men_n1244_));
  NA2        u1216(.A(men_men_n547_), .B(f), .Y(men_men_n1245_));
  OAI210     u1217(.A0(men_men_n1084_), .A1(men_men_n40_), .B0(men_men_n695_), .Y(men_men_n1246_));
  NA3        u1218(.A(men_men_n1246_), .B(men_men_n272_), .C(n), .Y(men_men_n1247_));
  AOI210     u1219(.A0(men_men_n1247_), .A1(men_men_n1245_), .B0(men_men_n1124_), .Y(men_men_n1248_));
  NO4        u1220(.A(men_men_n1248_), .B(men_men_n1244_), .C(men_men_n1241_), .D(men_men_n1147_), .Y(men_men_n1249_));
  NA3        u1221(.A(men_men_n176_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1250_));
  NA3        u1222(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1251_));
  NOi31      u1223(.An(n), .B(m), .C(i), .Y(men_men_n1252_));
  NA3        u1224(.A(men_men_n1252_), .B(men_men_n698_), .C(men_men_n51_), .Y(men_men_n1253_));
  OAI210     u1225(.A0(men_men_n1251_), .A1(men_men_n1250_), .B0(men_men_n1253_), .Y(men_men_n1254_));
  INV        u1226(.A(men_men_n619_), .Y(men_men_n1255_));
  NO4        u1227(.A(men_men_n1255_), .B(men_men_n1254_), .C(men_men_n1235_), .D(men_men_n991_), .Y(men_men_n1256_));
  NO4        u1228(.A(men_men_n523_), .B(men_men_n381_), .C(men_men_n1210_), .D(men_men_n59_), .Y(men_men_n1257_));
  NA3        u1229(.A(men_men_n411_), .B(men_men_n233_), .C(g), .Y(men_men_n1258_));
  OA220      u1230(.A0(men_men_n1258_), .A1(men_men_n1251_), .B0(men_men_n412_), .B1(men_men_n140_), .Y(men_men_n1259_));
  NO2        u1231(.A(h), .B(g), .Y(men_men_n1260_));
  NA4        u1232(.A(n), .B(men_men_n500_), .C(men_men_n1260_), .D(men_men_n1113_), .Y(men_men_n1261_));
  OAI220     u1233(.A0(men_men_n566_), .A1(men_men_n642_), .B0(men_men_n94_), .B1(men_men_n93_), .Y(men_men_n1262_));
  AOI220     u1234(.A0(men_men_n1262_), .A1(men_men_n575_), .B0(men_men_n1019_), .B1(men_men_n618_), .Y(men_men_n1263_));
  AOI220     u1235(.A0(men_men_n339_), .A1(men_men_n261_), .B0(men_men_n187_), .B1(men_men_n155_), .Y(men_men_n1264_));
  NA4        u1236(.A(men_men_n1264_), .B(men_men_n1263_), .C(men_men_n1261_), .D(men_men_n1259_), .Y(men_men_n1265_));
  NO3        u1237(.A(men_men_n1265_), .B(men_men_n1257_), .C(men_men_n282_), .Y(men_men_n1266_));
  INV        u1238(.A(men_men_n344_), .Y(men_men_n1267_));
  AOI210     u1239(.A0(men_men_n261_), .A1(men_men_n371_), .B0(men_men_n621_), .Y(men_men_n1268_));
  NA3        u1240(.A(men_men_n1268_), .B(men_men_n1267_), .C(men_men_n161_), .Y(men_men_n1269_));
  NO2        u1241(.A(men_men_n252_), .B(men_men_n191_), .Y(men_men_n1270_));
  NA2        u1242(.A(men_men_n1270_), .B(men_men_n457_), .Y(men_men_n1271_));
  NA3        u1243(.A(men_men_n189_), .B(men_men_n116_), .C(g), .Y(men_men_n1272_));
  NA3        u1244(.A(men_men_n500_), .B(men_men_n40_), .C(f), .Y(men_men_n1273_));
  NOi31      u1245(.An(men_men_n938_), .B(men_men_n1273_), .C(men_men_n1272_), .Y(men_men_n1274_));
  NAi31      u1246(.An(men_men_n196_), .B(men_men_n925_), .C(men_men_n500_), .Y(men_men_n1275_));
  NAi31      u1247(.An(men_men_n1274_), .B(men_men_n1275_), .C(men_men_n1271_), .Y(men_men_n1276_));
  NO2        u1248(.A(men_men_n292_), .B(men_men_n75_), .Y(men_men_n1277_));
  NO3        u1249(.A(men_men_n456_), .B(men_men_n896_), .C(n), .Y(men_men_n1278_));
  AOI210     u1250(.A0(men_men_n1278_), .A1(men_men_n1277_), .B0(men_men_n1162_), .Y(men_men_n1279_));
  NAi31      u1251(.An(men_men_n1127_), .B(men_men_n1279_), .C(men_men_n74_), .Y(men_men_n1280_));
  NO4        u1252(.A(men_men_n1280_), .B(men_men_n1276_), .C(men_men_n1269_), .D(men_men_n557_), .Y(men_men_n1281_));
  AN3        u1253(.A(men_men_n1281_), .B(men_men_n1266_), .C(men_men_n1256_), .Y(men_men_n1282_));
  NA2        u1254(.A(men_men_n575_), .B(men_men_n104_), .Y(men_men_n1283_));
  NA3        u1255(.A(men_men_n1194_), .B(men_men_n653_), .C(men_men_n499_), .Y(men_men_n1284_));
  NA4        u1256(.A(men_men_n1284_), .B(men_men_n602_), .C(men_men_n1283_), .D(men_men_n255_), .Y(men_men_n1285_));
  NA2        u1257(.A(men_men_n1187_), .B(men_men_n575_), .Y(men_men_n1286_));
  NA4        u1258(.A(men_men_n698_), .B(men_men_n217_), .C(men_men_n233_), .D(men_men_n170_), .Y(men_men_n1287_));
  NA3        u1259(.A(men_men_n1287_), .B(men_men_n1286_), .C(men_men_n315_), .Y(men_men_n1288_));
  OAI210     u1260(.A0(men_men_n498_), .A1(men_men_n124_), .B0(men_men_n931_), .Y(men_men_n1289_));
  AOI220     u1261(.A0(men_men_n1289_), .A1(men_men_n1228_), .B0(men_men_n601_), .B1(men_men_n438_), .Y(men_men_n1290_));
  OR4        u1262(.A(men_men_n1124_), .B(men_men_n288_), .C(men_men_n235_), .D(e), .Y(men_men_n1291_));
  NO2        u1263(.A(men_men_n229_), .B(men_men_n226_), .Y(men_men_n1292_));
  NA2        u1264(.A(n), .B(e), .Y(men_men_n1293_));
  NO2        u1265(.A(men_men_n1293_), .B(men_men_n153_), .Y(men_men_n1294_));
  AOI220     u1266(.A0(men_men_n1294_), .A1(men_men_n290_), .B0(men_men_n912_), .B1(men_men_n1292_), .Y(men_men_n1295_));
  OAI210     u1267(.A0(men_men_n382_), .A1(men_men_n333_), .B0(men_men_n479_), .Y(men_men_n1296_));
  NA4        u1268(.A(men_men_n1296_), .B(men_men_n1295_), .C(men_men_n1291_), .D(men_men_n1290_), .Y(men_men_n1297_));
  AOI210     u1269(.A0(men_men_n1294_), .A1(men_men_n916_), .B0(men_men_n884_), .Y(men_men_n1298_));
  AOI220     u1270(.A0(men_men_n1028_), .A1(men_men_n618_), .B0(men_men_n698_), .B1(men_men_n258_), .Y(men_men_n1299_));
  NO2        u1271(.A(men_men_n68_), .B(h), .Y(men_men_n1300_));
  NO3        u1272(.A(men_men_n1124_), .B(men_men_n1122_), .C(men_men_n782_), .Y(men_men_n1301_));
  NO2        u1273(.A(men_men_n1159_), .B(men_men_n137_), .Y(men_men_n1302_));
  AN2        u1274(.A(men_men_n1302_), .B(men_men_n1174_), .Y(men_men_n1303_));
  OAI210     u1275(.A0(men_men_n1303_), .A1(men_men_n1301_), .B0(men_men_n1300_), .Y(men_men_n1304_));
  NA4        u1276(.A(men_men_n1304_), .B(men_men_n1299_), .C(men_men_n1298_), .D(men_men_n933_), .Y(men_men_n1305_));
  NO4        u1277(.A(men_men_n1305_), .B(men_men_n1297_), .C(men_men_n1288_), .D(men_men_n1285_), .Y(men_men_n1306_));
  NA2        u1278(.A(men_men_n901_), .B(men_men_n815_), .Y(men_men_n1307_));
  NA4        u1279(.A(men_men_n1307_), .B(men_men_n1306_), .C(men_men_n1282_), .D(men_men_n1249_), .Y(men01));
  AN2        u1280(.A(men_men_n1102_), .B(men_men_n1100_), .Y(men_men_n1309_));
  NO4        u1281(.A(men_men_n864_), .B(men_men_n856_), .C(men_men_n514_), .D(men_men_n299_), .Y(men_men_n1310_));
  NO2        u1282(.A(men_men_n635_), .B(men_men_n308_), .Y(men_men_n1311_));
  OAI210     u1283(.A0(men_men_n1311_), .A1(men_men_n422_), .B0(i), .Y(men_men_n1312_));
  NA3        u1284(.A(men_men_n1312_), .B(men_men_n1310_), .C(men_men_n1309_), .Y(men_men_n1313_));
  NA2        u1285(.A(men_men_n631_), .B(men_men_n92_), .Y(men_men_n1314_));
  NA2        u1286(.A(men_men_n594_), .B(men_men_n287_), .Y(men_men_n1315_));
  NA2        u1287(.A(men_men_n1035_), .B(men_men_n1315_), .Y(men_men_n1316_));
  NA4        u1288(.A(men_men_n1316_), .B(men_men_n1314_), .C(men_men_n984_), .D(men_men_n356_), .Y(men_men_n1317_));
  NA2        u1289(.A(men_men_n45_), .B(f), .Y(men_men_n1318_));
  NA2        u1290(.A(men_men_n761_), .B(men_men_n99_), .Y(men_men_n1319_));
  OAI220     u1291(.A0(men_men_n1319_), .A1(men_men_n1318_), .B0(men_men_n378_), .B1(men_men_n303_), .Y(men_men_n1320_));
  OAI210     u1292(.A0(men_men_n842_), .A1(men_men_n648_), .B0(men_men_n1287_), .Y(men_men_n1321_));
  AOI210     u1293(.A0(men_men_n1320_), .A1(men_men_n684_), .B0(men_men_n1321_), .Y(men_men_n1322_));
  NA2        u1294(.A(men_men_n122_), .B(l), .Y(men_men_n1323_));
  OA220      u1295(.A0(men_men_n1323_), .A1(men_men_n628_), .B0(men_men_n711_), .B1(men_men_n396_), .Y(men_men_n1324_));
  NAi41      u1296(.An(men_men_n169_), .B(men_men_n1324_), .C(men_men_n1322_), .D(men_men_n967_), .Y(men_men_n1325_));
  NO3        u1297(.A(men_men_n843_), .B(men_men_n726_), .C(men_men_n550_), .Y(men_men_n1326_));
  NA4        u1298(.A(men_men_n761_), .B(men_men_n99_), .C(men_men_n45_), .D(men_men_n225_), .Y(men_men_n1327_));
  OA220      u1299(.A0(men_men_n1327_), .A1(men_men_n719_), .B0(men_men_n206_), .B1(men_men_n204_), .Y(men_men_n1328_));
  NA3        u1300(.A(men_men_n1328_), .B(men_men_n1326_), .C(men_men_n143_), .Y(men_men_n1329_));
  NO4        u1301(.A(men_men_n1329_), .B(men_men_n1325_), .C(men_men_n1317_), .D(men_men_n1313_), .Y(men_men_n1330_));
  NA2        u1302(.A(men_men_n1258_), .B(men_men_n218_), .Y(men_men_n1331_));
  OAI210     u1303(.A0(men_men_n1331_), .A1(men_men_n321_), .B0(men_men_n570_), .Y(men_men_n1332_));
  NA2        u1304(.A(men_men_n578_), .B(men_men_n424_), .Y(men_men_n1333_));
  NA2        u1305(.A(men_men_n76_), .B(i), .Y(men_men_n1334_));
  AOI210     u1306(.A0(men_men_n634_), .A1(men_men_n628_), .B0(men_men_n1334_), .Y(men_men_n1335_));
  NOi21      u1307(.An(men_men_n603_), .B(men_men_n625_), .Y(men_men_n1336_));
  AOI210     u1308(.A0(men_men_n1336_), .A1(men_men_n1333_), .B0(men_men_n1335_), .Y(men_men_n1337_));
  AOI210     u1309(.A0(men_men_n215_), .A1(men_men_n91_), .B0(men_men_n225_), .Y(men_men_n1338_));
  OAI210     u1310(.A0(men_men_n871_), .A1(men_men_n457_), .B0(men_men_n1338_), .Y(men_men_n1339_));
  AN3        u1311(.A(m), .B(l), .C(k), .Y(men_men_n1340_));
  OAI210     u1312(.A0(men_men_n384_), .A1(men_men_n34_), .B0(men_men_n1340_), .Y(men_men_n1341_));
  NA2        u1313(.A(men_men_n214_), .B(men_men_n34_), .Y(men_men_n1342_));
  AO210      u1314(.A0(men_men_n1342_), .A1(men_men_n1341_), .B0(men_men_n355_), .Y(men_men_n1343_));
  NA4        u1315(.A(men_men_n1343_), .B(men_men_n1339_), .C(men_men_n1337_), .D(men_men_n1332_), .Y(men_men_n1344_));
  AOI210     u1316(.A0(men_men_n640_), .A1(men_men_n122_), .B0(men_men_n646_), .Y(men_men_n1345_));
  OAI210     u1317(.A0(men_men_n1323_), .A1(men_men_n637_), .B0(men_men_n1345_), .Y(men_men_n1346_));
  NA2        u1318(.A(men_men_n298_), .B(men_men_n206_), .Y(men_men_n1347_));
  OAI210     u1319(.A0(men_men_n1347_), .A1(men_men_n413_), .B0(men_men_n716_), .Y(men_men_n1348_));
  NO3        u1320(.A(men_men_n883_), .B(men_men_n215_), .C(men_men_n436_), .Y(men_men_n1349_));
  NO2        u1321(.A(men_men_n1349_), .B(men_men_n1032_), .Y(men_men_n1350_));
  OAI210     u1322(.A0(men_men_n1320_), .A1(men_men_n349_), .B0(men_men_n727_), .Y(men_men_n1351_));
  NA4        u1323(.A(men_men_n1351_), .B(men_men_n1350_), .C(men_men_n1348_), .D(men_men_n846_), .Y(men_men_n1352_));
  NO3        u1324(.A(men_men_n1352_), .B(men_men_n1346_), .C(men_men_n1344_), .Y(men_men_n1353_));
  NA3        u1325(.A(men_men_n649_), .B(men_men_n29_), .C(f), .Y(men_men_n1354_));
  NO2        u1326(.A(men_men_n1354_), .B(men_men_n215_), .Y(men_men_n1355_));
  AOI210     u1327(.A0(men_men_n542_), .A1(men_men_n58_), .B0(men_men_n1355_), .Y(men_men_n1356_));
  OR3        u1328(.A(men_men_n1319_), .B(men_men_n650_), .C(men_men_n1318_), .Y(men_men_n1357_));
  NA3        u1329(.A(men_men_n796_), .B(men_men_n76_), .C(i), .Y(men_men_n1358_));
  AOI210     u1330(.A0(men_men_n1358_), .A1(men_men_n1327_), .B0(men_men_n1054_), .Y(men_men_n1359_));
  NO2        u1331(.A(men_men_n218_), .B(men_men_n115_), .Y(men_men_n1360_));
  NO3        u1332(.A(men_men_n1360_), .B(men_men_n1359_), .C(men_men_n1254_), .Y(men_men_n1361_));
  NA4        u1333(.A(men_men_n1361_), .B(men_men_n1357_), .C(men_men_n1356_), .D(men_men_n814_), .Y(men_men_n1362_));
  NO2        u1334(.A(men_men_n1041_), .B(men_men_n245_), .Y(men_men_n1363_));
  NO2        u1335(.A(men_men_n1042_), .B(men_men_n596_), .Y(men_men_n1364_));
  OAI210     u1336(.A0(men_men_n1364_), .A1(men_men_n1363_), .B0(men_men_n364_), .Y(men_men_n1365_));
  NA2        u1337(.A(men_men_n613_), .B(men_men_n611_), .Y(men_men_n1366_));
  NO3        u1338(.A(men_men_n81_), .B(men_men_n319_), .C(men_men_n45_), .Y(men_men_n1367_));
  NA2        u1339(.A(men_men_n1367_), .B(men_men_n593_), .Y(men_men_n1368_));
  NA3        u1340(.A(men_men_n1368_), .B(men_men_n1366_), .C(men_men_n721_), .Y(men_men_n1369_));
  OR2        u1341(.A(men_men_n1258_), .B(men_men_n1251_), .Y(men_men_n1370_));
  NO2        u1342(.A(men_men_n396_), .B(men_men_n73_), .Y(men_men_n1371_));
  AOI210     u1343(.A0(men_men_n787_), .A1(men_men_n664_), .B0(men_men_n1371_), .Y(men_men_n1372_));
  NA2        u1344(.A(men_men_n1367_), .B(men_men_n874_), .Y(men_men_n1373_));
  NA4        u1345(.A(men_men_n1373_), .B(men_men_n1372_), .C(men_men_n1370_), .D(men_men_n414_), .Y(men_men_n1374_));
  NOi41      u1346(.An(men_men_n1365_), .B(men_men_n1374_), .C(men_men_n1369_), .D(men_men_n1362_), .Y(men_men_n1375_));
  NO2        u1347(.A(men_men_n136_), .B(men_men_n45_), .Y(men_men_n1376_));
  AO220      u1348(.A0(i), .A1(men_men_n670_), .B0(men_men_n1376_), .B1(men_men_n759_), .Y(men_men_n1377_));
  NA2        u1349(.A(men_men_n1377_), .B(men_men_n364_), .Y(men_men_n1378_));
  NA2        u1350(.A(men_men_n493_), .B(men_men_n140_), .Y(men_men_n1379_));
  NO3        u1351(.A(men_men_n1172_), .B(men_men_n186_), .C(men_men_n89_), .Y(men_men_n1380_));
  AOI220     u1352(.A0(men_men_n1380_), .A1(men_men_n1379_), .B0(men_men_n1367_), .B1(men_men_n1045_), .Y(men_men_n1381_));
  NA2        u1353(.A(men_men_n1381_), .B(men_men_n1378_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n661_), .B(men_men_n660_), .Y(men_men_n1383_));
  NO4        u1355(.A(men_men_n1172_), .B(men_men_n1383_), .C(men_men_n184_), .D(men_men_n89_), .Y(men_men_n1384_));
  NO3        u1356(.A(men_men_n1384_), .B(men_men_n1382_), .C(men_men_n688_), .Y(men_men_n1385_));
  NA4        u1357(.A(men_men_n1385_), .B(men_men_n1375_), .C(men_men_n1353_), .D(men_men_n1330_), .Y(men06));
  NO2        u1358(.A(men_men_n437_), .B(men_men_n600_), .Y(men_men_n1387_));
  NO2        u1359(.A(men_men_n789_), .B(i), .Y(men_men_n1388_));
  OAI210     u1360(.A0(men_men_n1388_), .A1(men_men_n283_), .B0(men_men_n1387_), .Y(men_men_n1389_));
  NO2        u1361(.A(men_men_n237_), .B(men_men_n106_), .Y(men_men_n1390_));
  OAI210     u1362(.A0(men_men_n1390_), .A1(men_men_n1380_), .B0(men_men_n410_), .Y(men_men_n1391_));
  NO3        u1363(.A(men_men_n644_), .B(men_men_n869_), .C(men_men_n647_), .Y(men_men_n1392_));
  OR2        u1364(.A(men_men_n1392_), .B(men_men_n953_), .Y(men_men_n1393_));
  NA4        u1365(.A(men_men_n1393_), .B(men_men_n1391_), .C(men_men_n1389_), .D(men_men_n1365_), .Y(men_men_n1394_));
  NO3        u1366(.A(men_men_n1394_), .B(men_men_n1369_), .C(men_men_n271_), .Y(men_men_n1395_));
  NO2        u1367(.A(men_men_n319_), .B(men_men_n45_), .Y(men_men_n1396_));
  AOI210     u1368(.A0(men_men_n1396_), .A1(men_men_n1046_), .B0(men_men_n1363_), .Y(men_men_n1397_));
  AOI210     u1369(.A0(men_men_n1396_), .A1(men_men_n597_), .B0(men_men_n1377_), .Y(men_men_n1398_));
  AOI210     u1370(.A0(men_men_n1398_), .A1(men_men_n1397_), .B0(men_men_n361_), .Y(men_men_n1399_));
  OAI210     u1371(.A0(men_men_n91_), .A1(men_men_n40_), .B0(men_men_n725_), .Y(men_men_n1400_));
  NA2        u1372(.A(men_men_n1400_), .B(men_men_n387_), .Y(men_men_n1401_));
  NO2        u1373(.A(men_men_n553_), .B(men_men_n181_), .Y(men_men_n1402_));
  NOi21      u1374(.An(men_men_n142_), .B(men_men_n45_), .Y(men_men_n1403_));
  AOI210     u1375(.A0(men_men_n654_), .A1(men_men_n57_), .B0(men_men_n1195_), .Y(men_men_n1404_));
  OAI210     u1376(.A0(men_men_n493_), .A1(men_men_n262_), .B0(men_men_n978_), .Y(men_men_n1405_));
  NO4        u1377(.A(men_men_n1405_), .B(men_men_n1404_), .C(men_men_n1403_), .D(men_men_n1402_), .Y(men_men_n1406_));
  OR2        u1378(.A(men_men_n645_), .B(men_men_n643_), .Y(men_men_n1407_));
  NO2        u1379(.A(men_men_n395_), .B(men_men_n141_), .Y(men_men_n1408_));
  AOI210     u1380(.A0(men_men_n1408_), .A1(men_men_n631_), .B0(men_men_n1407_), .Y(men_men_n1409_));
  NA3        u1381(.A(men_men_n1409_), .B(men_men_n1406_), .C(men_men_n1401_), .Y(men_men_n1410_));
  NO2        u1382(.A(men_men_n805_), .B(men_men_n394_), .Y(men_men_n1411_));
  NO3        u1383(.A(men_men_n727_), .B(men_men_n816_), .C(men_men_n684_), .Y(men_men_n1412_));
  NOi21      u1384(.An(men_men_n1411_), .B(men_men_n1412_), .Y(men_men_n1413_));
  AN2        u1385(.A(men_men_n1028_), .B(men_men_n694_), .Y(men_men_n1414_));
  NO4        u1386(.A(men_men_n1414_), .B(men_men_n1413_), .C(men_men_n1410_), .D(men_men_n1399_), .Y(men_men_n1415_));
  NO2        u1387(.A(men_men_n863_), .B(men_men_n294_), .Y(men_men_n1416_));
  OAI220     u1388(.A0(men_men_n789_), .A1(men_men_n47_), .B0(men_men_n237_), .B1(men_men_n663_), .Y(men_men_n1417_));
  OAI210     u1389(.A0(men_men_n294_), .A1(c), .B0(men_men_n691_), .Y(men_men_n1418_));
  AOI220     u1390(.A0(men_men_n1418_), .A1(men_men_n1417_), .B0(men_men_n1416_), .B1(men_men_n283_), .Y(men_men_n1419_));
  NO3        u1391(.A(men_men_n257_), .B(men_men_n106_), .C(men_men_n301_), .Y(men_men_n1420_));
  OAI220     u1392(.A0(men_men_n752_), .A1(men_men_n262_), .B0(men_men_n549_), .B1(men_men_n553_), .Y(men_men_n1421_));
  OAI210     u1393(.A0(l), .A1(i), .B0(k), .Y(men_men_n1422_));
  NO3        u1394(.A(men_men_n1422_), .B(men_men_n642_), .C(j), .Y(men_men_n1423_));
  NOi21      u1395(.An(men_men_n1423_), .B(men_men_n719_), .Y(men_men_n1424_));
  NO4        u1396(.A(men_men_n1424_), .B(men_men_n1421_), .C(men_men_n1420_), .D(men_men_n1198_), .Y(men_men_n1425_));
  NA4        u1397(.A(men_men_n854_), .B(men_men_n853_), .C(men_men_n467_), .D(men_men_n945_), .Y(men_men_n1426_));
  NAi31      u1398(.An(men_men_n805_), .B(men_men_n1426_), .C(men_men_n214_), .Y(men_men_n1427_));
  NA4        u1399(.A(men_men_n1427_), .B(men_men_n1425_), .C(men_men_n1419_), .D(men_men_n1299_), .Y(men_men_n1428_));
  NOi31      u1400(.An(men_men_n1392_), .B(men_men_n497_), .C(men_men_n423_), .Y(men_men_n1429_));
  OR3        u1401(.A(men_men_n1429_), .B(men_men_n842_), .C(men_men_n581_), .Y(men_men_n1430_));
  OR3        u1402(.A(men_men_n398_), .B(men_men_n237_), .C(men_men_n663_), .Y(men_men_n1431_));
  AOI210     u1403(.A0(men_men_n613_), .A1(men_men_n479_), .B0(men_men_n400_), .Y(men_men_n1432_));
  NA2        u1404(.A(men_men_n1423_), .B(men_men_n850_), .Y(men_men_n1433_));
  NA4        u1405(.A(men_men_n1433_), .B(men_men_n1432_), .C(men_men_n1431_), .D(men_men_n1430_), .Y(men_men_n1434_));
  AOI220     u1406(.A0(men_men_n1411_), .A1(men_men_n815_), .B0(men_men_n1408_), .B1(men_men_n251_), .Y(men_men_n1435_));
  AO220      u1407(.A0(men_men_n1390_), .A1(men_men_n716_), .B0(men_men_n1000_), .B1(men_men_n999_), .Y(men_men_n1436_));
  NO4        u1408(.A(men_men_n1436_), .B(men_men_n943_), .C(men_men_n538_), .D(men_men_n517_), .Y(men_men_n1437_));
  NA3        u1409(.A(men_men_n1437_), .B(men_men_n1435_), .C(men_men_n1373_), .Y(men_men_n1438_));
  NAi21      u1410(.An(j), .B(i), .Y(men_men_n1439_));
  NO4        u1411(.A(men_men_n1383_), .B(men_men_n1439_), .C(men_men_n473_), .D(men_men_n248_), .Y(men_men_n1440_));
  NO4        u1412(.A(men_men_n1440_), .B(men_men_n1438_), .C(men_men_n1434_), .D(men_men_n1428_), .Y(men_men_n1441_));
  NA4        u1413(.A(men_men_n1441_), .B(men_men_n1415_), .C(men_men_n1395_), .D(men_men_n1385_), .Y(men07));
  NOi21      u1414(.An(j), .B(k), .Y(men_men_n1443_));
  NA4        u1415(.A(men_men_n189_), .B(men_men_n112_), .C(men_men_n1443_), .D(f), .Y(men_men_n1444_));
  NAi32      u1416(.An(m), .Bn(b), .C(n), .Y(men_men_n1445_));
  NO3        u1417(.A(men_men_n1445_), .B(g), .C(f), .Y(men_men_n1446_));
  OAI210     u1418(.A0(men_men_n343_), .A1(men_men_n519_), .B0(men_men_n1446_), .Y(men_men_n1447_));
  NAi21      u1419(.An(f), .B(c), .Y(men_men_n1448_));
  OR2        u1420(.A(e), .B(d), .Y(men_men_n1449_));
  OAI220     u1421(.A0(men_men_n1449_), .A1(men_men_n1448_), .B0(men_men_n676_), .B1(men_men_n345_), .Y(men_men_n1450_));
  NA3        u1422(.A(men_men_n1450_), .B(men_men_n1136_), .C(men_men_n189_), .Y(men_men_n1451_));
  NOi31      u1423(.An(n), .B(m), .C(b), .Y(men_men_n1452_));
  NO3        u1424(.A(men_men_n137_), .B(men_men_n481_), .C(h), .Y(men_men_n1453_));
  NA3        u1425(.A(men_men_n1451_), .B(men_men_n1447_), .C(men_men_n1444_), .Y(men_men_n1454_));
  NOi41      u1426(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1455_));
  NA3        u1427(.A(men_men_n1455_), .B(men_men_n935_), .C(men_men_n439_), .Y(men_men_n1456_));
  NOi21      u1428(.An(h), .B(k), .Y(men_men_n1457_));
  NO2        u1429(.A(men_men_n1456_), .B(men_men_n56_), .Y(men_men_n1458_));
  NO3        u1430(.A(men_men_n1130_), .B(men_men_n153_), .C(men_men_n226_), .Y(men_men_n1459_));
  OAI210     u1431(.A0(men_men_n1174_), .A1(men_men_n1459_), .B0(men_men_n233_), .Y(men_men_n1460_));
  NO2        u1432(.A(men_men_n1460_), .B(men_men_n61_), .Y(men_men_n1461_));
  NO2        u1433(.A(k), .B(i), .Y(men_men_n1462_));
  NA3        u1434(.A(men_men_n1462_), .B(men_men_n966_), .C(men_men_n189_), .Y(men_men_n1463_));
  NA2        u1435(.A(men_men_n89_), .B(men_men_n45_), .Y(men_men_n1464_));
  NO2        u1436(.A(men_men_n1130_), .B(men_men_n473_), .Y(men_men_n1465_));
  NA3        u1437(.A(men_men_n1465_), .B(men_men_n1464_), .C(men_men_n226_), .Y(men_men_n1466_));
  NO2        u1438(.A(men_men_n1144_), .B(men_men_n327_), .Y(men_men_n1467_));
  NA2        u1439(.A(men_men_n582_), .B(men_men_n82_), .Y(men_men_n1468_));
  NA2        u1440(.A(men_men_n1300_), .B(men_men_n309_), .Y(men_men_n1469_));
  NA4        u1441(.A(men_men_n1469_), .B(men_men_n1468_), .C(men_men_n1466_), .D(men_men_n1463_), .Y(men_men_n1470_));
  NO4        u1442(.A(men_men_n1470_), .B(men_men_n1461_), .C(men_men_n1458_), .D(men_men_n1454_), .Y(men_men_n1471_));
  NO3        u1443(.A(e), .B(d), .C(c), .Y(men_men_n1472_));
  AOI210     u1444(.A0(men_men_n1151_), .A1(men_men_n226_), .B0(men_men_n1472_), .Y(men_men_n1473_));
  OAI210     u1445(.A0(men_men_n137_), .A1(men_men_n226_), .B0(men_men_n651_), .Y(men_men_n1474_));
  NA2        u1446(.A(men_men_n1474_), .B(men_men_n1472_), .Y(men_men_n1475_));
  NO2        u1447(.A(men_men_n1475_), .B(men_men_n1473_), .Y(men_men_n1476_));
  OR2        u1448(.A(h), .B(f), .Y(men_men_n1477_));
  NO3        u1449(.A(n), .B(m), .C(i), .Y(men_men_n1478_));
  OAI210     u1450(.A0(men_men_n1196_), .A1(men_men_n164_), .B0(men_men_n1478_), .Y(men_men_n1479_));
  NO2        u1451(.A(i), .B(g), .Y(men_men_n1480_));
  OR3        u1452(.A(men_men_n1480_), .B(men_men_n1445_), .C(men_men_n72_), .Y(men_men_n1481_));
  OAI220     u1453(.A0(men_men_n1481_), .A1(men_men_n519_), .B0(men_men_n1479_), .B1(men_men_n1477_), .Y(men_men_n1482_));
  NA3        u1454(.A(men_men_n749_), .B(men_men_n735_), .C(men_men_n116_), .Y(men_men_n1483_));
  NA3        u1455(.A(men_men_n1452_), .B(men_men_n1139_), .C(men_men_n723_), .Y(men_men_n1484_));
  AOI210     u1456(.A0(men_men_n1484_), .A1(men_men_n1483_), .B0(men_men_n45_), .Y(men_men_n1485_));
  NA2        u1457(.A(men_men_n1478_), .B(men_men_n690_), .Y(men_men_n1486_));
  NO2        u1458(.A(l), .B(k), .Y(men_men_n1487_));
  NOi41      u1459(.An(men_men_n586_), .B(men_men_n1487_), .C(men_men_n512_), .D(men_men_n473_), .Y(men_men_n1488_));
  NO3        u1460(.A(men_men_n473_), .B(d), .C(c), .Y(men_men_n1489_));
  NO4        u1461(.A(men_men_n1488_), .B(men_men_n1485_), .C(men_men_n1482_), .D(men_men_n1476_), .Y(men_men_n1490_));
  NO2        u1462(.A(men_men_n154_), .B(h), .Y(men_men_n1491_));
  NO2        u1463(.A(g), .B(c), .Y(men_men_n1492_));
  NA3        u1464(.A(men_men_n1492_), .B(men_men_n148_), .C(men_men_n197_), .Y(men_men_n1493_));
  NO2        u1465(.A(men_men_n1493_), .B(men_men_n1668_), .Y(men_men_n1494_));
  NA2        u1466(.A(men_men_n1494_), .B(men_men_n189_), .Y(men_men_n1495_));
  OAI210     u1467(.A0(men_men_n1457_), .A1(men_men_n225_), .B0(men_men_n1154_), .Y(men_men_n1496_));
  NO2        u1468(.A(men_men_n484_), .B(a), .Y(men_men_n1497_));
  NA3        u1469(.A(men_men_n1497_), .B(men_men_n1496_), .C(men_men_n117_), .Y(men_men_n1498_));
  NO2        u1470(.A(i), .B(h), .Y(men_men_n1499_));
  NA2        u1471(.A(men_men_n1499_), .B(men_men_n233_), .Y(men_men_n1500_));
  AOI210     u1472(.A0(men_men_n272_), .A1(men_men_n120_), .B0(men_men_n570_), .Y(men_men_n1501_));
  NO2        u1473(.A(men_men_n1501_), .B(men_men_n1500_), .Y(men_men_n1502_));
  NO2        u1474(.A(men_men_n812_), .B(men_men_n198_), .Y(men_men_n1503_));
  NOi31      u1475(.An(m), .B(n), .C(b), .Y(men_men_n1504_));
  NOi31      u1476(.An(f), .B(d), .C(c), .Y(men_men_n1505_));
  NA2        u1477(.A(men_men_n1505_), .B(men_men_n1504_), .Y(men_men_n1506_));
  INV        u1478(.A(men_men_n1506_), .Y(men_men_n1507_));
  NO3        u1479(.A(men_men_n1507_), .B(men_men_n1503_), .C(men_men_n1502_), .Y(men_men_n1508_));
  NA2        u1480(.A(men_men_n1165_), .B(men_men_n500_), .Y(men_men_n1509_));
  NO4        u1481(.A(men_men_n1509_), .B(men_men_n1139_), .C(men_men_n473_), .D(men_men_n45_), .Y(men_men_n1510_));
  NO3        u1482(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1511_));
  INV        u1483(.A(men_men_n1510_), .Y(men_men_n1512_));
  AN4        u1484(.A(men_men_n1512_), .B(men_men_n1508_), .C(men_men_n1498_), .D(men_men_n1495_), .Y(men_men_n1513_));
  NA2        u1485(.A(men_men_n1452_), .B(men_men_n407_), .Y(men_men_n1514_));
  NO2        u1486(.A(men_men_n1514_), .B(men_men_n1121_), .Y(men_men_n1515_));
  NA2        u1487(.A(men_men_n1489_), .B(men_men_n227_), .Y(men_men_n1516_));
  NO2        u1488(.A(men_men_n198_), .B(b), .Y(men_men_n1517_));
  AOI220     u1489(.A0(men_men_n1252_), .A1(men_men_n1517_), .B0(men_men_n1173_), .B1(men_men_n1509_), .Y(men_men_n1518_));
  NO2        u1490(.A(i), .B(men_men_n225_), .Y(men_men_n1519_));
  NA4        u1491(.A(men_men_n1226_), .B(men_men_n1519_), .C(men_men_n107_), .D(m), .Y(men_men_n1520_));
  NAi41      u1492(.An(men_men_n1515_), .B(men_men_n1520_), .C(men_men_n1518_), .D(men_men_n1516_), .Y(men_men_n1521_));
  NO4        u1493(.A(men_men_n137_), .B(g), .C(f), .D(e), .Y(men_men_n1522_));
  NA3        u1494(.A(men_men_n1462_), .B(men_men_n310_), .C(h), .Y(men_men_n1523_));
  NA2        u1495(.A(men_men_n205_), .B(men_men_n101_), .Y(men_men_n1524_));
  OR2        u1496(.A(e), .B(a), .Y(men_men_n1525_));
  NO2        u1497(.A(men_men_n1449_), .B(men_men_n1448_), .Y(men_men_n1526_));
  AOI210     u1498(.A0(men_men_n30_), .A1(h), .B0(men_men_n1526_), .Y(men_men_n1527_));
  NO2        u1499(.A(men_men_n1527_), .B(men_men_n1161_), .Y(men_men_n1528_));
  NOi41      u1500(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1529_));
  NA2        u1501(.A(men_men_n1529_), .B(men_men_n117_), .Y(men_men_n1530_));
  INV        u1502(.A(men_men_n1530_), .Y(men_men_n1531_));
  OR3        u1503(.A(men_men_n581_), .B(men_men_n580_), .C(men_men_n116_), .Y(men_men_n1532_));
  NA2        u1504(.A(men_men_n1194_), .B(men_men_n436_), .Y(men_men_n1533_));
  OAI220     u1505(.A0(men_men_n1533_), .A1(men_men_n466_), .B0(men_men_n1532_), .B1(men_men_n319_), .Y(men_men_n1534_));
  AO210      u1506(.A0(men_men_n1534_), .A1(men_men_n120_), .B0(men_men_n1531_), .Y(men_men_n1535_));
  NO3        u1507(.A(men_men_n1535_), .B(men_men_n1528_), .C(men_men_n1521_), .Y(men_men_n1536_));
  NA4        u1508(.A(men_men_n1536_), .B(men_men_n1513_), .C(men_men_n1490_), .D(men_men_n1471_), .Y(men_men_n1537_));
  NO2        u1509(.A(men_men_n1210_), .B(men_men_n114_), .Y(men_men_n1538_));
  NA2        u1510(.A(men_men_n407_), .B(men_men_n56_), .Y(men_men_n1539_));
  AOI210     u1511(.A0(men_men_n1539_), .A1(men_men_n1130_), .B0(men_men_n1486_), .Y(men_men_n1540_));
  NA2        u1512(.A(men_men_n227_), .B(men_men_n189_), .Y(men_men_n1541_));
  AOI210     u1513(.A0(men_men_n1541_), .A1(men_men_n1272_), .B0(men_men_n1539_), .Y(men_men_n1542_));
  NO2        u1514(.A(men_men_n1166_), .B(men_men_n1161_), .Y(men_men_n1543_));
  NO3        u1515(.A(men_men_n1543_), .B(men_men_n1542_), .C(men_men_n1540_), .Y(men_men_n1544_));
  NO2        u1516(.A(men_men_n419_), .B(j), .Y(men_men_n1545_));
  NA3        u1517(.A(men_men_n1511_), .B(men_men_n1449_), .C(men_men_n1194_), .Y(men_men_n1546_));
  NAi41      u1518(.An(men_men_n1499_), .B(men_men_n1152_), .C(men_men_n177_), .D(men_men_n157_), .Y(men_men_n1547_));
  NA2        u1519(.A(men_men_n1547_), .B(men_men_n1546_), .Y(men_men_n1548_));
  NA3        u1520(.A(g), .B(men_men_n1545_), .C(men_men_n166_), .Y(men_men_n1549_));
  INV        u1521(.A(men_men_n1549_), .Y(men_men_n1550_));
  NO2        u1522(.A(men_men_n1550_), .B(men_men_n1548_), .Y(men_men_n1551_));
  NO3        u1523(.A(men_men_n1161_), .B(men_men_n625_), .C(g), .Y(men_men_n1552_));
  NOi21      u1524(.An(men_men_n1541_), .B(men_men_n1552_), .Y(men_men_n1553_));
  AOI210     u1525(.A0(men_men_n1553_), .A1(men_men_n1524_), .B0(men_men_n1130_), .Y(men_men_n1554_));
  OAI220     u1526(.A0(men_men_n717_), .A1(g), .B0(men_men_n237_), .B1(c), .Y(men_men_n1555_));
  AOI210     u1527(.A0(men_men_n1517_), .A1(men_men_n41_), .B0(men_men_n1555_), .Y(men_men_n1556_));
  NO2        u1528(.A(men_men_n137_), .B(l), .Y(men_men_n1557_));
  NO2        u1529(.A(men_men_n237_), .B(k), .Y(men_men_n1558_));
  OAI210     u1530(.A0(men_men_n1558_), .A1(men_men_n1499_), .B0(men_men_n1557_), .Y(men_men_n1559_));
  OAI220     u1531(.A0(men_men_n1559_), .A1(men_men_n31_), .B0(men_men_n1556_), .B1(men_men_n186_), .Y(men_men_n1560_));
  NO3        u1532(.A(men_men_n1532_), .B(men_men_n500_), .C(men_men_n378_), .Y(men_men_n1561_));
  NO3        u1533(.A(men_men_n1561_), .B(men_men_n1560_), .C(men_men_n1554_), .Y(men_men_n1562_));
  NO2        u1534(.A(men_men_n49_), .B(men_men_n625_), .Y(men_men_n1563_));
  NO3        u1535(.A(men_men_n1176_), .B(men_men_n1449_), .C(men_men_n49_), .Y(men_men_n1564_));
  AOI220     u1536(.A0(men_men_n1564_), .A1(men_men_n226_), .B0(men_men_n1177_), .B1(men_men_n1563_), .Y(men_men_n1565_));
  NO2        u1537(.A(men_men_n1161_), .B(h), .Y(men_men_n1566_));
  NA3        u1538(.A(men_men_n1566_), .B(d), .C(men_men_n1122_), .Y(men_men_n1567_));
  OAI220     u1539(.A0(men_men_n1567_), .A1(c), .B0(men_men_n1565_), .B1(j), .Y(men_men_n1568_));
  NA3        u1540(.A(men_men_n1538_), .B(men_men_n500_), .C(f), .Y(men_men_n1569_));
  NA2        u1541(.A(men_men_n189_), .B(men_men_n116_), .Y(men_men_n1570_));
  NO2        u1542(.A(men_men_n1443_), .B(men_men_n42_), .Y(men_men_n1571_));
  AOI210     u1543(.A0(men_men_n117_), .A1(men_men_n40_), .B0(men_men_n1571_), .Y(men_men_n1572_));
  NO2        u1544(.A(men_men_n1572_), .B(men_men_n1569_), .Y(men_men_n1573_));
  AOI210     u1545(.A0(men_men_n565_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1574_));
  NA2        u1546(.A(men_men_n1574_), .B(men_men_n1497_), .Y(men_men_n1575_));
  NO2        u1547(.A(men_men_n1439_), .B(men_men_n184_), .Y(men_men_n1576_));
  NOi21      u1548(.An(d), .B(f), .Y(men_men_n1577_));
  NO3        u1549(.A(men_men_n1505_), .B(men_men_n1577_), .C(men_men_n40_), .Y(men_men_n1578_));
  NA2        u1550(.A(men_men_n1578_), .B(men_men_n1576_), .Y(men_men_n1579_));
  NO2        u1551(.A(men_men_n1449_), .B(f), .Y(men_men_n1580_));
  NA2        u1552(.A(men_men_n1497_), .B(men_men_n1571_), .Y(men_men_n1581_));
  NO2        u1553(.A(men_men_n319_), .B(c), .Y(men_men_n1582_));
  NA2        u1554(.A(men_men_n1582_), .B(men_men_n582_), .Y(men_men_n1583_));
  NA4        u1555(.A(men_men_n1583_), .B(men_men_n1581_), .C(men_men_n1579_), .D(men_men_n1575_), .Y(men_men_n1584_));
  NO3        u1556(.A(men_men_n1584_), .B(men_men_n1573_), .C(men_men_n1568_), .Y(men_men_n1585_));
  NA4        u1557(.A(men_men_n1585_), .B(men_men_n1562_), .C(men_men_n1551_), .D(men_men_n1544_), .Y(men_men_n1586_));
  NO3        u1558(.A(men_men_n1165_), .B(men_men_n1151_), .C(men_men_n40_), .Y(men_men_n1587_));
  OAI220     u1559(.A0(men_men_n500_), .A1(men_men_n319_), .B0(men_men_n136_), .B1(men_men_n59_), .Y(men_men_n1588_));
  OAI210     u1560(.A0(men_men_n1588_), .A1(men_men_n1587_), .B0(men_men_n1467_), .Y(men_men_n1589_));
  OAI220     u1561(.A0(men_men_n1118_), .A1(men_men_n137_), .B0(men_men_n717_), .B1(men_men_n184_), .Y(men_men_n1590_));
  NA2        u1562(.A(men_men_n1590_), .B(men_men_n669_), .Y(men_men_n1591_));
  NA2        u1563(.A(men_men_n1591_), .B(men_men_n1589_), .Y(men_men_n1592_));
  NA2        u1564(.A(men_men_n1492_), .B(men_men_n1577_), .Y(men_men_n1593_));
  NO2        u1565(.A(men_men_n1593_), .B(m), .Y(men_men_n1594_));
  NA3        u1566(.A(men_men_n1174_), .B(men_men_n112_), .C(men_men_n233_), .Y(men_men_n1595_));
  OAI220     u1567(.A0(men_men_n158_), .A1(men_men_n191_), .B0(men_men_n481_), .B1(g), .Y(men_men_n1596_));
  OAI210     u1568(.A0(men_men_n1596_), .A1(men_men_n114_), .B0(men_men_n1504_), .Y(men_men_n1597_));
  NA2        u1569(.A(men_men_n1597_), .B(men_men_n1595_), .Y(men_men_n1598_));
  NO3        u1570(.A(men_men_n1598_), .B(men_men_n1594_), .C(men_men_n1592_), .Y(men_men_n1599_));
  NO2        u1571(.A(men_men_n1448_), .B(e), .Y(men_men_n1600_));
  NA2        u1572(.A(men_men_n1600_), .B(men_men_n434_), .Y(men_men_n1601_));
  NA2        u1573(.A(men_men_n1205_), .B(men_men_n680_), .Y(men_men_n1602_));
  OR3        u1574(.A(men_men_n1558_), .B(men_men_n1300_), .C(men_men_n137_), .Y(men_men_n1603_));
  OAI220     u1575(.A0(men_men_n1603_), .A1(men_men_n1601_), .B0(men_men_n1602_), .B1(men_men_n475_), .Y(men_men_n1604_));
  NO3        u1576(.A(men_men_n1532_), .B(men_men_n378_), .C(a), .Y(men_men_n1605_));
  NO2        u1577(.A(men_men_n1605_), .B(men_men_n1604_), .Y(men_men_n1606_));
  NO2        u1578(.A(men_men_n191_), .B(c), .Y(men_men_n1607_));
  OAI210     u1579(.A0(men_men_n1607_), .A1(men_men_n1600_), .B0(men_men_n189_), .Y(men_men_n1608_));
  AOI220     u1580(.A0(men_men_n1608_), .A1(men_men_n1153_), .B0(men_men_n572_), .B1(men_men_n394_), .Y(men_men_n1609_));
  NA2        u1581(.A(men_men_n580_), .B(g), .Y(men_men_n1610_));
  AOI210     u1582(.A0(men_men_n1610_), .A1(men_men_n1489_), .B0(men_men_n1564_), .Y(men_men_n1611_));
  NO2        u1583(.A(men_men_n1525_), .B(f), .Y(men_men_n1612_));
  AOI210     u1584(.A0(men_men_n1205_), .A1(a), .B0(men_men_n1612_), .Y(men_men_n1613_));
  OAI220     u1585(.A0(men_men_n1613_), .A1(men_men_n69_), .B0(men_men_n1611_), .B1(men_men_n225_), .Y(men_men_n1614_));
  AOI210     u1586(.A0(men_men_n971_), .A1(men_men_n446_), .B0(men_men_n108_), .Y(men_men_n1615_));
  OR2        u1587(.A(men_men_n1615_), .B(men_men_n580_), .Y(men_men_n1616_));
  NA2        u1588(.A(men_men_n1612_), .B(men_men_n1464_), .Y(men_men_n1617_));
  OAI220     u1589(.A0(men_men_n1617_), .A1(men_men_n49_), .B0(men_men_n1616_), .B1(men_men_n184_), .Y(men_men_n1618_));
  NA4        u1590(.A(men_men_n1174_), .B(men_men_n1171_), .C(men_men_n233_), .D(men_men_n68_), .Y(men_men_n1619_));
  NA2        u1591(.A(men_men_n1453_), .B(men_men_n192_), .Y(men_men_n1620_));
  NO2        u1592(.A(men_men_n49_), .B(l), .Y(men_men_n1621_));
  OAI210     u1593(.A0(men_men_n1525_), .A1(men_men_n927_), .B0(men_men_n519_), .Y(men_men_n1622_));
  OAI210     u1594(.A0(men_men_n1622_), .A1(men_men_n1177_), .B0(men_men_n1621_), .Y(men_men_n1623_));
  NO2        u1595(.A(men_men_n267_), .B(g), .Y(men_men_n1624_));
  NO2        u1596(.A(m), .B(i), .Y(men_men_n1625_));
  AOI220     u1597(.A0(men_men_n1625_), .A1(men_men_n1491_), .B0(men_men_n1152_), .B1(men_men_n1624_), .Y(men_men_n1626_));
  NA4        u1598(.A(men_men_n1626_), .B(men_men_n1623_), .C(men_men_n1620_), .D(men_men_n1619_), .Y(men_men_n1627_));
  NO4        u1599(.A(men_men_n1627_), .B(men_men_n1618_), .C(men_men_n1614_), .D(men_men_n1609_), .Y(men_men_n1628_));
  NA3        u1600(.A(men_men_n1628_), .B(men_men_n1606_), .C(men_men_n1599_), .Y(men_men_n1629_));
  NA3        u1601(.A(men_men_n1034_), .B(men_men_n144_), .C(men_men_n46_), .Y(men_men_n1630_));
  AOI210     u1602(.A0(men_men_n155_), .A1(c), .B0(men_men_n1630_), .Y(men_men_n1631_));
  OAI210     u1603(.A0(men_men_n625_), .A1(g), .B0(men_men_n195_), .Y(men_men_n1632_));
  NA2        u1604(.A(men_men_n1632_), .B(men_men_n1566_), .Y(men_men_n1633_));
  AO210      u1605(.A0(men_men_n138_), .A1(l), .B0(men_men_n1514_), .Y(men_men_n1634_));
  NO2        u1606(.A(men_men_n72_), .B(c), .Y(men_men_n1635_));
  NO4        u1607(.A(men_men_n1477_), .B(men_men_n196_), .C(men_men_n481_), .D(men_men_n45_), .Y(men_men_n1636_));
  AOI210     u1608(.A0(men_men_n1576_), .A1(men_men_n1635_), .B0(men_men_n1636_), .Y(men_men_n1637_));
  NA3        u1609(.A(men_men_n1637_), .B(men_men_n1634_), .C(men_men_n1633_), .Y(men_men_n1638_));
  NO2        u1610(.A(men_men_n1638_), .B(men_men_n1631_), .Y(men_men_n1639_));
  NO4        u1611(.A(men_men_n237_), .B(men_men_n196_), .C(men_men_n272_), .D(k), .Y(men_men_n1640_));
  AOI210     u1612(.A0(men_men_n164_), .A1(men_men_n56_), .B0(men_men_n1600_), .Y(men_men_n1641_));
  NO2        u1613(.A(men_men_n1641_), .B(men_men_n1570_), .Y(men_men_n1642_));
  NO2        u1614(.A(men_men_n1630_), .B(men_men_n114_), .Y(men_men_n1643_));
  NOi21      u1615(.An(men_men_n1453_), .B(e), .Y(men_men_n1644_));
  NO4        u1616(.A(men_men_n1644_), .B(men_men_n1643_), .C(men_men_n1642_), .D(men_men_n1640_), .Y(men_men_n1645_));
  AO220      u1617(.A0(men_men_n1174_), .A1(men_men_n1159_), .B0(men_men_n1459_), .B1(men_men_n820_), .Y(men_men_n1646_));
  AOI220     u1618(.A0(men_men_n1625_), .A1(men_men_n690_), .B0(men_men_n1136_), .B1(men_men_n167_), .Y(men_men_n1647_));
  NOi31      u1619(.An(men_men_n30_), .B(men_men_n1647_), .C(n), .Y(men_men_n1648_));
  AOI210     u1620(.A0(men_men_n1646_), .A1(men_men_n1252_), .B0(men_men_n1648_), .Y(men_men_n1649_));
  NO2        u1621(.A(men_men_n1569_), .B(men_men_n69_), .Y(men_men_n1650_));
  NA2        u1622(.A(men_men_n59_), .B(a), .Y(men_men_n1651_));
  NO2        u1623(.A(men_men_n1462_), .B(men_men_n122_), .Y(men_men_n1652_));
  OAI220     u1624(.A0(men_men_n1652_), .A1(men_men_n1514_), .B0(men_men_n1533_), .B1(men_men_n1651_), .Y(men_men_n1653_));
  NO2        u1625(.A(men_men_n1653_), .B(men_men_n1650_), .Y(men_men_n1654_));
  NA4        u1626(.A(men_men_n1654_), .B(men_men_n1649_), .C(men_men_n1645_), .D(men_men_n1639_), .Y(men_men_n1655_));
  OR4        u1627(.A(men_men_n1655_), .B(men_men_n1629_), .C(men_men_n1586_), .D(men_men_n1537_), .Y(men04));
  NOi31      u1628(.An(men_men_n1522_), .B(men_men_n1523_), .C(men_men_n1124_), .Y(men_men_n1657_));
  NA2        u1629(.A(men_men_n1580_), .B(men_men_n888_), .Y(men_men_n1658_));
  NO4        u1630(.A(men_men_n1658_), .B(men_men_n1114_), .C(men_men_n520_), .D(j), .Y(men_men_n1659_));
  OR3        u1631(.A(men_men_n1659_), .B(men_men_n1657_), .C(men_men_n1142_), .Y(men_men_n1660_));
  NO3        u1632(.A(men_men_n1464_), .B(men_men_n93_), .C(k), .Y(men_men_n1661_));
  AOI210     u1633(.A0(men_men_n1661_), .A1(men_men_n1135_), .B0(men_men_n1274_), .Y(men_men_n1662_));
  NA2        u1634(.A(men_men_n1662_), .B(men_men_n1304_), .Y(men_men_n1663_));
  NO4        u1635(.A(men_men_n1663_), .B(men_men_n1660_), .C(men_men_n1150_), .D(men_men_n1129_), .Y(men_men_n1664_));
  NA4        u1636(.A(men_men_n1664_), .B(men_men_n1207_), .C(men_men_n1192_), .D(men_men_n1180_), .Y(men05));
  INV        u1637(.A(l), .Y(men_men_n1668_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule