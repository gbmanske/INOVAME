//Benchmark atmr_alu4_1266_0.0625

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n136_, ori_ori_n137_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n56_));
  NO2        o034(.A(i_1_), .B(i_6_), .Y(ori_ori_n57_));
  NA2        o035(.A(i_8_), .B(i_7_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n57_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(i_12_), .Y(ori_ori_n60_));
  NAi21      o038(.An(i_2_), .B(i_7_), .Y(ori_ori_n61_));
  INV        o039(.A(i_1_), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n62_), .B(i_6_), .Y(ori_ori_n63_));
  NA3        o041(.A(ori_ori_n63_), .B(ori_ori_n61_), .C(ori_ori_n31_), .Y(ori_ori_n64_));
  NA2        o042(.A(i_1_), .B(i_10_), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n65_), .B(i_6_), .Y(ori_ori_n66_));
  NAi31      o044(.An(ori_ori_n66_), .B(ori_ori_n64_), .C(ori_ori_n60_), .Y(ori_ori_n67_));
  NA2        o045(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n69_));
  NA2        o047(.A(i_1_), .B(i_6_), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n70_), .B(ori_ori_n25_), .Y(ori_ori_n71_));
  INV        o049(.A(i_0_), .Y(ori_ori_n72_));
  NAi21      o050(.An(i_5_), .B(i_10_), .Y(ori_ori_n73_));
  NA2        o051(.A(i_5_), .B(i_9_), .Y(ori_ori_n74_));
  AOI210     o052(.A0(ori_ori_n74_), .A1(ori_ori_n73_), .B0(ori_ori_n72_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n75_), .B(ori_ori_n71_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n69_), .A1(ori_ori_n68_), .B0(ori_ori_n76_), .Y(ori_ori_n77_));
  OAI210     o055(.A0(ori_ori_n77_), .A1(ori_ori_n67_), .B0(i_0_), .Y(ori_ori_n78_));
  NA2        o056(.A(i_12_), .B(i_5_), .Y(ori_ori_n79_));
  NA2        o057(.A(i_2_), .B(i_8_), .Y(ori_ori_n80_));
  NO2        o058(.A(ori_ori_n80_), .B(ori_ori_n57_), .Y(ori_ori_n81_));
  NO2        o059(.A(i_3_), .B(i_9_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_3_), .B(i_7_), .Y(ori_ori_n83_));
  NO2        o061(.A(ori_ori_n82_), .B(ori_ori_n62_), .Y(ori_ori_n84_));
  INV        o062(.A(i_6_), .Y(ori_ori_n85_));
  NO2        o063(.A(i_2_), .B(i_7_), .Y(ori_ori_n86_));
  INV        o064(.A(ori_ori_n86_), .Y(ori_ori_n87_));
  OAI210     o065(.A0(ori_ori_n84_), .A1(ori_ori_n81_), .B0(ori_ori_n87_), .Y(ori_ori_n88_));
  NAi21      o066(.An(i_6_), .B(i_10_), .Y(ori_ori_n89_));
  NA2        o067(.A(i_6_), .B(i_9_), .Y(ori_ori_n90_));
  AOI210     o068(.A0(ori_ori_n90_), .A1(ori_ori_n89_), .B0(ori_ori_n62_), .Y(ori_ori_n91_));
  NA2        o069(.A(i_2_), .B(i_6_), .Y(ori_ori_n92_));
  INV        o070(.A(ori_ori_n91_), .Y(ori_ori_n93_));
  AOI210     o071(.A0(ori_ori_n93_), .A1(ori_ori_n88_), .B0(ori_ori_n79_), .Y(ori_ori_n94_));
  AN3        o072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n95_));
  NAi21      o073(.An(i_6_), .B(i_11_), .Y(ori_ori_n96_));
  NO2        o074(.A(i_5_), .B(i_8_), .Y(ori_ori_n97_));
  NOi21      o075(.An(ori_ori_n97_), .B(ori_ori_n96_), .Y(ori_ori_n98_));
  AOI220     o076(.A0(ori_ori_n98_), .A1(ori_ori_n61_), .B0(ori_ori_n95_), .B1(ori_ori_n32_), .Y(ori_ori_n99_));
  INV        o077(.A(i_7_), .Y(ori_ori_n100_));
  NA2        o078(.A(ori_ori_n46_), .B(ori_ori_n100_), .Y(ori_ori_n101_));
  NO2        o079(.A(i_0_), .B(i_5_), .Y(ori_ori_n102_));
  NO2        o080(.A(ori_ori_n102_), .B(ori_ori_n85_), .Y(ori_ori_n103_));
  NA2        o081(.A(i_12_), .B(i_3_), .Y(ori_ori_n104_));
  INV        o082(.A(ori_ori_n104_), .Y(ori_ori_n105_));
  NA3        o083(.A(ori_ori_n105_), .B(ori_ori_n103_), .C(ori_ori_n101_), .Y(ori_ori_n106_));
  NAi21      o084(.An(i_7_), .B(i_11_), .Y(ori_ori_n107_));
  AN2        o085(.A(i_2_), .B(i_10_), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n108_), .B(i_7_), .Y(ori_ori_n109_));
  OR2        o087(.A(ori_ori_n79_), .B(ori_ori_n57_), .Y(ori_ori_n110_));
  NO2        o088(.A(i_8_), .B(ori_ori_n100_), .Y(ori_ori_n111_));
  NO3        o089(.A(ori_ori_n111_), .B(ori_ori_n110_), .C(ori_ori_n109_), .Y(ori_ori_n112_));
  NA2        o090(.A(i_12_), .B(i_7_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n62_), .B(ori_ori_n26_), .Y(ori_ori_n114_));
  NA2        o092(.A(i_11_), .B(i_12_), .Y(ori_ori_n115_));
  INV        o093(.A(ori_ori_n115_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n116_), .B(ori_ori_n112_), .Y(ori_ori_n117_));
  NA3        o095(.A(ori_ori_n117_), .B(ori_ori_n106_), .C(ori_ori_n99_), .Y(ori_ori_n118_));
  NOi21      o096(.An(i_1_), .B(i_5_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(i_11_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n100_), .B(ori_ori_n37_), .Y(ori_ori_n121_));
  NA2        o099(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n122_), .B(ori_ori_n121_), .Y(ori_ori_n123_));
  NO2        o101(.A(ori_ori_n123_), .B(ori_ori_n46_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n90_), .B(ori_ori_n89_), .Y(ori_ori_n125_));
  NAi21      o103(.An(i_3_), .B(i_8_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n126_), .B(ori_ori_n61_), .Y(ori_ori_n127_));
  NOi31      o105(.An(ori_ori_n127_), .B(ori_ori_n125_), .C(ori_ori_n124_), .Y(ori_ori_n128_));
  NO2        o106(.A(i_1_), .B(ori_ori_n85_), .Y(ori_ori_n129_));
  NO2        o107(.A(i_6_), .B(i_5_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n130_), .B(i_3_), .Y(ori_ori_n131_));
  AO210      o109(.A0(ori_ori_n131_), .A1(ori_ori_n47_), .B0(ori_ori_n129_), .Y(ori_ori_n132_));
  OAI220     o110(.A0(ori_ori_n132_), .A1(ori_ori_n107_), .B0(ori_ori_n128_), .B1(ori_ori_n120_), .Y(ori_ori_n133_));
  NO3        o111(.A(ori_ori_n133_), .B(ori_ori_n118_), .C(ori_ori_n94_), .Y(ori_ori_n134_));
  NA3        o112(.A(ori_ori_n134_), .B(ori_ori_n78_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o113(.A(ori_ori_n62_), .B(ori_ori_n37_), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n646_), .B(ori_ori_n136_), .Y(ori_ori_n137_));
  NA4        o115(.A(ori_ori_n137_), .B(ori_ori_n76_), .C(ori_ori_n68_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o116(.A(i_8_), .B(i_7_), .Y(ori_ori_n139_));
  NA2        o117(.A(ori_ori_n139_), .B(i_6_), .Y(ori_ori_n140_));
  NO2        o118(.A(i_12_), .B(i_13_), .Y(ori_ori_n141_));
  NAi21      o119(.An(i_5_), .B(i_11_), .Y(ori_ori_n142_));
  NO2        o120(.A(i_0_), .B(i_1_), .Y(ori_ori_n143_));
  NA2        o121(.A(i_2_), .B(i_3_), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n144_), .B(i_4_), .Y(ori_ori_n145_));
  AN2        o123(.A(ori_ori_n141_), .B(ori_ori_n82_), .Y(ori_ori_n146_));
  NA2        o124(.A(i_1_), .B(i_5_), .Y(ori_ori_n147_));
  OR2        o125(.A(i_0_), .B(i_1_), .Y(ori_ori_n148_));
  NO3        o126(.A(ori_ori_n148_), .B(ori_ori_n79_), .C(i_13_), .Y(ori_ori_n149_));
  NAi32      o127(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n150_));
  NAi21      o128(.An(ori_ori_n150_), .B(ori_ori_n149_), .Y(ori_ori_n151_));
  NOi21      o129(.An(i_4_), .B(i_10_), .Y(ori_ori_n152_));
  NA2        o130(.A(ori_ori_n152_), .B(ori_ori_n40_), .Y(ori_ori_n153_));
  NOi21      o131(.An(i_4_), .B(i_9_), .Y(ori_ori_n154_));
  NOi21      o132(.An(i_11_), .B(i_13_), .Y(ori_ori_n155_));
  NA2        o133(.A(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n72_), .B(ori_ori_n62_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n72_), .B(i_5_), .Y(ori_ori_n158_));
  NO2        o136(.A(i_2_), .B(i_1_), .Y(ori_ori_n159_));
  NAi21      o137(.An(i_4_), .B(i_12_), .Y(ori_ori_n160_));
  INV        o138(.A(i_8_), .Y(ori_ori_n161_));
  NO2        o139(.A(i_3_), .B(i_8_), .Y(ori_ori_n162_));
  NO3        o140(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n163_));
  NO2        o141(.A(ori_ori_n102_), .B(ori_ori_n57_), .Y(ori_ori_n164_));
  NO2        o142(.A(i_13_), .B(i_9_), .Y(ori_ori_n165_));
  NAi21      o143(.An(i_12_), .B(i_3_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n167_));
  NAi21      o145(.An(i_12_), .B(i_7_), .Y(ori_ori_n168_));
  NA3        o146(.A(i_13_), .B(ori_ori_n161_), .C(i_10_), .Y(ori_ori_n169_));
  NA2        o147(.A(i_0_), .B(i_5_), .Y(ori_ori_n170_));
  NAi31      o148(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n171_));
  INV        o149(.A(i_13_), .Y(ori_ori_n172_));
  NO2        o150(.A(i_12_), .B(ori_ori_n172_), .Y(ori_ori_n173_));
  NO2        o151(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n174_));
  OR2        o152(.A(i_8_), .B(i_7_), .Y(ori_ori_n175_));
  INV        o153(.A(i_12_), .Y(ori_ori_n176_));
  NO2        o154(.A(ori_ori_n44_), .B(ori_ori_n176_), .Y(ori_ori_n177_));
  NO3        o155(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n178_));
  NA2        o156(.A(i_2_), .B(i_1_), .Y(ori_ori_n179_));
  NO3        o157(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n180_));
  NAi21      o158(.An(i_4_), .B(i_3_), .Y(ori_ori_n181_));
  NO2        o159(.A(i_0_), .B(i_6_), .Y(ori_ori_n182_));
  NOi41      o160(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n183_));
  NO2        o161(.A(i_11_), .B(ori_ori_n172_), .Y(ori_ori_n184_));
  NOi21      o162(.An(i_1_), .B(i_6_), .Y(ori_ori_n185_));
  NAi21      o163(.An(i_3_), .B(i_7_), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n176_), .B(i_9_), .Y(ori_ori_n187_));
  OR4        o165(.A(ori_ori_n187_), .B(ori_ori_n186_), .C(ori_ori_n185_), .D(ori_ori_n158_), .Y(ori_ori_n188_));
  NA2        o166(.A(ori_ori_n72_), .B(i_5_), .Y(ori_ori_n189_));
  NA2        o167(.A(i_3_), .B(i_9_), .Y(ori_ori_n190_));
  NAi21      o168(.An(i_7_), .B(i_10_), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n191_), .B(ori_ori_n190_), .Y(ori_ori_n192_));
  NA3        o170(.A(ori_ori_n192_), .B(ori_ori_n189_), .C(ori_ori_n63_), .Y(ori_ori_n193_));
  NA2        o171(.A(ori_ori_n193_), .B(ori_ori_n188_), .Y(ori_ori_n194_));
  INV        o172(.A(ori_ori_n140_), .Y(ori_ori_n195_));
  NA2        o173(.A(ori_ori_n176_), .B(i_13_), .Y(ori_ori_n196_));
  NO2        o174(.A(ori_ori_n196_), .B(ori_ori_n74_), .Y(ori_ori_n197_));
  AOI220     o175(.A0(ori_ori_n197_), .A1(ori_ori_n195_), .B0(ori_ori_n194_), .B1(ori_ori_n184_), .Y(ori_ori_n198_));
  NA2        o176(.A(i_12_), .B(i_6_), .Y(ori_ori_n199_));
  OR2        o177(.A(i_13_), .B(i_9_), .Y(ori_ori_n200_));
  NO2        o178(.A(ori_ori_n181_), .B(i_2_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n184_), .B(i_9_), .Y(ori_ori_n202_));
  NO3        o180(.A(i_11_), .B(ori_ori_n172_), .C(ori_ori_n25_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n186_), .B(i_8_), .Y(ori_ori_n204_));
  NO3        o182(.A(i_12_), .B(ori_ori_n172_), .C(ori_ori_n37_), .Y(ori_ori_n205_));
  NO2        o183(.A(i_2_), .B(ori_ori_n100_), .Y(ori_ori_n206_));
  AN2        o184(.A(i_3_), .B(i_10_), .Y(ori_ori_n207_));
  NO2        o185(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n208_));
  NO2        o186(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n209_));
  NO3        o187(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n210_));
  NO2        o188(.A(i_2_), .B(i_3_), .Y(ori_ori_n211_));
  OR2        o189(.A(i_0_), .B(i_5_), .Y(ori_ori_n212_));
  NO2        o190(.A(i_12_), .B(i_10_), .Y(ori_ori_n213_));
  NOi21      o191(.An(i_5_), .B(i_0_), .Y(ori_ori_n214_));
  NO2        o192(.A(i_1_), .B(i_7_), .Y(ori_ori_n215_));
  NOi21      o193(.An(ori_ori_n147_), .B(ori_ori_n103_), .Y(ori_ori_n216_));
  NO2        o194(.A(ori_ori_n216_), .B(ori_ori_n122_), .Y(ori_ori_n217_));
  NA2        o195(.A(ori_ori_n217_), .B(i_3_), .Y(ori_ori_n218_));
  NO2        o196(.A(ori_ori_n161_), .B(i_9_), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n219_), .B(ori_ori_n164_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n220_), .B(ori_ori_n46_), .Y(ori_ori_n221_));
  INV        o199(.A(ori_ori_n221_), .Y(ori_ori_n222_));
  AOI210     o200(.A0(ori_ori_n222_), .A1(ori_ori_n218_), .B0(ori_ori_n153_), .Y(ori_ori_n223_));
  INV        o201(.A(ori_ori_n223_), .Y(ori_ori_n224_));
  NOi32      o202(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n225_));
  INV        o203(.A(ori_ori_n225_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n150_), .B(ori_ori_n148_), .Y(ori_ori_n227_));
  NOi32      o205(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n228_));
  NAi21      o206(.An(i_6_), .B(i_1_), .Y(ori_ori_n229_));
  NO2        o207(.A(i_1_), .B(ori_ori_n100_), .Y(ori_ori_n230_));
  NAi21      o208(.An(i_3_), .B(i_4_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n231_), .B(i_9_), .Y(ori_ori_n232_));
  AN2        o210(.A(i_6_), .B(i_7_), .Y(ori_ori_n233_));
  OAI210     o211(.A0(ori_ori_n233_), .A1(ori_ori_n230_), .B0(ori_ori_n232_), .Y(ori_ori_n234_));
  NA2        o212(.A(i_2_), .B(i_7_), .Y(ori_ori_n235_));
  NO2        o213(.A(ori_ori_n231_), .B(i_10_), .Y(ori_ori_n236_));
  NA3        o214(.A(ori_ori_n236_), .B(ori_ori_n235_), .C(ori_ori_n182_), .Y(ori_ori_n237_));
  AOI210     o215(.A0(ori_ori_n237_), .A1(ori_ori_n234_), .B0(ori_ori_n158_), .Y(ori_ori_n238_));
  AOI210     o216(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n239_));
  OAI210     o217(.A0(ori_ori_n239_), .A1(ori_ori_n159_), .B0(ori_ori_n236_), .Y(ori_ori_n240_));
  AOI220     o218(.A0(ori_ori_n236_), .A1(ori_ori_n215_), .B0(ori_ori_n178_), .B1(ori_ori_n159_), .Y(ori_ori_n241_));
  AOI210     o219(.A0(ori_ori_n241_), .A1(ori_ori_n240_), .B0(i_5_), .Y(ori_ori_n242_));
  NO3        o220(.A(ori_ori_n242_), .B(ori_ori_n238_), .C(ori_ori_n227_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n243_), .B(ori_ori_n226_), .Y(ori_ori_n244_));
  AN2        o222(.A(i_12_), .B(i_5_), .Y(ori_ori_n245_));
  NO2        o223(.A(i_11_), .B(i_6_), .Y(ori_ori_n246_));
  NO2        o224(.A(i_5_), .B(i_10_), .Y(ori_ori_n247_));
  NO2        o225(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n248_));
  NO3        o226(.A(ori_ori_n85_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n249_));
  NO2        o227(.A(i_11_), .B(i_12_), .Y(ori_ori_n250_));
  NAi21      o228(.An(i_13_), .B(i_0_), .Y(ori_ori_n251_));
  NO3        o229(.A(i_1_), .B(i_12_), .C(ori_ori_n85_), .Y(ori_ori_n252_));
  NO2        o230(.A(i_0_), .B(i_11_), .Y(ori_ori_n253_));
  AN2        o231(.A(i_1_), .B(i_6_), .Y(ori_ori_n254_));
  NOi21      o232(.An(i_2_), .B(i_12_), .Y(ori_ori_n255_));
  NAi21      o233(.An(i_9_), .B(i_4_), .Y(ori_ori_n256_));
  OR2        o234(.A(i_13_), .B(i_10_), .Y(ori_ori_n257_));
  NO3        o235(.A(ori_ori_n257_), .B(ori_ori_n115_), .C(ori_ori_n256_), .Y(ori_ori_n258_));
  NO2        o236(.A(ori_ori_n156_), .B(ori_ori_n121_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n100_), .B(ori_ori_n25_), .Y(ori_ori_n260_));
  NA2        o238(.A(ori_ori_n205_), .B(ori_ori_n260_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n261_), .B(ori_ori_n216_), .Y(ori_ori_n262_));
  INV        o240(.A(ori_ori_n262_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n263_), .B(ori_ori_n26_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n161_), .B(i_10_), .Y(ori_ori_n265_));
  NA3        o243(.A(ori_ori_n189_), .B(ori_ori_n63_), .C(i_2_), .Y(ori_ori_n266_));
  NO2        o244(.A(ori_ori_n266_), .B(ori_ori_n265_), .Y(ori_ori_n267_));
  INV        o245(.A(ori_ori_n267_), .Y(ori_ori_n268_));
  NO2        o246(.A(ori_ori_n268_), .B(ori_ori_n202_), .Y(ori_ori_n269_));
  NO3        o247(.A(ori_ori_n269_), .B(ori_ori_n264_), .C(ori_ori_n244_), .Y(ori_ori_n270_));
  NO2        o248(.A(ori_ori_n72_), .B(i_13_), .Y(ori_ori_n271_));
  NO2        o249(.A(i_10_), .B(i_9_), .Y(ori_ori_n272_));
  NAi21      o250(.An(i_12_), .B(i_8_), .Y(ori_ori_n273_));
  NO2        o251(.A(ori_ori_n273_), .B(i_3_), .Y(ori_ori_n274_));
  NO3        o252(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n275_));
  NA2        o253(.A(ori_ori_n199_), .B(ori_ori_n96_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n276_), .B(ori_ori_n275_), .Y(ori_ori_n277_));
  NA2        o255(.A(i_8_), .B(i_9_), .Y(ori_ori_n278_));
  AOI210     o256(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n279_));
  OR2        o257(.A(ori_ori_n279_), .B(ori_ori_n278_), .Y(ori_ori_n280_));
  NA2        o258(.A(ori_ori_n205_), .B(ori_ori_n164_), .Y(ori_ori_n281_));
  NO2        o259(.A(ori_ori_n281_), .B(ori_ori_n280_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n184_), .B(ori_ori_n208_), .Y(ori_ori_n283_));
  NO3        o261(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n284_));
  INV        o262(.A(ori_ori_n284_), .Y(ori_ori_n285_));
  NA3        o263(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n286_));
  NA4        o264(.A(ori_ori_n142_), .B(ori_ori_n114_), .C(ori_ori_n79_), .D(ori_ori_n23_), .Y(ori_ori_n287_));
  OAI220     o265(.A0(ori_ori_n287_), .A1(ori_ori_n286_), .B0(ori_ori_n285_), .B1(ori_ori_n283_), .Y(ori_ori_n288_));
  NO2        o266(.A(ori_ori_n288_), .B(ori_ori_n282_), .Y(ori_ori_n289_));
  NA2        o267(.A(ori_ori_n95_), .B(i_13_), .Y(ori_ori_n290_));
  NO2        o268(.A(i_11_), .B(i_1_), .Y(ori_ori_n291_));
  NOi21      o269(.An(i_2_), .B(i_7_), .Y(ori_ori_n292_));
  NO2        o270(.A(i_6_), .B(i_10_), .Y(ori_ori_n293_));
  NA3        o271(.A(ori_ori_n183_), .B(ori_ori_n155_), .C(ori_ori_n130_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n295_));
  NO2        o273(.A(ori_ori_n148_), .B(i_3_), .Y(ori_ori_n296_));
  NAi31      o274(.An(ori_ori_n295_), .B(ori_ori_n296_), .C(ori_ori_n173_), .Y(ori_ori_n297_));
  NA3        o275(.A(ori_ori_n248_), .B(ori_ori_n157_), .C(ori_ori_n145_), .Y(ori_ori_n298_));
  NA3        o276(.A(ori_ori_n298_), .B(ori_ori_n297_), .C(ori_ori_n294_), .Y(ori_ori_n299_));
  INV        o277(.A(ori_ori_n299_), .Y(ori_ori_n300_));
  NA2        o278(.A(ori_ori_n275_), .B(ori_ori_n245_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n284_), .B(ori_ori_n247_), .Y(ori_ori_n302_));
  NAi21      o280(.An(ori_ori_n169_), .B(ori_ori_n250_), .Y(ori_ori_n303_));
  NA2        o281(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n304_));
  NA2        o282(.A(ori_ori_n210_), .B(ori_ori_n178_), .Y(ori_ori_n305_));
  OAI220     o283(.A0(ori_ori_n305_), .A1(ori_ori_n266_), .B0(ori_ori_n304_), .B1(ori_ori_n290_), .Y(ori_ori_n306_));
  INV        o284(.A(ori_ori_n306_), .Y(ori_ori_n307_));
  NA3        o285(.A(ori_ori_n307_), .B(ori_ori_n300_), .C(ori_ori_n289_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n245_), .B(ori_ori_n172_), .Y(ori_ori_n309_));
  NA2        o287(.A(ori_ori_n233_), .B(ori_ori_n228_), .Y(ori_ori_n310_));
  OR2        o288(.A(ori_ori_n309_), .B(ori_ori_n310_), .Y(ori_ori_n311_));
  NO2        o289(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n312_));
  AOI210     o290(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n258_), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n313_), .B(ori_ori_n311_), .Y(ori_ori_n314_));
  INV        o292(.A(ori_ori_n314_), .Y(ori_ori_n315_));
  INV        o293(.A(ori_ori_n132_), .Y(ori_ori_n316_));
  NA2        o294(.A(ori_ori_n316_), .B(ori_ori_n259_), .Y(ori_ori_n317_));
  NA2        o295(.A(ori_ori_n317_), .B(ori_ori_n315_), .Y(ori_ori_n318_));
  NO2        o296(.A(i_12_), .B(ori_ori_n161_), .Y(ori_ori_n319_));
  NA2        o297(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n320_));
  NO2        o298(.A(ori_ori_n320_), .B(i_6_), .Y(ori_ori_n321_));
  NO2        o299(.A(ori_ori_n148_), .B(i_5_), .Y(ori_ori_n322_));
  NA3        o300(.A(ori_ori_n170_), .B(ori_ori_n70_), .C(ori_ori_n44_), .Y(ori_ori_n323_));
  NA2        o301(.A(ori_ori_n205_), .B(ori_ori_n83_), .Y(ori_ori_n324_));
  NO2        o302(.A(ori_ori_n323_), .B(ori_ori_n324_), .Y(ori_ori_n325_));
  AOI210     o303(.A0(ori_ori_n229_), .A1(ori_ori_n46_), .B0(ori_ori_n230_), .Y(ori_ori_n326_));
  NA2        o304(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n327_));
  NA3        o305(.A(ori_ori_n319_), .B(ori_ori_n203_), .C(ori_ori_n327_), .Y(ori_ori_n328_));
  NO2        o306(.A(ori_ori_n326_), .B(ori_ori_n328_), .Y(ori_ori_n329_));
  NO2        o307(.A(ori_ori_n329_), .B(ori_ori_n325_), .Y(ori_ori_n330_));
  NO3        o308(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n331_));
  NO2        o309(.A(ori_ori_n257_), .B(i_1_), .Y(ori_ori_n332_));
  NOi31      o310(.An(ori_ori_n332_), .B(ori_ori_n276_), .C(ori_ori_n72_), .Y(ori_ori_n333_));
  NOi21      o311(.An(i_10_), .B(i_6_), .Y(ori_ori_n334_));
  NO2        o312(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n113_), .B(ori_ori_n23_), .Y(ori_ori_n336_));
  NO2        o314(.A(i_12_), .B(ori_ori_n85_), .Y(ori_ori_n337_));
  OR2        o315(.A(i_2_), .B(i_5_), .Y(ori_ori_n338_));
  OR2        o316(.A(ori_ori_n338_), .B(ori_ori_n254_), .Y(ori_ori_n339_));
  NA2        o317(.A(ori_ori_n235_), .B(ori_ori_n182_), .Y(ori_ori_n340_));
  AOI210     o318(.A0(ori_ori_n340_), .A1(ori_ori_n339_), .B0(ori_ori_n303_), .Y(ori_ori_n341_));
  INV        o319(.A(ori_ori_n341_), .Y(ori_ori_n342_));
  NA2        o320(.A(ori_ori_n342_), .B(ori_ori_n330_), .Y(ori_ori_n343_));
  NO3        o321(.A(ori_ori_n343_), .B(ori_ori_n318_), .C(ori_ori_n308_), .Y(ori_ori_n344_));
  NA4        o322(.A(ori_ori_n344_), .B(ori_ori_n270_), .C(ori_ori_n224_), .D(ori_ori_n198_), .Y(ori7));
  NO2        o323(.A(ori_ori_n92_), .B(ori_ori_n54_), .Y(ori_ori_n346_));
  NA2        o324(.A(ori_ori_n293_), .B(ori_ori_n83_), .Y(ori_ori_n347_));
  NA2        o325(.A(i_11_), .B(ori_ori_n161_), .Y(ori_ori_n348_));
  NA2        o326(.A(ori_ori_n141_), .B(ori_ori_n348_), .Y(ori_ori_n349_));
  NO2        o327(.A(ori_ori_n349_), .B(ori_ori_n347_), .Y(ori_ori_n350_));
  NA3        o328(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n351_));
  NO2        o329(.A(ori_ori_n176_), .B(i_4_), .Y(ori_ori_n352_));
  NA2        o330(.A(ori_ori_n352_), .B(i_8_), .Y(ori_ori_n353_));
  NO2        o331(.A(ori_ori_n104_), .B(ori_ori_n351_), .Y(ori_ori_n354_));
  NA2        o332(.A(i_2_), .B(ori_ori_n85_), .Y(ori_ori_n355_));
  OAI210     o333(.A0(ori_ori_n86_), .A1(ori_ori_n162_), .B0(ori_ori_n163_), .Y(ori_ori_n356_));
  NO2        o334(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n357_));
  NA2        o335(.A(i_4_), .B(i_8_), .Y(ori_ori_n358_));
  AOI210     o336(.A0(ori_ori_n358_), .A1(ori_ori_n207_), .B0(ori_ori_n357_), .Y(ori_ori_n359_));
  OAI220     o337(.A0(ori_ori_n359_), .A1(ori_ori_n355_), .B0(ori_ori_n356_), .B1(i_13_), .Y(ori_ori_n360_));
  NO4        o338(.A(ori_ori_n360_), .B(ori_ori_n354_), .C(ori_ori_n350_), .D(ori_ori_n346_), .Y(ori_ori_n361_));
  AOI210     o339(.A0(ori_ori_n126_), .A1(ori_ori_n61_), .B0(i_10_), .Y(ori_ori_n362_));
  AOI210     o340(.A0(ori_ori_n362_), .A1(ori_ori_n176_), .B0(ori_ori_n152_), .Y(ori_ori_n363_));
  OR2        o341(.A(i_6_), .B(i_10_), .Y(ori_ori_n364_));
  OR3        o342(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n365_));
  OR2        o343(.A(ori_ori_n363_), .B(ori_ori_n200_), .Y(ori_ori_n366_));
  AOI210     o344(.A0(ori_ori_n366_), .A1(ori_ori_n361_), .B0(ori_ori_n62_), .Y(ori_ori_n367_));
  NOi21      o345(.An(i_11_), .B(i_7_), .Y(ori_ori_n368_));
  AO210      o346(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n369_));
  NO2        o347(.A(ori_ori_n369_), .B(ori_ori_n368_), .Y(ori_ori_n370_));
  NA2        o348(.A(ori_ori_n370_), .B(ori_ori_n165_), .Y(ori_ori_n371_));
  NA3        o349(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n372_));
  NO2        o350(.A(ori_ori_n371_), .B(ori_ori_n62_), .Y(ori_ori_n373_));
  OR2        o351(.A(ori_ori_n241_), .B(ori_ori_n41_), .Y(ori_ori_n374_));
  NA2        o352(.A(ori_ori_n173_), .B(ori_ori_n62_), .Y(ori_ori_n375_));
  OR2        o353(.A(ori_ori_n166_), .B(ori_ori_n107_), .Y(ori_ori_n376_));
  NO2        o354(.A(i_1_), .B(i_12_), .Y(ori_ori_n377_));
  NA2        o355(.A(ori_ori_n375_), .B(ori_ori_n374_), .Y(ori_ori_n378_));
  OAI210     o356(.A0(ori_ori_n378_), .A1(ori_ori_n373_), .B0(i_6_), .Y(ori_ori_n379_));
  NO2        o357(.A(ori_ori_n372_), .B(ori_ori_n107_), .Y(ori_ori_n380_));
  NA2        o358(.A(ori_ori_n380_), .B(ori_ori_n337_), .Y(ori_ori_n381_));
  NO2        o359(.A(i_6_), .B(i_11_), .Y(ori_ori_n382_));
  NA2        o360(.A(ori_ori_n381_), .B(ori_ori_n277_), .Y(ori_ori_n383_));
  NO3        o361(.A(ori_ori_n364_), .B(ori_ori_n175_), .C(ori_ori_n23_), .Y(ori_ori_n384_));
  AOI210     o362(.A0(i_1_), .A1(ori_ori_n192_), .B0(ori_ori_n384_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n385_), .B(ori_ori_n44_), .Y(ori_ori_n386_));
  INV        o364(.A(i_2_), .Y(ori_ori_n387_));
  NA2        o365(.A(ori_ori_n136_), .B(i_9_), .Y(ori_ori_n388_));
  NO2        o366(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n389_));
  NO2        o367(.A(ori_ori_n388_), .B(ori_ori_n387_), .Y(ori_ori_n390_));
  AOI210     o368(.A0(ori_ori_n291_), .A1(ori_ori_n260_), .B0(ori_ori_n180_), .Y(ori_ori_n391_));
  NO2        o369(.A(ori_ori_n391_), .B(ori_ori_n355_), .Y(ori_ori_n392_));
  NO2        o370(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n393_));
  OR2        o371(.A(ori_ori_n392_), .B(ori_ori_n390_), .Y(ori_ori_n394_));
  NO3        o372(.A(ori_ori_n394_), .B(ori_ori_n386_), .C(ori_ori_n383_), .Y(ori_ori_n395_));
  NO2        o373(.A(ori_ori_n176_), .B(ori_ori_n100_), .Y(ori_ori_n396_));
  NO2        o374(.A(ori_ori_n396_), .B(ori_ori_n368_), .Y(ori_ori_n397_));
  NA2        o375(.A(ori_ori_n397_), .B(i_1_), .Y(ori_ori_n398_));
  NO2        o376(.A(ori_ori_n398_), .B(ori_ori_n365_), .Y(ori_ori_n399_));
  NO2        o377(.A(ori_ori_n256_), .B(ori_ori_n85_), .Y(ori_ori_n400_));
  NA2        o378(.A(ori_ori_n399_), .B(ori_ori_n46_), .Y(ori_ori_n401_));
  NA2        o379(.A(i_3_), .B(ori_ori_n161_), .Y(ori_ori_n402_));
  NO2        o380(.A(ori_ori_n402_), .B(ori_ori_n113_), .Y(ori_ori_n403_));
  AN2        o381(.A(ori_ori_n403_), .B(ori_ori_n321_), .Y(ori_ori_n404_));
  NO2        o382(.A(ori_ori_n175_), .B(ori_ori_n44_), .Y(ori_ori_n405_));
  NO3        o383(.A(ori_ori_n405_), .B(ori_ori_n209_), .C(ori_ori_n177_), .Y(ori_ori_n406_));
  NO2        o384(.A(ori_ori_n115_), .B(ori_ori_n37_), .Y(ori_ori_n407_));
  NO2        o385(.A(ori_ori_n407_), .B(i_6_), .Y(ori_ori_n408_));
  NO2        o386(.A(ori_ori_n85_), .B(i_9_), .Y(ori_ori_n409_));
  NO2        o387(.A(ori_ori_n409_), .B(ori_ori_n62_), .Y(ori_ori_n410_));
  NO2        o388(.A(ori_ori_n410_), .B(ori_ori_n377_), .Y(ori_ori_n411_));
  NO4        o389(.A(ori_ori_n411_), .B(ori_ori_n408_), .C(ori_ori_n406_), .D(i_4_), .Y(ori_ori_n412_));
  NA2        o390(.A(i_1_), .B(i_3_), .Y(ori_ori_n413_));
  NO2        o391(.A(ori_ori_n278_), .B(ori_ori_n92_), .Y(ori_ori_n414_));
  AOI210     o392(.A0(ori_ori_n405_), .A1(ori_ori_n334_), .B0(ori_ori_n414_), .Y(ori_ori_n415_));
  NO2        o393(.A(ori_ori_n415_), .B(ori_ori_n413_), .Y(ori_ori_n416_));
  NO3        o394(.A(ori_ori_n416_), .B(ori_ori_n412_), .C(ori_ori_n404_), .Y(ori_ori_n417_));
  NA4        o395(.A(ori_ori_n417_), .B(ori_ori_n401_), .C(ori_ori_n395_), .D(ori_ori_n379_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n233_), .B(ori_ori_n232_), .Y(ori_ori_n419_));
  INV        o397(.A(ori_ori_n419_), .Y(ori_ori_n420_));
  NA2        o398(.A(ori_ori_n420_), .B(i_1_), .Y(ori_ori_n421_));
  AOI210     o399(.A0(ori_ori_n199_), .A1(ori_ori_n96_), .B0(i_1_), .Y(ori_ori_n422_));
  NO2        o400(.A(ori_ori_n231_), .B(i_2_), .Y(ori_ori_n423_));
  NA2        o401(.A(ori_ori_n423_), .B(ori_ori_n422_), .Y(ori_ori_n424_));
  AOI210     o402(.A0(ori_ori_n424_), .A1(ori_ori_n421_), .B0(i_13_), .Y(ori_ori_n425_));
  OR2        o403(.A(i_11_), .B(i_7_), .Y(ori_ori_n426_));
  NO2        o404(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n427_));
  NO2        o405(.A(ori_ori_n292_), .B(ori_ori_n24_), .Y(ori_ori_n428_));
  NA2        o406(.A(ori_ori_n428_), .B(ori_ori_n400_), .Y(ori_ori_n429_));
  OAI220     o407(.A0(ori_ori_n429_), .A1(ori_ori_n41_), .B0(ori_ori_n645_), .B1(ori_ori_n92_), .Y(ori_ori_n430_));
  INV        o408(.A(ori_ori_n430_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n246_), .B(ori_ori_n389_), .Y(ori_ori_n432_));
  NO2        o410(.A(ori_ori_n432_), .B(ori_ori_n181_), .Y(ori_ori_n433_));
  AOI210     o411(.A0(ori_ori_n273_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n434_));
  NOi31      o412(.An(ori_ori_n434_), .B(ori_ori_n347_), .C(ori_ori_n44_), .Y(ori_ori_n435_));
  NA2        o413(.A(ori_ori_n125_), .B(i_13_), .Y(ori_ori_n436_));
  NO2        o414(.A(ori_ori_n436_), .B(ori_ori_n422_), .Y(ori_ori_n437_));
  NA2        o415(.A(ori_ori_n26_), .B(ori_ori_n161_), .Y(ori_ori_n438_));
  NA2        o416(.A(ori_ori_n438_), .B(i_7_), .Y(ori_ori_n439_));
  AOI220     o417(.A0(ori_ori_n246_), .A1(ori_ori_n389_), .B0(ori_ori_n91_), .B1(ori_ori_n101_), .Y(ori_ori_n440_));
  NO2        o418(.A(ori_ori_n440_), .B(ori_ori_n353_), .Y(ori_ori_n441_));
  NO4        o419(.A(ori_ori_n441_), .B(ori_ori_n437_), .C(ori_ori_n435_), .D(ori_ori_n433_), .Y(ori_ori_n442_));
  OR2        o420(.A(i_11_), .B(i_6_), .Y(ori_ori_n443_));
  NA3        o421(.A(ori_ori_n352_), .B(ori_ori_n438_), .C(i_7_), .Y(ori_ori_n444_));
  NO2        o422(.A(ori_ori_n444_), .B(ori_ori_n443_), .Y(ori_ori_n445_));
  NA3        o423(.A(ori_ori_n255_), .B(ori_ori_n357_), .C(ori_ori_n96_), .Y(ori_ori_n446_));
  NA2        o424(.A(ori_ori_n382_), .B(i_13_), .Y(ori_ori_n447_));
  NAi21      o425(.An(i_11_), .B(i_12_), .Y(ori_ori_n448_));
  NOi41      o426(.An(ori_ori_n109_), .B(ori_ori_n448_), .C(i_13_), .D(ori_ori_n85_), .Y(ori_ori_n449_));
  NA2        o427(.A(ori_ori_n449_), .B(ori_ori_n46_), .Y(ori_ori_n450_));
  NA3        o428(.A(ori_ori_n450_), .B(ori_ori_n447_), .C(ori_ori_n446_), .Y(ori_ori_n451_));
  OAI210     o429(.A0(ori_ori_n451_), .A1(ori_ori_n445_), .B0(ori_ori_n62_), .Y(ori_ori_n452_));
  NO2        o430(.A(i_2_), .B(i_12_), .Y(ori_ori_n453_));
  NA2        o431(.A(ori_ori_n230_), .B(ori_ori_n453_), .Y(ori_ori_n454_));
  NA2        o432(.A(ori_ori_n232_), .B(ori_ori_n230_), .Y(ori_ori_n455_));
  NA2        o433(.A(ori_ori_n455_), .B(ori_ori_n454_), .Y(ori_ori_n456_));
  NA3        o434(.A(ori_ori_n456_), .B(ori_ori_n45_), .C(ori_ori_n172_), .Y(ori_ori_n457_));
  NA4        o435(.A(ori_ori_n457_), .B(ori_ori_n452_), .C(ori_ori_n442_), .D(ori_ori_n431_), .Y(ori_ori_n458_));
  OR4        o436(.A(ori_ori_n458_), .B(ori_ori_n425_), .C(ori_ori_n418_), .D(ori_ori_n367_), .Y(ori5));
  NA2        o437(.A(ori_ori_n397_), .B(ori_ori_n201_), .Y(ori_ori_n460_));
  AN2        o438(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n461_));
  NA3        o439(.A(ori_ori_n461_), .B(ori_ori_n453_), .C(ori_ori_n107_), .Y(ori_ori_n462_));
  NO2        o440(.A(ori_ori_n353_), .B(i_11_), .Y(ori_ori_n463_));
  NA2        o441(.A(ori_ori_n86_), .B(ori_ori_n463_), .Y(ori_ori_n464_));
  NA3        o442(.A(ori_ori_n464_), .B(ori_ori_n462_), .C(ori_ori_n460_), .Y(ori_ori_n465_));
  NO3        o443(.A(i_11_), .B(ori_ori_n176_), .C(i_13_), .Y(ori_ori_n466_));
  NO2        o444(.A(ori_ori_n122_), .B(ori_ori_n23_), .Y(ori_ori_n467_));
  NA2        o445(.A(i_12_), .B(i_8_), .Y(ori_ori_n468_));
  OAI210     o446(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n468_), .Y(ori_ori_n469_));
  INV        o447(.A(ori_ori_n272_), .Y(ori_ori_n470_));
  AOI220     o448(.A0(ori_ori_n211_), .A1(ori_ori_n336_), .B0(ori_ori_n469_), .B1(ori_ori_n467_), .Y(ori_ori_n471_));
  INV        o449(.A(ori_ori_n471_), .Y(ori_ori_n472_));
  NO2        o450(.A(ori_ori_n472_), .B(ori_ori_n465_), .Y(ori_ori_n473_));
  INV        o451(.A(ori_ori_n155_), .Y(ori_ori_n474_));
  INV        o452(.A(ori_ori_n183_), .Y(ori_ori_n475_));
  OAI210     o453(.A0(ori_ori_n423_), .A1(ori_ori_n274_), .B0(ori_ori_n109_), .Y(ori_ori_n476_));
  AOI210     o454(.A0(ori_ori_n476_), .A1(ori_ori_n475_), .B0(ori_ori_n474_), .Y(ori_ori_n477_));
  NO2        o455(.A(ori_ori_n278_), .B(ori_ori_n26_), .Y(ori_ori_n478_));
  NO2        o456(.A(ori_ori_n478_), .B(ori_ori_n260_), .Y(ori_ori_n479_));
  NA2        o457(.A(ori_ori_n479_), .B(i_2_), .Y(ori_ori_n480_));
  INV        o458(.A(ori_ori_n480_), .Y(ori_ori_n481_));
  AOI210     o459(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n257_), .Y(ori_ori_n482_));
  AOI210     o460(.A0(ori_ori_n482_), .A1(ori_ori_n481_), .B0(ori_ori_n477_), .Y(ori_ori_n483_));
  NO2        o461(.A(ori_ori_n160_), .B(ori_ori_n123_), .Y(ori_ori_n484_));
  OAI210     o462(.A0(ori_ori_n484_), .A1(ori_ori_n467_), .B0(i_2_), .Y(ori_ori_n485_));
  INV        o463(.A(ori_ori_n156_), .Y(ori_ori_n486_));
  NO3        o464(.A(ori_ori_n369_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n487_));
  AOI210     o465(.A0(ori_ori_n486_), .A1(ori_ori_n86_), .B0(ori_ori_n487_), .Y(ori_ori_n488_));
  AOI210     o466(.A0(ori_ori_n488_), .A1(ori_ori_n485_), .B0(ori_ori_n161_), .Y(ori_ori_n489_));
  OA210      o467(.A0(ori_ori_n370_), .A1(ori_ori_n124_), .B0(i_13_), .Y(ori_ori_n490_));
  NA2        o468(.A(ori_ori_n146_), .B(ori_ori_n348_), .Y(ori_ori_n491_));
  NO2        o469(.A(ori_ori_n491_), .B(ori_ori_n235_), .Y(ori_ori_n492_));
  AOI210     o470(.A0(ori_ori_n166_), .A1(ori_ori_n144_), .B0(ori_ori_n312_), .Y(ori_ori_n493_));
  NA2        o471(.A(ori_ori_n493_), .B(ori_ori_n260_), .Y(ori_ori_n494_));
  NO2        o472(.A(ori_ori_n101_), .B(ori_ori_n44_), .Y(ori_ori_n495_));
  INV        o473(.A(ori_ori_n206_), .Y(ori_ori_n496_));
  NA4        o474(.A(ori_ori_n496_), .B(ori_ori_n207_), .C(ori_ori_n122_), .D(ori_ori_n42_), .Y(ori_ori_n497_));
  OAI210     o475(.A0(ori_ori_n497_), .A1(ori_ori_n495_), .B0(ori_ori_n494_), .Y(ori_ori_n498_));
  NO4        o476(.A(ori_ori_n498_), .B(ori_ori_n492_), .C(ori_ori_n490_), .D(ori_ori_n489_), .Y(ori_ori_n499_));
  NA2        o477(.A(ori_ori_n336_), .B(ori_ori_n28_), .Y(ori_ori_n500_));
  NA2        o478(.A(ori_ori_n466_), .B(ori_ori_n204_), .Y(ori_ori_n501_));
  NA2        o479(.A(ori_ori_n501_), .B(ori_ori_n500_), .Y(ori_ori_n502_));
  NO2        o480(.A(ori_ori_n61_), .B(i_12_), .Y(ori_ori_n503_));
  NO2        o481(.A(ori_ori_n503_), .B(ori_ori_n124_), .Y(ori_ori_n504_));
  NO2        o482(.A(ori_ori_n504_), .B(ori_ori_n348_), .Y(ori_ori_n505_));
  AOI220     o483(.A0(ori_ori_n505_), .A1(ori_ori_n36_), .B0(ori_ori_n502_), .B1(ori_ori_n46_), .Y(ori_ori_n506_));
  NA4        o484(.A(ori_ori_n506_), .B(ori_ori_n499_), .C(ori_ori_n483_), .D(ori_ori_n473_), .Y(ori6));
  NO2        o485(.A(ori_ori_n171_), .B(ori_ori_n295_), .Y(ori_ori_n508_));
  OR2        o486(.A(ori_ori_n647_), .B(i_12_), .Y(ori_ori_n509_));
  NA2        o487(.A(ori_ori_n337_), .B(ori_ori_n62_), .Y(ori_ori_n510_));
  INV        o488(.A(ori_ori_n510_), .Y(ori_ori_n511_));
  NA2        o489(.A(ori_ori_n511_), .B(ori_ori_n72_), .Y(ori_ori_n512_));
  INV        o490(.A(ori_ori_n213_), .Y(ori_ori_n513_));
  NA2        o491(.A(ori_ori_n74_), .B(ori_ori_n129_), .Y(ori_ori_n514_));
  INV        o492(.A(ori_ori_n122_), .Y(ori_ori_n515_));
  NA2        o493(.A(ori_ori_n515_), .B(ori_ori_n46_), .Y(ori_ori_n516_));
  AOI210     o494(.A0(ori_ori_n516_), .A1(ori_ori_n514_), .B0(ori_ori_n513_), .Y(ori_ori_n517_));
  NO2        o495(.A(ori_ori_n185_), .B(i_9_), .Y(ori_ori_n518_));
  NA2        o496(.A(ori_ori_n518_), .B(ori_ori_n503_), .Y(ori_ori_n519_));
  AOI210     o497(.A0(ori_ori_n519_), .A1(ori_ori_n310_), .B0(ori_ori_n158_), .Y(ori_ori_n520_));
  NAi32      o498(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n521_));
  NO2        o499(.A(ori_ori_n443_), .B(ori_ori_n521_), .Y(ori_ori_n522_));
  OR3        o500(.A(ori_ori_n522_), .B(ori_ori_n520_), .C(ori_ori_n517_), .Y(ori_ori_n523_));
  NO2        o501(.A(ori_ori_n426_), .B(i_2_), .Y(ori_ori_n524_));
  BUFFER     o502(.A(ori_ori_n370_), .Y(ori_ori_n525_));
  NA3        o503(.A(ori_ori_n525_), .B(ori_ori_n143_), .C(ori_ori_n68_), .Y(ori_ori_n526_));
  AO210      o504(.A0(ori_ori_n302_), .A1(ori_ori_n470_), .B0(ori_ori_n36_), .Y(ori_ori_n527_));
  NA2        o505(.A(ori_ori_n527_), .B(ori_ori_n526_), .Y(ori_ori_n528_));
  NO2        o506(.A(i_6_), .B(i_11_), .Y(ori_ori_n529_));
  AOI220     o507(.A0(ori_ori_n529_), .A1(ori_ori_n331_), .B0(ori_ori_n508_), .B1(ori_ori_n439_), .Y(ori_ori_n530_));
  NA3        o508(.A(ori_ori_n235_), .B(ori_ori_n178_), .C(ori_ori_n143_), .Y(ori_ori_n531_));
  NA2        o509(.A(ori_ori_n249_), .B(ori_ori_n69_), .Y(ori_ori_n532_));
  NA4        o510(.A(ori_ori_n532_), .B(ori_ori_n531_), .C(ori_ori_n530_), .D(ori_ori_n356_), .Y(ori_ori_n533_));
  NA2        o511(.A(ori_ori_n274_), .B(ori_ori_n272_), .Y(ori_ori_n534_));
  NO2        o512(.A(ori_ori_n364_), .B(ori_ori_n101_), .Y(ori_ori_n535_));
  OAI210     o513(.A0(ori_ori_n535_), .A1(ori_ori_n110_), .B0(ori_ori_n253_), .Y(ori_ori_n536_));
  INV        o514(.A(ori_ori_n339_), .Y(ori_ori_n537_));
  NA3        o515(.A(ori_ori_n537_), .B(ori_ori_n213_), .C(i_7_), .Y(ori_ori_n538_));
  NA3        o516(.A(ori_ori_n538_), .B(ori_ori_n536_), .C(ori_ori_n534_), .Y(ori_ori_n539_));
  NO4        o517(.A(ori_ori_n539_), .B(ori_ori_n533_), .C(ori_ori_n528_), .D(ori_ori_n523_), .Y(ori_ori_n540_));
  NA4        o518(.A(ori_ori_n540_), .B(ori_ori_n512_), .C(ori_ori_n509_), .D(ori_ori_n243_), .Y(ori3));
  NA2        o519(.A(i_12_), .B(i_10_), .Y(ori_ori_n542_));
  NO2        o520(.A(i_11_), .B(ori_ori_n176_), .Y(ori_ori_n543_));
  NA3        o521(.A(ori_ori_n531_), .B(ori_ori_n356_), .C(ori_ori_n234_), .Y(ori_ori_n544_));
  NA2        o522(.A(ori_ori_n544_), .B(ori_ori_n40_), .Y(ori_ori_n545_));
  NOi21      o523(.An(ori_ori_n95_), .B(ori_ori_n479_), .Y(ori_ori_n546_));
  NO3        o524(.A(ori_ori_n376_), .B(ori_ori_n278_), .C(ori_ori_n129_), .Y(ori_ori_n547_));
  NA2        o525(.A(ori_ori_n255_), .B(ori_ori_n45_), .Y(ori_ori_n548_));
  AN2        o526(.A(ori_ori_n276_), .B(ori_ori_n55_), .Y(ori_ori_n549_));
  NO3        o527(.A(ori_ori_n549_), .B(ori_ori_n547_), .C(ori_ori_n546_), .Y(ori_ori_n550_));
  AOI210     o528(.A0(ori_ori_n550_), .A1(ori_ori_n545_), .B0(ori_ori_n48_), .Y(ori_ori_n551_));
  NO4        o529(.A(ori_ori_n239_), .B(ori_ori_n245_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n552_));
  NA2        o530(.A(ori_ori_n158_), .B(ori_ori_n334_), .Y(ori_ori_n553_));
  NOi21      o531(.An(ori_ori_n553_), .B(ori_ori_n552_), .Y(ori_ori_n554_));
  NO2        o532(.A(ori_ori_n554_), .B(ori_ori_n62_), .Y(ori_ori_n555_));
  NOi21      o533(.An(i_5_), .B(i_9_), .Y(ori_ori_n556_));
  NA2        o534(.A(ori_ori_n556_), .B(ori_ori_n271_), .Y(ori_ori_n557_));
  BUFFER     o535(.A(ori_ori_n199_), .Y(ori_ori_n558_));
  NA2        o536(.A(ori_ori_n558_), .B(ori_ori_n291_), .Y(ori_ori_n559_));
  NO2        o537(.A(ori_ori_n559_), .B(ori_ori_n557_), .Y(ori_ori_n560_));
  NO3        o538(.A(ori_ori_n560_), .B(ori_ori_n555_), .C(ori_ori_n551_), .Y(ori_ori_n561_));
  NA2        o539(.A(ori_ori_n335_), .B(i_0_), .Y(ori_ori_n562_));
  NO4        o540(.A(ori_ori_n338_), .B(ori_ori_n168_), .C(ori_ori_n257_), .D(ori_ori_n254_), .Y(ori_ori_n563_));
  NA2        o541(.A(ori_ori_n563_), .B(i_11_), .Y(ori_ori_n564_));
  NA2        o542(.A(ori_ori_n466_), .B(ori_ori_n214_), .Y(ori_ori_n565_));
  AOI210     o543(.A0(ori_ori_n293_), .A1(ori_ori_n86_), .B0(ori_ori_n57_), .Y(ori_ori_n566_));
  NO2        o544(.A(ori_ori_n566_), .B(ori_ori_n565_), .Y(ori_ori_n567_));
  NO2        o545(.A(ori_ori_n187_), .B(ori_ori_n147_), .Y(ori_ori_n568_));
  NA2        o546(.A(i_0_), .B(i_10_), .Y(ori_ori_n569_));
  INV        o547(.A(ori_ori_n320_), .Y(ori_ori_n570_));
  NO4        o548(.A(ori_ori_n113_), .B(ori_ori_n57_), .C(ori_ori_n402_), .D(i_5_), .Y(ori_ori_n571_));
  AO220      o549(.A0(ori_ori_n571_), .A1(ori_ori_n570_), .B0(ori_ori_n568_), .B1(i_6_), .Y(ori_ori_n572_));
  NO2        o550(.A(ori_ori_n572_), .B(ori_ori_n567_), .Y(ori_ori_n573_));
  NA2        o551(.A(ori_ori_n573_), .B(ori_ori_n564_), .Y(ori_ori_n574_));
  NO2        o552(.A(ori_ori_n102_), .B(ori_ori_n37_), .Y(ori_ori_n575_));
  NA2        o553(.A(i_11_), .B(i_9_), .Y(ori_ori_n576_));
  NO3        o554(.A(i_12_), .B(ori_ori_n576_), .C(ori_ori_n355_), .Y(ori_ori_n577_));
  AN2        o555(.A(ori_ori_n577_), .B(ori_ori_n575_), .Y(ori_ori_n578_));
  NA2        o556(.A(ori_ori_n248_), .B(ori_ori_n157_), .Y(ori_ori_n579_));
  NA2        o557(.A(ori_ori_n579_), .B(ori_ori_n151_), .Y(ori_ori_n580_));
  NO2        o558(.A(ori_ori_n576_), .B(ori_ori_n72_), .Y(ori_ori_n581_));
  INV        o559(.A(ori_ori_n252_), .Y(ori_ori_n582_));
  NO2        o560(.A(ori_ori_n582_), .B(ori_ori_n557_), .Y(ori_ori_n583_));
  NO3        o561(.A(ori_ori_n583_), .B(ori_ori_n580_), .C(ori_ori_n578_), .Y(ori_ori_n584_));
  NA2        o562(.A(ori_ori_n393_), .B(ori_ori_n119_), .Y(ori_ori_n585_));
  NO2        o563(.A(i_6_), .B(ori_ori_n585_), .Y(ori_ori_n586_));
  NA2        o564(.A(ori_ori_n155_), .B(ori_ori_n102_), .Y(ori_ori_n587_));
  INV        o565(.A(ori_ori_n586_), .Y(ori_ori_n588_));
  INV        o566(.A(ori_ori_n212_), .Y(ori_ori_n589_));
  NA2        o567(.A(ori_ori_n588_), .B(ori_ori_n584_), .Y(ori_ori_n590_));
  NO2        o568(.A(ori_ori_n542_), .B(ori_ori_n211_), .Y(ori_ori_n591_));
  NA2        o569(.A(ori_ori_n591_), .B(ori_ori_n581_), .Y(ori_ori_n592_));
  NA2        o570(.A(ori_ori_n428_), .B(ori_ori_n322_), .Y(ori_ori_n593_));
  NAi21      o571(.An(i_9_), .B(i_5_), .Y(ori_ori_n594_));
  NO2        o572(.A(ori_ori_n594_), .B(ori_ori_n251_), .Y(ori_ori_n595_));
  NA2        o573(.A(ori_ori_n595_), .B(ori_ori_n370_), .Y(ori_ori_n596_));
  OAI220     o574(.A0(ori_ori_n596_), .A1(ori_ori_n85_), .B0(ori_ori_n593_), .B1(ori_ori_n156_), .Y(ori_ori_n597_));
  NO2        o575(.A(ori_ori_n597_), .B(ori_ori_n314_), .Y(ori_ori_n598_));
  NA2        o576(.A(ori_ori_n598_), .B(ori_ori_n592_), .Y(ori_ori_n599_));
  NO3        o577(.A(ori_ori_n599_), .B(ori_ori_n590_), .C(ori_ori_n574_), .Y(ori_ori_n600_));
  AOI210     o578(.A0(ori_ori_n510_), .A1(ori_ori_n419_), .B0(ori_ori_n587_), .Y(ori_ori_n601_));
  INV        o579(.A(ori_ori_n601_), .Y(ori_ori_n602_));
  NA2        o580(.A(ori_ori_n182_), .B(ori_ori_n174_), .Y(ori_ori_n603_));
  AOI210     o581(.A0(ori_ori_n603_), .A1(ori_ori_n562_), .B0(ori_ori_n147_), .Y(ori_ori_n604_));
  INV        o582(.A(ori_ori_n604_), .Y(ori_ori_n605_));
  NA2        o583(.A(ori_ori_n605_), .B(ori_ori_n602_), .Y(ori_ori_n606_));
  NO3        o584(.A(ori_ori_n569_), .B(ori_ori_n556_), .C(ori_ori_n160_), .Y(ori_ori_n607_));
  AOI220     o585(.A0(ori_ori_n607_), .A1(i_11_), .B0(ori_ori_n333_), .B1(ori_ori_n74_), .Y(ori_ori_n608_));
  NO3        o586(.A(ori_ori_n167_), .B(ori_ori_n245_), .C(i_0_), .Y(ori_ori_n609_));
  OAI210     o587(.A0(ori_ori_n609_), .A1(ori_ori_n75_), .B0(i_13_), .Y(ori_ori_n610_));
  NA2        o588(.A(ori_ori_n610_), .B(ori_ori_n608_), .Y(ori_ori_n611_));
  NO3        o589(.A(ori_ori_n548_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n612_));
  NA2        o590(.A(ori_ori_n301_), .B(ori_ori_n294_), .Y(ori_ori_n613_));
  NO2        o591(.A(ori_ori_n613_), .B(ori_ori_n612_), .Y(ori_ori_n614_));
  NA3        o592(.A(ori_ori_n247_), .B(ori_ori_n155_), .C(ori_ori_n154_), .Y(ori_ori_n615_));
  INV        o593(.A(ori_ori_n615_), .Y(ori_ori_n616_));
  NO3        o594(.A(ori_ori_n576_), .B(ori_ori_n170_), .C(ori_ori_n160_), .Y(ori_ori_n617_));
  NO2        o595(.A(ori_ori_n617_), .B(ori_ori_n616_), .Y(ori_ori_n618_));
  NA2        o596(.A(ori_ori_n618_), .B(ori_ori_n614_), .Y(ori_ori_n619_));
  NO2        o597(.A(ori_ori_n85_), .B(i_5_), .Y(ori_ori_n620_));
  NA3        o598(.A(ori_ori_n543_), .B(ori_ori_n108_), .C(ori_ori_n122_), .Y(ori_ori_n621_));
  INV        o599(.A(ori_ori_n621_), .Y(ori_ori_n622_));
  NA2        o600(.A(ori_ori_n622_), .B(ori_ori_n620_), .Y(ori_ori_n623_));
  NAi21      o601(.An(ori_ori_n180_), .B(ori_ori_n181_), .Y(ori_ori_n624_));
  NO4        o602(.A(ori_ori_n179_), .B(ori_ori_n167_), .C(i_0_), .D(i_12_), .Y(ori_ori_n625_));
  NA2        o603(.A(ori_ori_n625_), .B(ori_ori_n624_), .Y(ori_ori_n626_));
  NA2        o604(.A(ori_ori_n626_), .B(ori_ori_n623_), .Y(ori_ori_n627_));
  NO4        o605(.A(ori_ori_n627_), .B(ori_ori_n619_), .C(ori_ori_n611_), .D(ori_ori_n606_), .Y(ori_ori_n628_));
  NA2        o606(.A(ori_ori_n524_), .B(ori_ori_n37_), .Y(ori_ori_n629_));
  NA2        o607(.A(ori_ori_n629_), .B(ori_ori_n363_), .Y(ori_ori_n630_));
  NA2        o608(.A(ori_ori_n630_), .B(ori_ori_n165_), .Y(ori_ori_n631_));
  NAi31      o609(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n632_));
  NO2        o610(.A(ori_ori_n69_), .B(ori_ori_n632_), .Y(ori_ori_n633_));
  AOI210     o611(.A0(ori_ori_n633_), .A1(ori_ori_n48_), .B0(ori_ori_n563_), .Y(ori_ori_n634_));
  AOI210     o612(.A0(ori_ori_n634_), .A1(ori_ori_n631_), .B0(ori_ori_n72_), .Y(ori_ori_n635_));
  INV        o613(.A(ori_ori_n242_), .Y(ori_ori_n636_));
  NO2        o614(.A(ori_ori_n636_), .B(ori_ori_n474_), .Y(ori_ori_n637_));
  NO3        o615(.A(ori_ori_n58_), .B(ori_ori_n57_), .C(i_4_), .Y(ori_ori_n638_));
  OAI210     o616(.A0(ori_ori_n589_), .A1(ori_ori_n208_), .B0(ori_ori_n638_), .Y(ori_ori_n639_));
  NO2        o617(.A(ori_ori_n639_), .B(ori_ori_n448_), .Y(ori_ori_n640_));
  NO3        o618(.A(ori_ori_n640_), .B(ori_ori_n637_), .C(ori_ori_n635_), .Y(ori_ori_n641_));
  NA4        o619(.A(ori_ori_n641_), .B(ori_ori_n628_), .C(ori_ori_n600_), .D(ori_ori_n561_), .Y(ori4));
  INV        o620(.A(ori_ori_n427_), .Y(ori_ori_n645_));
  INV        o621(.A(i_6_), .Y(ori_ori_n646_));
  INV        o622(.A(ori_ori_n214_), .Y(ori_ori_n647_));
  NAi21      m0000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m0001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m0002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m0003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m0004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m0005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m0006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m0007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m0008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m0010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m0011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m0012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m0013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m0014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m0015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m0016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m0017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m0018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m0019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m0021(.A(mai_mai_n35_), .Y(mai1));
  INV        m0022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m0023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m0024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m0025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m0026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m0027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m0028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m0029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m0030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m0031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m0032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NA2        m0033(.A(mai_mai_n53_), .B(mai_mai_n46_), .Y(mai_mai_n56_));
  NA3        m0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n57_));
  NO2        m0035(.A(i_1_), .B(i_6_), .Y(mai_mai_n58_));
  NA2        m0036(.A(i_8_), .B(i_7_), .Y(mai_mai_n59_));
  OAI210     m0037(.A0(mai_mai_n59_), .A1(mai_mai_n58_), .B0(mai_mai_n57_), .Y(mai_mai_n60_));
  NA2        m0038(.A(mai_mai_n60_), .B(i_12_), .Y(mai_mai_n61_));
  NAi21      m0039(.An(i_2_), .B(i_7_), .Y(mai_mai_n62_));
  INV        m0040(.A(i_1_), .Y(mai_mai_n63_));
  NA2        m0041(.A(mai_mai_n63_), .B(i_6_), .Y(mai_mai_n64_));
  NA3        m0042(.A(mai_mai_n64_), .B(mai_mai_n62_), .C(mai_mai_n31_), .Y(mai_mai_n65_));
  NA2        m0043(.A(i_1_), .B(i_10_), .Y(mai_mai_n66_));
  NO2        m0044(.A(mai_mai_n66_), .B(i_6_), .Y(mai_mai_n67_));
  NAi31      m0045(.An(mai_mai_n67_), .B(mai_mai_n65_), .C(mai_mai_n61_), .Y(mai_mai_n68_));
  NA2        m0046(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n69_));
  AOI210     m0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n70_));
  NA2        m0048(.A(i_1_), .B(i_6_), .Y(mai_mai_n71_));
  NO2        m0049(.A(mai_mai_n71_), .B(mai_mai_n25_), .Y(mai_mai_n72_));
  INV        m0050(.A(i_0_), .Y(mai_mai_n73_));
  NAi21      m0051(.An(i_5_), .B(i_10_), .Y(mai_mai_n74_));
  NA2        m0052(.A(i_5_), .B(i_9_), .Y(mai_mai_n75_));
  AOI210     m0053(.A0(mai_mai_n75_), .A1(mai_mai_n74_), .B0(mai_mai_n73_), .Y(mai_mai_n76_));
  NO2        m0054(.A(mai_mai_n76_), .B(mai_mai_n72_), .Y(mai_mai_n77_));
  OAI210     m0055(.A0(mai_mai_n70_), .A1(mai_mai_n69_), .B0(mai_mai_n77_), .Y(mai_mai_n78_));
  OAI210     m0056(.A0(mai_mai_n78_), .A1(mai_mai_n68_), .B0(i_0_), .Y(mai_mai_n79_));
  NA2        m0057(.A(i_12_), .B(i_5_), .Y(mai_mai_n80_));
  NA2        m0058(.A(i_2_), .B(i_8_), .Y(mai_mai_n81_));
  NO2        m0059(.A(mai_mai_n81_), .B(mai_mai_n58_), .Y(mai_mai_n82_));
  NO2        m0060(.A(i_3_), .B(i_9_), .Y(mai_mai_n83_));
  NO2        m0061(.A(i_3_), .B(i_7_), .Y(mai_mai_n84_));
  INV        m0062(.A(i_6_), .Y(mai_mai_n85_));
  OR4        m0063(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n86_));
  INV        m0064(.A(mai_mai_n86_), .Y(mai_mai_n87_));
  NO2        m0065(.A(i_2_), .B(i_7_), .Y(mai_mai_n88_));
  NAi21      m0066(.An(i_6_), .B(i_10_), .Y(mai_mai_n89_));
  NA2        m0067(.A(i_6_), .B(i_9_), .Y(mai_mai_n90_));
  AOI210     m0068(.A0(mai_mai_n90_), .A1(mai_mai_n89_), .B0(mai_mai_n63_), .Y(mai_mai_n91_));
  NA2        m0069(.A(i_2_), .B(i_6_), .Y(mai_mai_n92_));
  NO3        m0070(.A(mai_mai_n92_), .B(mai_mai_n50_), .C(mai_mai_n25_), .Y(mai_mai_n93_));
  NO2        m0071(.A(mai_mai_n93_), .B(mai_mai_n91_), .Y(mai_mai_n94_));
  AOI210     m0072(.A0(mai_mai_n94_), .A1(mai_mai_n1027_), .B0(mai_mai_n80_), .Y(mai_mai_n95_));
  AN3        m0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n96_));
  NAi21      m0074(.An(i_6_), .B(i_11_), .Y(mai_mai_n97_));
  NO2        m0075(.A(i_5_), .B(i_8_), .Y(mai_mai_n98_));
  NOi21      m0076(.An(mai_mai_n98_), .B(mai_mai_n97_), .Y(mai_mai_n99_));
  AOI220     m0077(.A0(mai_mai_n99_), .A1(mai_mai_n62_), .B0(mai_mai_n96_), .B1(mai_mai_n32_), .Y(mai_mai_n100_));
  INV        m0078(.A(i_7_), .Y(mai_mai_n101_));
  NA2        m0079(.A(mai_mai_n47_), .B(mai_mai_n101_), .Y(mai_mai_n102_));
  NO2        m0080(.A(i_0_), .B(i_5_), .Y(mai_mai_n103_));
  NO2        m0081(.A(mai_mai_n103_), .B(mai_mai_n85_), .Y(mai_mai_n104_));
  NA2        m0082(.A(i_12_), .B(i_3_), .Y(mai_mai_n105_));
  INV        m0083(.A(mai_mai_n105_), .Y(mai_mai_n106_));
  NA3        m0084(.A(mai_mai_n106_), .B(mai_mai_n104_), .C(mai_mai_n102_), .Y(mai_mai_n107_));
  NAi21      m0085(.An(i_7_), .B(i_11_), .Y(mai_mai_n108_));
  NO3        m0086(.A(mai_mai_n108_), .B(mai_mai_n89_), .C(mai_mai_n54_), .Y(mai_mai_n109_));
  AN2        m0087(.A(i_2_), .B(i_10_), .Y(mai_mai_n110_));
  NO2        m0088(.A(mai_mai_n110_), .B(i_7_), .Y(mai_mai_n111_));
  OR2        m0089(.A(mai_mai_n80_), .B(mai_mai_n58_), .Y(mai_mai_n112_));
  NO2        m0090(.A(i_8_), .B(mai_mai_n101_), .Y(mai_mai_n113_));
  NO3        m0091(.A(mai_mai_n113_), .B(mai_mai_n112_), .C(mai_mai_n111_), .Y(mai_mai_n114_));
  NA2        m0092(.A(i_12_), .B(i_7_), .Y(mai_mai_n115_));
  NO2        m0093(.A(mai_mai_n63_), .B(mai_mai_n26_), .Y(mai_mai_n116_));
  NA2        m0094(.A(mai_mai_n116_), .B(i_0_), .Y(mai_mai_n117_));
  NA2        m0095(.A(i_11_), .B(i_12_), .Y(mai_mai_n118_));
  OAI210     m0096(.A0(mai_mai_n117_), .A1(mai_mai_n115_), .B0(mai_mai_n118_), .Y(mai_mai_n119_));
  NO2        m0097(.A(mai_mai_n119_), .B(mai_mai_n114_), .Y(mai_mai_n120_));
  NAi41      m0098(.An(mai_mai_n109_), .B(mai_mai_n120_), .C(mai_mai_n107_), .D(mai_mai_n100_), .Y(mai_mai_n121_));
  NOi21      m0099(.An(i_1_), .B(i_5_), .Y(mai_mai_n122_));
  NA2        m0100(.A(mai_mai_n122_), .B(i_11_), .Y(mai_mai_n123_));
  NA2        m0101(.A(mai_mai_n101_), .B(mai_mai_n37_), .Y(mai_mai_n124_));
  NA2        m0102(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n125_));
  NA2        m0103(.A(mai_mai_n125_), .B(mai_mai_n124_), .Y(mai_mai_n126_));
  NO2        m0104(.A(mai_mai_n126_), .B(mai_mai_n47_), .Y(mai_mai_n127_));
  NA2        m0105(.A(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n128_));
  NAi21      m0106(.An(i_3_), .B(i_8_), .Y(mai_mai_n129_));
  NA2        m0107(.A(mai_mai_n129_), .B(mai_mai_n62_), .Y(mai_mai_n130_));
  NOi31      m0108(.An(mai_mai_n130_), .B(mai_mai_n128_), .C(mai_mai_n127_), .Y(mai_mai_n131_));
  NO2        m0109(.A(i_1_), .B(mai_mai_n85_), .Y(mai_mai_n132_));
  NO2        m0110(.A(i_6_), .B(i_5_), .Y(mai_mai_n133_));
  NA2        m0111(.A(mai_mai_n133_), .B(i_3_), .Y(mai_mai_n134_));
  OAI220     m0112(.A0(mai_mai_n134_), .A1(mai_mai_n108_), .B0(mai_mai_n131_), .B1(mai_mai_n123_), .Y(mai_mai_n135_));
  NO3        m0113(.A(mai_mai_n135_), .B(mai_mai_n121_), .C(mai_mai_n95_), .Y(mai_mai_n136_));
  NA3        m0114(.A(mai_mai_n136_), .B(mai_mai_n79_), .C(mai_mai_n56_), .Y(mai2));
  NO2        m0115(.A(mai_mai_n63_), .B(mai_mai_n37_), .Y(mai_mai_n138_));
  NA2        m0116(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n139_));
  NA2        m0117(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n140_));
  NA4        m0118(.A(mai_mai_n140_), .B(mai_mai_n77_), .C(mai_mai_n69_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m0119(.A(i_8_), .B(i_7_), .Y(mai_mai_n142_));
  NA2        m0120(.A(mai_mai_n142_), .B(i_6_), .Y(mai_mai_n143_));
  NO2        m0121(.A(i_12_), .B(i_13_), .Y(mai_mai_n144_));
  NAi21      m0122(.An(i_5_), .B(i_11_), .Y(mai_mai_n145_));
  NOi21      m0123(.An(mai_mai_n144_), .B(mai_mai_n145_), .Y(mai_mai_n146_));
  NO2        m0124(.A(i_0_), .B(i_1_), .Y(mai_mai_n147_));
  NA2        m0125(.A(i_2_), .B(i_3_), .Y(mai_mai_n148_));
  NO2        m0126(.A(mai_mai_n148_), .B(i_4_), .Y(mai_mai_n149_));
  NA2        m0127(.A(mai_mai_n149_), .B(mai_mai_n146_), .Y(mai_mai_n150_));
  AN2        m0128(.A(mai_mai_n144_), .B(mai_mai_n83_), .Y(mai_mai_n151_));
  NO2        m0129(.A(mai_mai_n151_), .B(mai_mai_n27_), .Y(mai_mai_n152_));
  NA2        m0130(.A(i_1_), .B(i_5_), .Y(mai_mai_n153_));
  NO2        m0131(.A(mai_mai_n73_), .B(mai_mai_n47_), .Y(mai_mai_n154_));
  NA2        m0132(.A(mai_mai_n154_), .B(mai_mai_n36_), .Y(mai_mai_n155_));
  NO3        m0133(.A(mai_mai_n155_), .B(mai_mai_n153_), .C(mai_mai_n152_), .Y(mai_mai_n156_));
  OR2        m0134(.A(i_0_), .B(i_1_), .Y(mai_mai_n157_));
  NO3        m0135(.A(mai_mai_n157_), .B(mai_mai_n80_), .C(i_13_), .Y(mai_mai_n158_));
  NAi32      m0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n159_));
  NAi21      m0137(.An(mai_mai_n159_), .B(mai_mai_n158_), .Y(mai_mai_n160_));
  NOi21      m0138(.An(i_4_), .B(i_10_), .Y(mai_mai_n161_));
  NA2        m0139(.A(mai_mai_n161_), .B(mai_mai_n40_), .Y(mai_mai_n162_));
  NO2        m0140(.A(i_3_), .B(i_5_), .Y(mai_mai_n163_));
  NO3        m0141(.A(mai_mai_n73_), .B(i_2_), .C(i_1_), .Y(mai_mai_n164_));
  NA2        m0142(.A(mai_mai_n164_), .B(mai_mai_n163_), .Y(mai_mai_n165_));
  OAI210     m0143(.A0(mai_mai_n165_), .A1(mai_mai_n162_), .B0(mai_mai_n160_), .Y(mai_mai_n166_));
  NO2        m0144(.A(mai_mai_n166_), .B(mai_mai_n156_), .Y(mai_mai_n167_));
  AOI210     m0145(.A0(mai_mai_n167_), .A1(mai_mai_n150_), .B0(mai_mai_n143_), .Y(mai_mai_n168_));
  NA2        m0146(.A(mai_mai_n73_), .B(i_1_), .Y(mai_mai_n169_));
  NA2        m0147(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n170_));
  NOi21      m0148(.An(i_4_), .B(i_9_), .Y(mai_mai_n171_));
  NOi21      m0149(.An(i_11_), .B(i_13_), .Y(mai_mai_n172_));
  NA2        m0150(.A(mai_mai_n172_), .B(mai_mai_n171_), .Y(mai_mai_n173_));
  OR2        m0151(.A(mai_mai_n173_), .B(mai_mai_n170_), .Y(mai_mai_n174_));
  NO2        m0152(.A(i_4_), .B(i_5_), .Y(mai_mai_n175_));
  NAi21      m0153(.An(i_12_), .B(i_11_), .Y(mai_mai_n176_));
  NO2        m0154(.A(mai_mai_n176_), .B(i_13_), .Y(mai_mai_n177_));
  NA3        m0155(.A(mai_mai_n177_), .B(mai_mai_n175_), .C(mai_mai_n83_), .Y(mai_mai_n178_));
  AOI210     m0156(.A0(mai_mai_n178_), .A1(mai_mai_n174_), .B0(mai_mai_n169_), .Y(mai_mai_n179_));
  NO2        m0157(.A(mai_mai_n73_), .B(mai_mai_n63_), .Y(mai_mai_n180_));
  NA2        m0158(.A(mai_mai_n180_), .B(mai_mai_n47_), .Y(mai_mai_n181_));
  NA2        m0159(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n182_));
  NAi31      m0160(.An(mai_mai_n182_), .B(mai_mai_n151_), .C(i_11_), .Y(mai_mai_n183_));
  NA2        m0161(.A(i_3_), .B(i_5_), .Y(mai_mai_n184_));
  OR2        m0162(.A(mai_mai_n184_), .B(mai_mai_n173_), .Y(mai_mai_n185_));
  AOI210     m0163(.A0(mai_mai_n185_), .A1(mai_mai_n183_), .B0(mai_mai_n181_), .Y(mai_mai_n186_));
  NO2        m0164(.A(mai_mai_n73_), .B(i_5_), .Y(mai_mai_n187_));
  NO2        m0165(.A(i_13_), .B(i_10_), .Y(mai_mai_n188_));
  NA3        m0166(.A(mai_mai_n188_), .B(mai_mai_n187_), .C(mai_mai_n45_), .Y(mai_mai_n189_));
  NO2        m0167(.A(i_2_), .B(i_1_), .Y(mai_mai_n190_));
  NA2        m0168(.A(mai_mai_n190_), .B(i_3_), .Y(mai_mai_n191_));
  NAi21      m0169(.An(i_4_), .B(i_12_), .Y(mai_mai_n192_));
  NO4        m0170(.A(mai_mai_n192_), .B(mai_mai_n191_), .C(mai_mai_n189_), .D(mai_mai_n25_), .Y(mai_mai_n193_));
  NO3        m0171(.A(mai_mai_n193_), .B(mai_mai_n186_), .C(mai_mai_n179_), .Y(mai_mai_n194_));
  INV        m0172(.A(i_8_), .Y(mai_mai_n195_));
  NA2        m0173(.A(i_8_), .B(i_6_), .Y(mai_mai_n196_));
  NO3        m0174(.A(i_3_), .B(mai_mai_n85_), .C(mai_mai_n49_), .Y(mai_mai_n197_));
  NA2        m0175(.A(mai_mai_n197_), .B(mai_mai_n113_), .Y(mai_mai_n198_));
  NO3        m0176(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n199_));
  NA3        m0177(.A(mai_mai_n199_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n200_));
  NO3        m0178(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n201_));
  OAI210     m0179(.A0(mai_mai_n96_), .A1(i_12_), .B0(mai_mai_n201_), .Y(mai_mai_n202_));
  AOI210     m0180(.A0(mai_mai_n202_), .A1(mai_mai_n200_), .B0(mai_mai_n198_), .Y(mai_mai_n203_));
  NO2        m0181(.A(i_3_), .B(i_8_), .Y(mai_mai_n204_));
  NO3        m0182(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n205_));
  NA3        m0183(.A(mai_mai_n205_), .B(mai_mai_n204_), .C(mai_mai_n40_), .Y(mai_mai_n206_));
  NO2        m0184(.A(i_13_), .B(i_9_), .Y(mai_mai_n207_));
  NA2        m0185(.A(mai_mai_n207_), .B(i_6_), .Y(mai_mai_n208_));
  NAi21      m0186(.An(i_12_), .B(i_3_), .Y(mai_mai_n209_));
  NO2        m0187(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n210_));
  NO3        m0188(.A(i_0_), .B(i_2_), .C(mai_mai_n63_), .Y(mai_mai_n211_));
  NA3        m0189(.A(mai_mai_n211_), .B(mai_mai_n210_), .C(i_10_), .Y(mai_mai_n212_));
  OAI220     m0190(.A0(mai_mai_n212_), .A1(mai_mai_n208_), .B0(mai_mai_n58_), .B1(mai_mai_n206_), .Y(mai_mai_n213_));
  AOI210     m0191(.A0(mai_mai_n213_), .A1(i_7_), .B0(mai_mai_n203_), .Y(mai_mai_n214_));
  OAI220     m0192(.A0(mai_mai_n214_), .A1(i_4_), .B0(mai_mai_n196_), .B1(mai_mai_n194_), .Y(mai_mai_n215_));
  NAi21      m0193(.An(i_12_), .B(i_7_), .Y(mai_mai_n216_));
  NA3        m0194(.A(i_13_), .B(mai_mai_n195_), .C(i_10_), .Y(mai_mai_n217_));
  NO2        m0195(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  NA2        m0196(.A(i_0_), .B(i_5_), .Y(mai_mai_n219_));
  OAI220     m0197(.A0(mai_mai_n85_), .A1(mai_mai_n191_), .B0(mai_mai_n181_), .B1(mai_mai_n134_), .Y(mai_mai_n220_));
  NAi31      m0198(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n221_));
  NO2        m0199(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n222_));
  NO2        m0200(.A(mai_mai_n73_), .B(mai_mai_n26_), .Y(mai_mai_n223_));
  NO2        m0201(.A(mai_mai_n47_), .B(mai_mai_n63_), .Y(mai_mai_n224_));
  NA3        m0202(.A(mai_mai_n224_), .B(mai_mai_n223_), .C(mai_mai_n222_), .Y(mai_mai_n225_));
  INV        m0203(.A(i_13_), .Y(mai_mai_n226_));
  NO2        m0204(.A(i_12_), .B(mai_mai_n226_), .Y(mai_mai_n227_));
  NA3        m0205(.A(mai_mai_n227_), .B(mai_mai_n199_), .C(mai_mai_n197_), .Y(mai_mai_n228_));
  OAI210     m0206(.A0(mai_mai_n225_), .A1(mai_mai_n221_), .B0(mai_mai_n228_), .Y(mai_mai_n229_));
  AOI220     m0207(.A0(mai_mai_n229_), .A1(mai_mai_n142_), .B0(mai_mai_n220_), .B1(mai_mai_n218_), .Y(mai_mai_n230_));
  NO2        m0208(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n231_));
  NO2        m0209(.A(mai_mai_n184_), .B(i_4_), .Y(mai_mai_n232_));
  NA2        m0210(.A(mai_mai_n232_), .B(mai_mai_n231_), .Y(mai_mai_n233_));
  OR2        m0211(.A(i_8_), .B(i_7_), .Y(mai_mai_n234_));
  NO2        m0212(.A(mai_mai_n234_), .B(mai_mai_n85_), .Y(mai_mai_n235_));
  NO2        m0213(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n236_));
  NA2        m0214(.A(mai_mai_n236_), .B(mai_mai_n235_), .Y(mai_mai_n237_));
  INV        m0215(.A(i_12_), .Y(mai_mai_n238_));
  NO2        m0216(.A(mai_mai_n45_), .B(mai_mai_n238_), .Y(mai_mai_n239_));
  NO3        m0217(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n240_));
  NA2        m0218(.A(i_2_), .B(i_1_), .Y(mai_mai_n241_));
  NO2        m0219(.A(mai_mai_n237_), .B(mai_mai_n233_), .Y(mai_mai_n242_));
  NO3        m0220(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n243_));
  NAi21      m0221(.An(i_4_), .B(i_3_), .Y(mai_mai_n244_));
  INV        m0222(.A(mai_mai_n75_), .Y(mai_mai_n245_));
  NO2        m0223(.A(i_0_), .B(i_6_), .Y(mai_mai_n246_));
  NOi41      m0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n247_));
  NA2        m0225(.A(mai_mai_n247_), .B(mai_mai_n246_), .Y(mai_mai_n248_));
  NO2        m0226(.A(mai_mai_n241_), .B(mai_mai_n184_), .Y(mai_mai_n249_));
  NAi21      m0227(.An(mai_mai_n248_), .B(mai_mai_n249_), .Y(mai_mai_n250_));
  INV        m0228(.A(mai_mai_n250_), .Y(mai_mai_n251_));
  AOI210     m0229(.A0(mai_mai_n251_), .A1(mai_mai_n40_), .B0(mai_mai_n242_), .Y(mai_mai_n252_));
  NO2        m0230(.A(i_11_), .B(mai_mai_n226_), .Y(mai_mai_n253_));
  NOi21      m0231(.An(i_1_), .B(i_6_), .Y(mai_mai_n254_));
  NAi21      m0232(.An(i_3_), .B(i_7_), .Y(mai_mai_n255_));
  NO2        m0233(.A(i_12_), .B(i_3_), .Y(mai_mai_n256_));
  NA2        m0234(.A(mai_mai_n73_), .B(i_5_), .Y(mai_mai_n257_));
  NAi21      m0235(.An(i_7_), .B(i_10_), .Y(mai_mai_n258_));
  NA3        m0236(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n259_));
  INV        m0237(.A(mai_mai_n143_), .Y(mai_mai_n260_));
  NA2        m0238(.A(mai_mai_n238_), .B(i_13_), .Y(mai_mai_n261_));
  NO2        m0239(.A(mai_mai_n261_), .B(mai_mai_n75_), .Y(mai_mai_n262_));
  NA2        m0240(.A(mai_mai_n262_), .B(mai_mai_n260_), .Y(mai_mai_n263_));
  NO2        m0241(.A(mai_mai_n234_), .B(mai_mai_n37_), .Y(mai_mai_n264_));
  NA2        m0242(.A(i_12_), .B(i_6_), .Y(mai_mai_n265_));
  OR2        m0243(.A(i_13_), .B(i_9_), .Y(mai_mai_n266_));
  NO3        m0244(.A(mai_mai_n266_), .B(mai_mai_n265_), .C(mai_mai_n49_), .Y(mai_mai_n267_));
  NO2        m0245(.A(mai_mai_n244_), .B(i_2_), .Y(mai_mai_n268_));
  NA3        m0246(.A(mai_mai_n268_), .B(mai_mai_n267_), .C(mai_mai_n45_), .Y(mai_mai_n269_));
  NA2        m0247(.A(mai_mai_n253_), .B(i_9_), .Y(mai_mai_n270_));
  NA2        m0248(.A(mai_mai_n257_), .B(mai_mai_n64_), .Y(mai_mai_n271_));
  OAI210     m0249(.A0(mai_mai_n271_), .A1(mai_mai_n270_), .B0(mai_mai_n269_), .Y(mai_mai_n272_));
  NA2        m0250(.A(mai_mai_n154_), .B(mai_mai_n63_), .Y(mai_mai_n273_));
  NO3        m0251(.A(i_11_), .B(mai_mai_n226_), .C(mai_mai_n25_), .Y(mai_mai_n274_));
  NO2        m0252(.A(mai_mai_n255_), .B(i_8_), .Y(mai_mai_n275_));
  NO2        m0253(.A(i_6_), .B(mai_mai_n49_), .Y(mai_mai_n276_));
  NA3        m0254(.A(mai_mai_n276_), .B(mai_mai_n275_), .C(mai_mai_n274_), .Y(mai_mai_n277_));
  NO3        m0255(.A(mai_mai_n26_), .B(mai_mai_n85_), .C(i_5_), .Y(mai_mai_n278_));
  NA3        m0256(.A(mai_mai_n278_), .B(mai_mai_n264_), .C(mai_mai_n227_), .Y(mai_mai_n279_));
  AOI210     m0257(.A0(mai_mai_n279_), .A1(mai_mai_n277_), .B0(mai_mai_n273_), .Y(mai_mai_n280_));
  AOI210     m0258(.A0(mai_mai_n272_), .A1(mai_mai_n264_), .B0(mai_mai_n280_), .Y(mai_mai_n281_));
  NA4        m0259(.A(mai_mai_n281_), .B(mai_mai_n263_), .C(mai_mai_n252_), .D(mai_mai_n230_), .Y(mai_mai_n282_));
  NO3        m0260(.A(i_12_), .B(mai_mai_n226_), .C(mai_mai_n37_), .Y(mai_mai_n283_));
  INV        m0261(.A(mai_mai_n283_), .Y(mai_mai_n284_));
  NA2        m0262(.A(i_8_), .B(mai_mai_n101_), .Y(mai_mai_n285_));
  NO3        m0263(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n286_));
  AOI220     m0264(.A0(mai_mai_n286_), .A1(mai_mai_n197_), .B0(mai_mai_n163_), .B1(mai_mai_n236_), .Y(mai_mai_n287_));
  NO2        m0265(.A(mai_mai_n287_), .B(mai_mai_n285_), .Y(mai_mai_n288_));
  NO2        m0266(.A(mai_mai_n241_), .B(i_0_), .Y(mai_mai_n289_));
  AOI220     m0267(.A0(mai_mai_n289_), .A1(i_8_), .B0(i_1_), .B1(mai_mai_n142_), .Y(mai_mai_n290_));
  NA2        m0268(.A(mai_mai_n276_), .B(mai_mai_n26_), .Y(mai_mai_n291_));
  NO2        m0269(.A(mai_mai_n291_), .B(mai_mai_n290_), .Y(mai_mai_n292_));
  NA2        m0270(.A(i_0_), .B(i_1_), .Y(mai_mai_n293_));
  NO2        m0271(.A(mai_mai_n293_), .B(i_2_), .Y(mai_mai_n294_));
  NO2        m0272(.A(mai_mai_n59_), .B(i_6_), .Y(mai_mai_n295_));
  NA3        m0273(.A(mai_mai_n295_), .B(mai_mai_n294_), .C(mai_mai_n163_), .Y(mai_mai_n296_));
  OAI210     m0274(.A0(mai_mai_n165_), .A1(mai_mai_n143_), .B0(mai_mai_n296_), .Y(mai_mai_n297_));
  NO3        m0275(.A(mai_mai_n297_), .B(mai_mai_n292_), .C(mai_mai_n288_), .Y(mai_mai_n298_));
  NO2        m0276(.A(i_3_), .B(i_10_), .Y(mai_mai_n299_));
  NA3        m0277(.A(mai_mai_n299_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n300_));
  NO2        m0278(.A(i_2_), .B(mai_mai_n101_), .Y(mai_mai_n301_));
  NA2        m0279(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n302_));
  NO2        m0280(.A(mai_mai_n302_), .B(i_8_), .Y(mai_mai_n303_));
  NA2        m0281(.A(mai_mai_n303_), .B(mai_mai_n301_), .Y(mai_mai_n304_));
  AN2        m0282(.A(i_3_), .B(i_10_), .Y(mai_mai_n305_));
  NA4        m0283(.A(mai_mai_n305_), .B(mai_mai_n199_), .C(mai_mai_n177_), .D(mai_mai_n175_), .Y(mai_mai_n306_));
  NO2        m0284(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n307_));
  NO2        m0285(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n308_));
  OR2        m0286(.A(mai_mai_n304_), .B(mai_mai_n300_), .Y(mai_mai_n309_));
  OAI220     m0287(.A0(mai_mai_n309_), .A1(i_6_), .B0(mai_mai_n298_), .B1(mai_mai_n284_), .Y(mai_mai_n310_));
  NO4        m0288(.A(mai_mai_n310_), .B(mai_mai_n282_), .C(mai_mai_n215_), .D(mai_mai_n168_), .Y(mai_mai_n311_));
  NO3        m0289(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n312_));
  NO2        m0290(.A(mai_mai_n59_), .B(mai_mai_n85_), .Y(mai_mai_n313_));
  NO3        m0291(.A(i_6_), .B(mai_mai_n195_), .C(i_7_), .Y(mai_mai_n314_));
  NA2        m0292(.A(mai_mai_n314_), .B(mai_mai_n199_), .Y(mai_mai_n315_));
  INV        m0293(.A(mai_mai_n315_), .Y(mai_mai_n316_));
  NO2        m0294(.A(i_2_), .B(i_3_), .Y(mai_mai_n317_));
  OR2        m0295(.A(i_0_), .B(i_5_), .Y(mai_mai_n318_));
  NA3        m0296(.A(mai_mai_n235_), .B(mai_mai_n317_), .C(i_1_), .Y(mai_mai_n319_));
  NA3        m0297(.A(mai_mai_n289_), .B(mai_mai_n163_), .C(mai_mai_n113_), .Y(mai_mai_n320_));
  NAi21      m0298(.An(i_8_), .B(i_7_), .Y(mai_mai_n321_));
  NO2        m0299(.A(mai_mai_n321_), .B(i_6_), .Y(mai_mai_n322_));
  NO2        m0300(.A(mai_mai_n157_), .B(mai_mai_n47_), .Y(mai_mai_n323_));
  NA3        m0301(.A(mai_mai_n323_), .B(mai_mai_n322_), .C(mai_mai_n163_), .Y(mai_mai_n324_));
  NA3        m0302(.A(mai_mai_n324_), .B(mai_mai_n320_), .C(mai_mai_n319_), .Y(mai_mai_n325_));
  OAI210     m0303(.A0(mai_mai_n325_), .A1(mai_mai_n316_), .B0(i_4_), .Y(mai_mai_n326_));
  NO2        m0304(.A(i_12_), .B(i_10_), .Y(mai_mai_n327_));
  NOi21      m0305(.An(i_5_), .B(i_0_), .Y(mai_mai_n328_));
  NO3        m0306(.A(mai_mai_n302_), .B(mai_mai_n328_), .C(mai_mai_n129_), .Y(mai_mai_n329_));
  NA4        m0307(.A(mai_mai_n84_), .B(mai_mai_n36_), .C(mai_mai_n85_), .D(i_8_), .Y(mai_mai_n330_));
  NA2        m0308(.A(mai_mai_n329_), .B(mai_mai_n327_), .Y(mai_mai_n331_));
  NO2        m0309(.A(i_6_), .B(i_8_), .Y(mai_mai_n332_));
  NOi21      m0310(.An(i_0_), .B(i_2_), .Y(mai_mai_n333_));
  AN2        m0311(.A(mai_mai_n333_), .B(mai_mai_n332_), .Y(mai_mai_n334_));
  NO2        m0312(.A(i_1_), .B(i_7_), .Y(mai_mai_n335_));
  AO220      m0313(.A0(mai_mai_n335_), .A1(mai_mai_n334_), .B0(mai_mai_n322_), .B1(mai_mai_n236_), .Y(mai_mai_n336_));
  NA2        m0314(.A(mai_mai_n336_), .B(mai_mai_n42_), .Y(mai_mai_n337_));
  NA3        m0315(.A(mai_mai_n337_), .B(mai_mai_n331_), .C(mai_mai_n326_), .Y(mai_mai_n338_));
  NO3        m0316(.A(mai_mai_n234_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n339_));
  NO3        m0317(.A(mai_mai_n321_), .B(i_2_), .C(i_1_), .Y(mai_mai_n340_));
  OAI210     m0318(.A0(mai_mai_n340_), .A1(mai_mai_n339_), .B0(i_6_), .Y(mai_mai_n341_));
  NA2        m0319(.A(mai_mai_n254_), .B(mai_mai_n301_), .Y(mai_mai_n342_));
  NA2        m0320(.A(mai_mai_n342_), .B(mai_mai_n341_), .Y(mai_mai_n343_));
  NA2        m0321(.A(mai_mai_n343_), .B(i_3_), .Y(mai_mai_n344_));
  INV        m0322(.A(mai_mai_n84_), .Y(mai_mai_n345_));
  NO2        m0323(.A(mai_mai_n293_), .B(mai_mai_n81_), .Y(mai_mai_n346_));
  NA2        m0324(.A(mai_mai_n346_), .B(mai_mai_n133_), .Y(mai_mai_n347_));
  NO2        m0325(.A(mai_mai_n92_), .B(mai_mai_n195_), .Y(mai_mai_n348_));
  NA2        m0326(.A(mai_mai_n348_), .B(mai_mai_n63_), .Y(mai_mai_n349_));
  AOI210     m0327(.A0(mai_mai_n349_), .A1(mai_mai_n347_), .B0(mai_mai_n345_), .Y(mai_mai_n350_));
  NO2        m0328(.A(mai_mai_n195_), .B(i_9_), .Y(mai_mai_n351_));
  NA2        m0329(.A(mai_mai_n351_), .B(i_6_), .Y(mai_mai_n352_));
  NO2        m0330(.A(mai_mai_n350_), .B(mai_mai_n292_), .Y(mai_mai_n353_));
  AOI210     m0331(.A0(mai_mai_n353_), .A1(mai_mai_n344_), .B0(mai_mai_n162_), .Y(mai_mai_n354_));
  AOI210     m0332(.A0(mai_mai_n338_), .A1(mai_mai_n312_), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  NOi32      m0333(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n356_));
  INV        m0334(.A(mai_mai_n356_), .Y(mai_mai_n357_));
  NAi21      m0335(.An(i_0_), .B(i_6_), .Y(mai_mai_n358_));
  NAi21      m0336(.An(i_1_), .B(i_5_), .Y(mai_mai_n359_));
  NA2        m0337(.A(mai_mai_n359_), .B(mai_mai_n358_), .Y(mai_mai_n360_));
  NA2        m0338(.A(mai_mai_n360_), .B(mai_mai_n25_), .Y(mai_mai_n361_));
  OAI210     m0339(.A0(mai_mai_n361_), .A1(mai_mai_n159_), .B0(mai_mai_n248_), .Y(mai_mai_n362_));
  NAi41      m0340(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n363_));
  OAI220     m0341(.A0(mai_mai_n363_), .A1(mai_mai_n359_), .B0(mai_mai_n221_), .B1(mai_mai_n159_), .Y(mai_mai_n364_));
  AOI210     m0342(.A0(mai_mai_n363_), .A1(mai_mai_n159_), .B0(mai_mai_n157_), .Y(mai_mai_n365_));
  NOi32      m0343(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n366_));
  NAi21      m0344(.An(i_6_), .B(i_1_), .Y(mai_mai_n367_));
  NA3        m0345(.A(mai_mai_n367_), .B(mai_mai_n366_), .C(mai_mai_n47_), .Y(mai_mai_n368_));
  NO2        m0346(.A(mai_mai_n368_), .B(i_0_), .Y(mai_mai_n369_));
  OR3        m0347(.A(mai_mai_n369_), .B(mai_mai_n365_), .C(mai_mai_n364_), .Y(mai_mai_n370_));
  NO2        m0348(.A(i_1_), .B(mai_mai_n101_), .Y(mai_mai_n371_));
  NAi21      m0349(.An(i_3_), .B(i_4_), .Y(mai_mai_n372_));
  NA2        m0350(.A(i_2_), .B(i_7_), .Y(mai_mai_n373_));
  NO2        m0351(.A(mai_mai_n372_), .B(i_10_), .Y(mai_mai_n374_));
  AOI210     m0352(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n375_));
  OAI210     m0353(.A0(mai_mai_n375_), .A1(mai_mai_n190_), .B0(mai_mai_n374_), .Y(mai_mai_n376_));
  AOI220     m0354(.A0(mai_mai_n374_), .A1(mai_mai_n335_), .B0(mai_mai_n240_), .B1(mai_mai_n190_), .Y(mai_mai_n377_));
  AOI210     m0355(.A0(mai_mai_n377_), .A1(mai_mai_n376_), .B0(i_5_), .Y(mai_mai_n378_));
  NO3        m0356(.A(mai_mai_n378_), .B(mai_mai_n370_), .C(mai_mai_n362_), .Y(mai_mai_n379_));
  NO2        m0357(.A(mai_mai_n379_), .B(mai_mai_n357_), .Y(mai_mai_n380_));
  NO2        m0358(.A(mai_mai_n59_), .B(mai_mai_n25_), .Y(mai_mai_n381_));
  AN2        m0359(.A(i_12_), .B(i_5_), .Y(mai_mai_n382_));
  NA2        m0360(.A(i_3_), .B(mai_mai_n382_), .Y(mai_mai_n383_));
  NO2        m0361(.A(i_11_), .B(i_6_), .Y(mai_mai_n384_));
  NA3        m0362(.A(mai_mai_n384_), .B(mai_mai_n323_), .C(mai_mai_n226_), .Y(mai_mai_n385_));
  NO2        m0363(.A(mai_mai_n385_), .B(mai_mai_n383_), .Y(mai_mai_n386_));
  NO2        m0364(.A(mai_mai_n244_), .B(i_5_), .Y(mai_mai_n387_));
  NO2        m0365(.A(i_5_), .B(i_10_), .Y(mai_mai_n388_));
  AOI220     m0366(.A0(mai_mai_n388_), .A1(mai_mai_n268_), .B0(mai_mai_n387_), .B1(mai_mai_n199_), .Y(mai_mai_n389_));
  NA2        m0367(.A(mai_mai_n144_), .B(mai_mai_n46_), .Y(mai_mai_n390_));
  NO2        m0368(.A(mai_mai_n390_), .B(mai_mai_n389_), .Y(mai_mai_n391_));
  OAI210     m0369(.A0(mai_mai_n391_), .A1(mai_mai_n386_), .B0(mai_mai_n381_), .Y(mai_mai_n392_));
  NO2        m0370(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n393_));
  NA2        m0371(.A(mai_mai_n386_), .B(mai_mai_n393_), .Y(mai_mai_n394_));
  NO3        m0372(.A(mai_mai_n85_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n395_));
  NA2        m0373(.A(mai_mai_n299_), .B(mai_mai_n90_), .Y(mai_mai_n396_));
  NO2        m0374(.A(i_11_), .B(i_12_), .Y(mai_mai_n397_));
  NA2        m0375(.A(mai_mai_n397_), .B(mai_mai_n36_), .Y(mai_mai_n398_));
  NO2        m0376(.A(mai_mai_n396_), .B(mai_mai_n398_), .Y(mai_mai_n399_));
  NA2        m0377(.A(mai_mai_n388_), .B(mai_mai_n238_), .Y(mai_mai_n400_));
  NA2        m0378(.A(mai_mai_n42_), .B(i_11_), .Y(mai_mai_n401_));
  NO2        m0379(.A(mai_mai_n401_), .B(mai_mai_n221_), .Y(mai_mai_n402_));
  NAi21      m0380(.An(i_13_), .B(i_0_), .Y(mai_mai_n403_));
  NO2        m0381(.A(mai_mai_n403_), .B(mai_mai_n241_), .Y(mai_mai_n404_));
  OAI210     m0382(.A0(mai_mai_n402_), .A1(mai_mai_n399_), .B0(mai_mai_n404_), .Y(mai_mai_n405_));
  NA3        m0383(.A(mai_mai_n405_), .B(mai_mai_n394_), .C(mai_mai_n392_), .Y(mai_mai_n406_));
  NA2        m0384(.A(mai_mai_n45_), .B(mai_mai_n226_), .Y(mai_mai_n407_));
  NO2        m0385(.A(i_0_), .B(i_11_), .Y(mai_mai_n408_));
  AN2        m0386(.A(i_1_), .B(i_6_), .Y(mai_mai_n409_));
  NOi21      m0387(.An(i_2_), .B(i_12_), .Y(mai_mai_n410_));
  NA2        m0388(.A(mai_mai_n410_), .B(mai_mai_n409_), .Y(mai_mai_n411_));
  INV        m0389(.A(mai_mai_n411_), .Y(mai_mai_n412_));
  NA2        m0390(.A(mai_mai_n142_), .B(i_9_), .Y(mai_mai_n413_));
  NO2        m0391(.A(mai_mai_n413_), .B(i_4_), .Y(mai_mai_n414_));
  NA2        m0392(.A(mai_mai_n412_), .B(mai_mai_n414_), .Y(mai_mai_n415_));
  NAi21      m0393(.An(i_9_), .B(i_4_), .Y(mai_mai_n416_));
  OR2        m0394(.A(i_13_), .B(i_10_), .Y(mai_mai_n417_));
  NO3        m0395(.A(mai_mai_n417_), .B(mai_mai_n118_), .C(mai_mai_n416_), .Y(mai_mai_n418_));
  NO2        m0396(.A(mai_mai_n173_), .B(mai_mai_n124_), .Y(mai_mai_n419_));
  OR2        m0397(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n420_));
  NO2        m0398(.A(mai_mai_n101_), .B(mai_mai_n25_), .Y(mai_mai_n421_));
  NA2        m0399(.A(mai_mai_n276_), .B(mai_mai_n211_), .Y(mai_mai_n422_));
  NO2        m0400(.A(mai_mai_n422_), .B(mai_mai_n420_), .Y(mai_mai_n423_));
  INV        m0401(.A(mai_mai_n423_), .Y(mai_mai_n424_));
  AOI210     m0402(.A0(mai_mai_n424_), .A1(mai_mai_n415_), .B0(mai_mai_n26_), .Y(mai_mai_n425_));
  NA2        m0403(.A(mai_mai_n320_), .B(mai_mai_n319_), .Y(mai_mai_n426_));
  AOI220     m0404(.A0(mai_mai_n295_), .A1(mai_mai_n286_), .B0(mai_mai_n289_), .B1(mai_mai_n313_), .Y(mai_mai_n427_));
  NO2        m0405(.A(mai_mai_n427_), .B(mai_mai_n170_), .Y(mai_mai_n428_));
  NO2        m0406(.A(mai_mai_n184_), .B(mai_mai_n85_), .Y(mai_mai_n429_));
  AOI220     m0407(.A0(mai_mai_n429_), .A1(mai_mai_n294_), .B0(mai_mai_n278_), .B1(mai_mai_n211_), .Y(mai_mai_n430_));
  NO2        m0408(.A(mai_mai_n430_), .B(mai_mai_n285_), .Y(mai_mai_n431_));
  NO3        m0409(.A(mai_mai_n431_), .B(mai_mai_n428_), .C(mai_mai_n426_), .Y(mai_mai_n432_));
  NA2        m0410(.A(mai_mai_n197_), .B(mai_mai_n96_), .Y(mai_mai_n433_));
  NA3        m0411(.A(mai_mai_n323_), .B(mai_mai_n163_), .C(mai_mai_n85_), .Y(mai_mai_n434_));
  AOI210     m0412(.A0(mai_mai_n434_), .A1(mai_mai_n433_), .B0(mai_mai_n321_), .Y(mai_mai_n435_));
  NA2        m0413(.A(mai_mai_n295_), .B(mai_mai_n236_), .Y(mai_mai_n436_));
  NO2        m0414(.A(mai_mai_n436_), .B(mai_mai_n184_), .Y(mai_mai_n437_));
  NO2        m0415(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n438_));
  NA3        m0416(.A(mai_mai_n335_), .B(mai_mai_n334_), .C(mai_mai_n438_), .Y(mai_mai_n439_));
  INV        m0417(.A(mai_mai_n314_), .Y(mai_mai_n440_));
  OAI210     m0418(.A0(mai_mai_n440_), .A1(mai_mai_n191_), .B0(mai_mai_n439_), .Y(mai_mai_n441_));
  NO3        m0419(.A(mai_mai_n441_), .B(mai_mai_n437_), .C(mai_mai_n435_), .Y(mai_mai_n442_));
  AOI210     m0420(.A0(mai_mai_n442_), .A1(mai_mai_n432_), .B0(mai_mai_n270_), .Y(mai_mai_n443_));
  NO4        m0421(.A(mai_mai_n443_), .B(mai_mai_n425_), .C(mai_mai_n406_), .D(mai_mai_n380_), .Y(mai_mai_n444_));
  NO2        m0422(.A(mai_mai_n73_), .B(i_13_), .Y(mai_mai_n445_));
  NO2        m0423(.A(i_10_), .B(i_9_), .Y(mai_mai_n446_));
  NAi21      m0424(.An(i_12_), .B(i_8_), .Y(mai_mai_n447_));
  NO2        m0425(.A(mai_mai_n447_), .B(i_3_), .Y(mai_mai_n448_));
  NO2        m0426(.A(mai_mai_n47_), .B(i_4_), .Y(mai_mai_n449_));
  NA2        m0427(.A(mai_mai_n449_), .B(mai_mai_n104_), .Y(mai_mai_n450_));
  NO2        m0428(.A(mai_mai_n450_), .B(mai_mai_n206_), .Y(mai_mai_n451_));
  NA2        m0429(.A(mai_mai_n308_), .B(i_0_), .Y(mai_mai_n452_));
  NO3        m0430(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n453_));
  NA2        m0431(.A(mai_mai_n265_), .B(mai_mai_n97_), .Y(mai_mai_n454_));
  NA2        m0432(.A(mai_mai_n454_), .B(mai_mai_n453_), .Y(mai_mai_n455_));
  NA2        m0433(.A(i_8_), .B(i_9_), .Y(mai_mai_n456_));
  NO2        m0434(.A(mai_mai_n455_), .B(mai_mai_n452_), .Y(mai_mai_n457_));
  NA2        m0435(.A(mai_mai_n253_), .B(mai_mai_n307_), .Y(mai_mai_n458_));
  NO3        m0436(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n459_));
  INV        m0437(.A(mai_mai_n459_), .Y(mai_mai_n460_));
  NA3        m0438(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n461_));
  NA4        m0439(.A(mai_mai_n145_), .B(mai_mai_n116_), .C(mai_mai_n80_), .D(mai_mai_n23_), .Y(mai_mai_n462_));
  OAI220     m0440(.A0(mai_mai_n462_), .A1(mai_mai_n461_), .B0(mai_mai_n460_), .B1(mai_mai_n458_), .Y(mai_mai_n463_));
  NO3        m0441(.A(mai_mai_n463_), .B(mai_mai_n457_), .C(mai_mai_n451_), .Y(mai_mai_n464_));
  OR2        m0442(.A(mai_mai_n293_), .B(mai_mai_n208_), .Y(mai_mai_n465_));
  OA210      m0443(.A0(mai_mai_n352_), .A1(mai_mai_n101_), .B0(mai_mai_n296_), .Y(mai_mai_n466_));
  OA220      m0444(.A0(mai_mai_n466_), .A1(mai_mai_n162_), .B0(mai_mai_n465_), .B1(mai_mai_n233_), .Y(mai_mai_n467_));
  NA2        m0445(.A(mai_mai_n96_), .B(i_13_), .Y(mai_mai_n468_));
  NA2        m0446(.A(mai_mai_n429_), .B(mai_mai_n381_), .Y(mai_mai_n469_));
  NO2        m0447(.A(i_2_), .B(i_13_), .Y(mai_mai_n470_));
  NA3        m0448(.A(mai_mai_n470_), .B(mai_mai_n161_), .C(mai_mai_n99_), .Y(mai_mai_n471_));
  NO2        m0449(.A(mai_mai_n469_), .B(mai_mai_n468_), .Y(mai_mai_n472_));
  NO3        m0450(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n473_));
  NO2        m0451(.A(i_6_), .B(i_7_), .Y(mai_mai_n474_));
  NA2        m0452(.A(mai_mai_n474_), .B(mai_mai_n473_), .Y(mai_mai_n475_));
  NO2        m0453(.A(i_11_), .B(i_1_), .Y(mai_mai_n476_));
  OR2        m0454(.A(i_11_), .B(i_8_), .Y(mai_mai_n477_));
  NOi21      m0455(.An(i_2_), .B(i_7_), .Y(mai_mai_n478_));
  NAi31      m0456(.An(mai_mai_n477_), .B(mai_mai_n478_), .C(i_0_), .Y(mai_mai_n479_));
  NO2        m0457(.A(mai_mai_n417_), .B(i_6_), .Y(mai_mai_n480_));
  NA2        m0458(.A(mai_mai_n480_), .B(i_1_), .Y(mai_mai_n481_));
  NO2        m0459(.A(mai_mai_n481_), .B(mai_mai_n479_), .Y(mai_mai_n482_));
  NO2        m0460(.A(i_3_), .B(mai_mai_n195_), .Y(mai_mai_n483_));
  NO2        m0461(.A(i_6_), .B(i_10_), .Y(mai_mai_n484_));
  NA4        m0462(.A(mai_mai_n484_), .B(mai_mai_n312_), .C(mai_mai_n483_), .D(mai_mai_n238_), .Y(mai_mai_n485_));
  NO2        m0463(.A(mai_mai_n485_), .B(mai_mai_n155_), .Y(mai_mai_n486_));
  NA2        m0464(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n487_));
  NO2        m0465(.A(mai_mai_n157_), .B(i_3_), .Y(mai_mai_n488_));
  NAi31      m0466(.An(mai_mai_n487_), .B(mai_mai_n488_), .C(mai_mai_n227_), .Y(mai_mai_n489_));
  NA3        m0467(.A(mai_mai_n393_), .B(mai_mai_n180_), .C(mai_mai_n149_), .Y(mai_mai_n490_));
  NA2        m0468(.A(mai_mai_n490_), .B(mai_mai_n489_), .Y(mai_mai_n491_));
  NO4        m0469(.A(mai_mai_n491_), .B(mai_mai_n486_), .C(mai_mai_n482_), .D(mai_mai_n472_), .Y(mai_mai_n492_));
  NA2        m0470(.A(mai_mai_n453_), .B(mai_mai_n382_), .Y(mai_mai_n493_));
  NAi21      m0471(.An(mai_mai_n217_), .B(mai_mai_n397_), .Y(mai_mai_n494_));
  NA2        m0472(.A(mai_mai_n335_), .B(mai_mai_n219_), .Y(mai_mai_n495_));
  NA3        m0473(.A(i_6_), .B(i_3_), .C(mai_mai_n142_), .Y(mai_mai_n496_));
  OR3        m0474(.A(mai_mai_n302_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n497_));
  OAI220     m0475(.A0(mai_mai_n497_), .A1(mai_mai_n496_), .B0(mai_mai_n495_), .B1(mai_mai_n494_), .Y(mai_mai_n498_));
  NA3        m0476(.A(mai_mai_n305_), .B(mai_mai_n224_), .C(mai_mai_n73_), .Y(mai_mai_n499_));
  NO2        m0477(.A(mai_mai_n499_), .B(mai_mai_n475_), .Y(mai_mai_n500_));
  NO2        m0478(.A(mai_mai_n500_), .B(mai_mai_n498_), .Y(mai_mai_n501_));
  NA4        m0479(.A(mai_mai_n501_), .B(mai_mai_n492_), .C(mai_mai_n467_), .D(mai_mai_n464_), .Y(mai_mai_n502_));
  NA3        m0480(.A(mai_mai_n305_), .B(mai_mai_n177_), .C(mai_mai_n175_), .Y(mai_mai_n503_));
  INV        m0481(.A(mai_mai_n503_), .Y(mai_mai_n504_));
  BUFFER     m0482(.A(mai_mai_n286_), .Y(mai_mai_n505_));
  NA2        m0483(.A(mai_mai_n505_), .B(mai_mai_n504_), .Y(mai_mai_n506_));
  NA2        m0484(.A(mai_mai_n123_), .B(mai_mai_n112_), .Y(mai_mai_n507_));
  AO220      m0485(.A0(mai_mai_n507_), .A1(mai_mai_n453_), .B0(mai_mai_n418_), .B1(i_6_), .Y(mai_mai_n508_));
  NA2        m0486(.A(mai_mai_n312_), .B(mai_mai_n164_), .Y(mai_mai_n509_));
  OAI210     m0487(.A0(mai_mai_n509_), .A1(mai_mai_n233_), .B0(mai_mai_n306_), .Y(mai_mai_n510_));
  AOI220     m0488(.A0(mai_mai_n510_), .A1(mai_mai_n322_), .B0(mai_mai_n508_), .B1(mai_mai_n308_), .Y(mai_mai_n511_));
  NA2        m0489(.A(mai_mai_n356_), .B(mai_mai_n73_), .Y(mai_mai_n512_));
  NO2        m0490(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n513_));
  AOI210     m0491(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n418_), .Y(mai_mai_n514_));
  NA2        m0492(.A(mai_mai_n257_), .B(mai_mai_n64_), .Y(mai_mai_n515_));
  OAI210     m0493(.A0(i_8_), .A1(mai_mai_n515_), .B0(mai_mai_n134_), .Y(mai_mai_n516_));
  NO2        m0494(.A(i_7_), .B(mai_mai_n200_), .Y(mai_mai_n517_));
  OR2        m0495(.A(mai_mai_n184_), .B(i_4_), .Y(mai_mai_n518_));
  NO2        m0496(.A(mai_mai_n518_), .B(mai_mai_n85_), .Y(mai_mai_n519_));
  AOI220     m0497(.A0(mai_mai_n519_), .A1(mai_mai_n517_), .B0(mai_mai_n516_), .B1(mai_mai_n419_), .Y(mai_mai_n520_));
  NA4        m0498(.A(mai_mai_n520_), .B(mai_mai_n514_), .C(mai_mai_n511_), .D(mai_mai_n506_), .Y(mai_mai_n521_));
  NA2        m0499(.A(mai_mai_n387_), .B(mai_mai_n294_), .Y(mai_mai_n522_));
  OAI210     m0500(.A0(mai_mai_n383_), .A1(mai_mai_n169_), .B0(mai_mai_n522_), .Y(mai_mai_n523_));
  NA2        m0501(.A(mai_mai_n1026_), .B(mai_mai_n226_), .Y(mai_mai_n524_));
  NA2        m0502(.A(mai_mai_n484_), .B(mai_mai_n27_), .Y(mai_mai_n525_));
  NO2        m0503(.A(mai_mai_n525_), .B(mai_mai_n524_), .Y(mai_mai_n526_));
  NOi31      m0504(.An(mai_mai_n314_), .B(mai_mai_n417_), .C(mai_mai_n38_), .Y(mai_mai_n527_));
  OAI210     m0505(.A0(mai_mai_n527_), .A1(mai_mai_n526_), .B0(mai_mai_n523_), .Y(mai_mai_n528_));
  NO2        m0506(.A(i_8_), .B(i_7_), .Y(mai_mai_n529_));
  OAI210     m0507(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n530_));
  NA2        m0508(.A(mai_mai_n530_), .B(mai_mai_n224_), .Y(mai_mai_n531_));
  OAI220     m0509(.A0(mai_mai_n47_), .A1(mai_mai_n518_), .B0(mai_mai_n531_), .B1(mai_mai_n244_), .Y(mai_mai_n532_));
  NA2        m0510(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n533_));
  NO2        m0511(.A(mai_mai_n533_), .B(i_6_), .Y(mai_mai_n534_));
  NA3        m0512(.A(mai_mai_n534_), .B(mai_mai_n532_), .C(mai_mai_n529_), .Y(mai_mai_n535_));
  AOI220     m0513(.A0(mai_mai_n429_), .A1(mai_mai_n323_), .B0(mai_mai_n249_), .B1(mai_mai_n246_), .Y(mai_mai_n536_));
  OAI220     m0514(.A0(mai_mai_n536_), .A1(mai_mai_n261_), .B0(mai_mai_n468_), .B1(mai_mai_n134_), .Y(mai_mai_n537_));
  NA2        m0515(.A(mai_mai_n537_), .B(mai_mai_n264_), .Y(mai_mai_n538_));
  NOi31      m0516(.An(mai_mai_n289_), .B(mai_mai_n300_), .C(mai_mai_n182_), .Y(mai_mai_n539_));
  NA3        m0517(.A(mai_mai_n305_), .B(mai_mai_n175_), .C(mai_mai_n96_), .Y(mai_mai_n540_));
  NO2        m0518(.A(mai_mai_n222_), .B(mai_mai_n45_), .Y(mai_mai_n541_));
  NO2        m0519(.A(mai_mai_n157_), .B(i_5_), .Y(mai_mai_n542_));
  NA3        m0520(.A(mai_mai_n542_), .B(mai_mai_n407_), .C(mai_mai_n317_), .Y(mai_mai_n543_));
  OAI210     m0521(.A0(mai_mai_n543_), .A1(mai_mai_n541_), .B0(mai_mai_n540_), .Y(mai_mai_n544_));
  OAI210     m0522(.A0(mai_mai_n544_), .A1(mai_mai_n539_), .B0(mai_mai_n459_), .Y(mai_mai_n545_));
  NA4        m0523(.A(mai_mai_n545_), .B(mai_mai_n538_), .C(mai_mai_n535_), .D(mai_mai_n528_), .Y(mai_mai_n546_));
  NA2        m0524(.A(mai_mai_n283_), .B(mai_mai_n84_), .Y(mai_mai_n547_));
  NO2        m0525(.A(mai_mai_n347_), .B(mai_mai_n547_), .Y(mai_mai_n548_));
  NA2        m0526(.A(mai_mai_n295_), .B(mai_mai_n286_), .Y(mai_mai_n549_));
  NO2        m0527(.A(mai_mai_n549_), .B(mai_mai_n174_), .Y(mai_mai_n550_));
  NA2        m0528(.A(mai_mai_n224_), .B(mai_mai_n223_), .Y(mai_mai_n551_));
  NA2        m0529(.A(mai_mai_n446_), .B(mai_mai_n222_), .Y(mai_mai_n552_));
  NO2        m0530(.A(mai_mai_n551_), .B(mai_mai_n552_), .Y(mai_mai_n553_));
  NO3        m0531(.A(mai_mai_n553_), .B(mai_mai_n550_), .C(mai_mai_n548_), .Y(mai_mai_n554_));
  NO4        m0532(.A(mai_mai_n254_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n555_));
  NO3        m0533(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n556_));
  NO2        m0534(.A(mai_mai_n234_), .B(mai_mai_n36_), .Y(mai_mai_n557_));
  AN2        m0535(.A(mai_mai_n557_), .B(mai_mai_n556_), .Y(mai_mai_n558_));
  OA210      m0536(.A0(mai_mai_n558_), .A1(mai_mai_n555_), .B0(mai_mai_n356_), .Y(mai_mai_n559_));
  NO2        m0537(.A(mai_mai_n417_), .B(i_1_), .Y(mai_mai_n560_));
  NOi31      m0538(.An(mai_mai_n560_), .B(mai_mai_n454_), .C(mai_mai_n73_), .Y(mai_mai_n561_));
  AN4        m0539(.A(mai_mai_n561_), .B(mai_mai_n414_), .C(i_3_), .D(i_2_), .Y(mai_mai_n562_));
  NO2        m0540(.A(mai_mai_n427_), .B(mai_mai_n178_), .Y(mai_mai_n563_));
  NO3        m0541(.A(mai_mai_n563_), .B(mai_mai_n562_), .C(mai_mai_n559_), .Y(mai_mai_n564_));
  NOi21      m0542(.An(i_10_), .B(i_6_), .Y(mai_mai_n565_));
  NO2        m0543(.A(mai_mai_n85_), .B(mai_mai_n25_), .Y(mai_mai_n566_));
  AOI220     m0544(.A0(mai_mai_n283_), .A1(mai_mai_n566_), .B0(mai_mai_n274_), .B1(mai_mai_n565_), .Y(mai_mai_n567_));
  NO2        m0545(.A(mai_mai_n567_), .B(mai_mai_n452_), .Y(mai_mai_n568_));
  NO2        m0546(.A(mai_mai_n115_), .B(mai_mai_n23_), .Y(mai_mai_n569_));
  NA2        m0547(.A(mai_mai_n314_), .B(mai_mai_n164_), .Y(mai_mai_n570_));
  AOI220     m0548(.A0(mai_mai_n570_), .A1(mai_mai_n436_), .B0(mai_mai_n185_), .B1(mai_mai_n183_), .Y(mai_mai_n571_));
  NOi21      m0549(.An(mai_mai_n146_), .B(mai_mai_n330_), .Y(mai_mai_n572_));
  NO3        m0550(.A(mai_mai_n572_), .B(mai_mai_n571_), .C(mai_mai_n568_), .Y(mai_mai_n573_));
  NO2        m0551(.A(mai_mai_n512_), .B(mai_mai_n377_), .Y(mai_mai_n574_));
  INV        m0552(.A(mai_mai_n317_), .Y(mai_mai_n575_));
  NO2        m0553(.A(i_12_), .B(mai_mai_n85_), .Y(mai_mai_n576_));
  NA3        m0554(.A(mai_mai_n576_), .B(mai_mai_n274_), .C(i_5_), .Y(mai_mai_n577_));
  NA3        m0555(.A(mai_mai_n384_), .B(mai_mai_n283_), .C(mai_mai_n219_), .Y(mai_mai_n578_));
  AOI210     m0556(.A0(mai_mai_n578_), .A1(mai_mai_n577_), .B0(mai_mai_n575_), .Y(mai_mai_n579_));
  NO3        m0557(.A(i_4_), .B(mai_mai_n341_), .C(mai_mai_n300_), .Y(mai_mai_n580_));
  NO3        m0558(.A(mai_mai_n580_), .B(mai_mai_n579_), .C(mai_mai_n574_), .Y(mai_mai_n581_));
  NA4        m0559(.A(mai_mai_n581_), .B(mai_mai_n573_), .C(mai_mai_n564_), .D(mai_mai_n554_), .Y(mai_mai_n582_));
  NO4        m0560(.A(mai_mai_n582_), .B(mai_mai_n546_), .C(mai_mai_n521_), .D(mai_mai_n502_), .Y(mai_mai_n583_));
  NA4        m0561(.A(mai_mai_n583_), .B(mai_mai_n444_), .C(mai_mai_n355_), .D(mai_mai_n311_), .Y(mai7));
  NO2        m0562(.A(mai_mai_n92_), .B(mai_mai_n55_), .Y(mai_mai_n585_));
  NO2        m0563(.A(mai_mai_n108_), .B(mai_mai_n89_), .Y(mai_mai_n586_));
  NA2        m0564(.A(i_3_), .B(mai_mai_n586_), .Y(mai_mai_n587_));
  NA2        m0565(.A(i_11_), .B(mai_mai_n195_), .Y(mai_mai_n588_));
  INV        m0566(.A(mai_mai_n587_), .Y(mai_mai_n589_));
  NA3        m0567(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n590_));
  NO2        m0568(.A(mai_mai_n238_), .B(i_4_), .Y(mai_mai_n591_));
  NA2        m0569(.A(mai_mai_n591_), .B(i_8_), .Y(mai_mai_n592_));
  NO2        m0570(.A(mai_mai_n105_), .B(mai_mai_n590_), .Y(mai_mai_n593_));
  NA2        m0571(.A(i_2_), .B(mai_mai_n85_), .Y(mai_mai_n594_));
  OAI210     m0572(.A0(mai_mai_n88_), .A1(mai_mai_n204_), .B0(mai_mai_n205_), .Y(mai_mai_n595_));
  NO2        m0573(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n596_));
  NA2        m0574(.A(i_4_), .B(i_8_), .Y(mai_mai_n597_));
  AOI210     m0575(.A0(mai_mai_n597_), .A1(mai_mai_n305_), .B0(mai_mai_n596_), .Y(mai_mai_n598_));
  OAI220     m0576(.A0(mai_mai_n598_), .A1(mai_mai_n594_), .B0(mai_mai_n595_), .B1(i_13_), .Y(mai_mai_n599_));
  NO4        m0577(.A(mai_mai_n599_), .B(mai_mai_n593_), .C(mai_mai_n589_), .D(mai_mai_n585_), .Y(mai_mai_n600_));
  AOI210     m0578(.A0(mai_mai_n129_), .A1(mai_mai_n62_), .B0(i_10_), .Y(mai_mai_n601_));
  AOI210     m0579(.A0(mai_mai_n601_), .A1(mai_mai_n238_), .B0(mai_mai_n161_), .Y(mai_mai_n602_));
  OR2        m0580(.A(i_6_), .B(i_10_), .Y(mai_mai_n603_));
  NO2        m0581(.A(mai_mai_n603_), .B(mai_mai_n23_), .Y(mai_mai_n604_));
  OR3        m0582(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n605_));
  NO3        m0583(.A(mai_mai_n605_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n606_));
  INV        m0584(.A(mai_mai_n201_), .Y(mai_mai_n607_));
  NO2        m0585(.A(mai_mai_n606_), .B(mai_mai_n604_), .Y(mai_mai_n608_));
  OA220      m0586(.A0(mai_mai_n608_), .A1(mai_mai_n575_), .B0(mai_mai_n602_), .B1(mai_mai_n266_), .Y(mai_mai_n609_));
  AOI210     m0587(.A0(mai_mai_n609_), .A1(mai_mai_n600_), .B0(mai_mai_n63_), .Y(mai_mai_n610_));
  NOi21      m0588(.An(i_11_), .B(i_7_), .Y(mai_mai_n611_));
  AO210      m0589(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n612_));
  NO2        m0590(.A(mai_mai_n612_), .B(mai_mai_n611_), .Y(mai_mai_n613_));
  NA2        m0591(.A(mai_mai_n613_), .B(mai_mai_n207_), .Y(mai_mai_n614_));
  NA3        m0592(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n615_));
  NAi31      m0593(.An(mai_mai_n615_), .B(mai_mai_n216_), .C(i_11_), .Y(mai_mai_n616_));
  AOI210     m0594(.A0(mai_mai_n616_), .A1(mai_mai_n614_), .B0(mai_mai_n63_), .Y(mai_mai_n617_));
  NA2        m0595(.A(mai_mai_n87_), .B(mai_mai_n63_), .Y(mai_mai_n618_));
  AO210      m0596(.A0(mai_mai_n618_), .A1(mai_mai_n377_), .B0(mai_mai_n41_), .Y(mai_mai_n619_));
  NO3        m0597(.A(mai_mai_n258_), .B(mai_mai_n209_), .C(mai_mai_n588_), .Y(mai_mai_n620_));
  OAI210     m0598(.A0(mai_mai_n620_), .A1(mai_mai_n227_), .B0(mai_mai_n63_), .Y(mai_mai_n621_));
  NA2        m0599(.A(mai_mai_n410_), .B(mai_mai_n31_), .Y(mai_mai_n622_));
  OR2        m0600(.A(mai_mai_n209_), .B(mai_mai_n108_), .Y(mai_mai_n623_));
  NA2        m0601(.A(mai_mai_n623_), .B(mai_mai_n622_), .Y(mai_mai_n624_));
  NO2        m0602(.A(mai_mai_n63_), .B(i_9_), .Y(mai_mai_n625_));
  NO2        m0603(.A(mai_mai_n625_), .B(i_4_), .Y(mai_mai_n626_));
  NA2        m0604(.A(mai_mai_n626_), .B(mai_mai_n624_), .Y(mai_mai_n627_));
  NO2        m0605(.A(i_1_), .B(i_12_), .Y(mai_mai_n628_));
  NA3        m0606(.A(mai_mai_n628_), .B(mai_mai_n110_), .C(mai_mai_n24_), .Y(mai_mai_n629_));
  NA4        m0607(.A(mai_mai_n629_), .B(mai_mai_n627_), .C(mai_mai_n621_), .D(mai_mai_n619_), .Y(mai_mai_n630_));
  OAI210     m0608(.A0(mai_mai_n630_), .A1(mai_mai_n617_), .B0(i_6_), .Y(mai_mai_n631_));
  NO2        m0609(.A(i_6_), .B(i_11_), .Y(mai_mai_n632_));
  INV        m0610(.A(mai_mai_n455_), .Y(mai_mai_n633_));
  NO4        m0611(.A(mai_mai_n216_), .B(mai_mai_n129_), .C(i_13_), .D(mai_mai_n85_), .Y(mai_mai_n634_));
  NA2        m0612(.A(mai_mai_n634_), .B(mai_mai_n625_), .Y(mai_mai_n635_));
  INV        m0613(.A(mai_mai_n635_), .Y(mai_mai_n636_));
  NA3        m0614(.A(mai_mai_n529_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n637_));
  NA2        m0615(.A(mai_mai_n138_), .B(i_9_), .Y(mai_mai_n638_));
  NA3        m0616(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n639_));
  NO2        m0617(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n640_));
  NA3        m0618(.A(mai_mai_n640_), .B(mai_mai_n265_), .C(mai_mai_n45_), .Y(mai_mai_n641_));
  OAI220     m0619(.A0(mai_mai_n641_), .A1(mai_mai_n639_), .B0(mai_mai_n638_), .B1(mai_mai_n1024_), .Y(mai_mai_n642_));
  NA3        m0620(.A(mai_mai_n625_), .B(mai_mai_n317_), .C(i_6_), .Y(mai_mai_n643_));
  NO2        m0621(.A(mai_mai_n643_), .B(mai_mai_n23_), .Y(mai_mai_n644_));
  AOI210     m0622(.A0(mai_mai_n476_), .A1(mai_mai_n421_), .B0(mai_mai_n243_), .Y(mai_mai_n645_));
  NO2        m0623(.A(mai_mai_n645_), .B(mai_mai_n594_), .Y(mai_mai_n646_));
  NAi21      m0624(.An(mai_mai_n637_), .B(mai_mai_n91_), .Y(mai_mai_n647_));
  NA2        m0625(.A(mai_mai_n640_), .B(mai_mai_n265_), .Y(mai_mai_n648_));
  NO2        m0626(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n649_));
  NA2        m0627(.A(mai_mai_n649_), .B(mai_mai_n24_), .Y(mai_mai_n650_));
  OAI210     m0628(.A0(mai_mai_n650_), .A1(mai_mai_n648_), .B0(mai_mai_n647_), .Y(mai_mai_n651_));
  OR4        m0629(.A(mai_mai_n651_), .B(mai_mai_n646_), .C(mai_mai_n644_), .D(mai_mai_n642_), .Y(mai_mai_n652_));
  NO3        m0630(.A(mai_mai_n652_), .B(mai_mai_n636_), .C(mai_mai_n633_), .Y(mai_mai_n653_));
  NO2        m0631(.A(mai_mai_n238_), .B(mai_mai_n101_), .Y(mai_mai_n654_));
  NO2        m0632(.A(mai_mai_n654_), .B(mai_mai_n611_), .Y(mai_mai_n655_));
  NA2        m0633(.A(mai_mai_n655_), .B(i_1_), .Y(mai_mai_n656_));
  NO2        m0634(.A(mai_mai_n656_), .B(mai_mai_n605_), .Y(mai_mai_n657_));
  NA2        m0635(.A(mai_mai_n657_), .B(mai_mai_n47_), .Y(mai_mai_n658_));
  NO2        m0636(.A(mai_mai_n234_), .B(mai_mai_n45_), .Y(mai_mai_n659_));
  NO3        m0637(.A(mai_mai_n659_), .B(mai_mai_n308_), .C(mai_mai_n239_), .Y(mai_mai_n660_));
  NO2        m0638(.A(mai_mai_n118_), .B(mai_mai_n37_), .Y(mai_mai_n661_));
  NO2        m0639(.A(mai_mai_n661_), .B(i_6_), .Y(mai_mai_n662_));
  NO2        m0640(.A(mai_mai_n85_), .B(i_9_), .Y(mai_mai_n663_));
  NO2        m0641(.A(mai_mai_n663_), .B(mai_mai_n63_), .Y(mai_mai_n664_));
  NO2        m0642(.A(mai_mai_n664_), .B(mai_mai_n628_), .Y(mai_mai_n665_));
  NO4        m0643(.A(mai_mai_n665_), .B(mai_mai_n662_), .C(mai_mai_n660_), .D(i_4_), .Y(mai_mai_n666_));
  NA2        m0644(.A(i_1_), .B(i_3_), .Y(mai_mai_n667_));
  INV        m0645(.A(mai_mai_n666_), .Y(mai_mai_n668_));
  NA4        m0646(.A(mai_mai_n668_), .B(mai_mai_n658_), .C(mai_mai_n653_), .D(mai_mai_n631_), .Y(mai_mai_n669_));
  NO3        m0647(.A(mai_mai_n477_), .B(i_3_), .C(i_7_), .Y(mai_mai_n670_));
  NOi21      m0648(.An(mai_mai_n670_), .B(i_10_), .Y(mai_mai_n671_));
  OA210      m0649(.A0(mai_mai_n671_), .A1(mai_mai_n247_), .B0(mai_mai_n85_), .Y(mai_mai_n672_));
  NA3        m0650(.A(mai_mai_n484_), .B(mai_mai_n513_), .C(mai_mai_n47_), .Y(mai_mai_n673_));
  NO3        m0651(.A(mai_mai_n478_), .B(mai_mai_n597_), .C(mai_mai_n85_), .Y(mai_mai_n674_));
  NA2        m0652(.A(mai_mai_n674_), .B(mai_mai_n25_), .Y(mai_mai_n675_));
  NA3        m0653(.A(mai_mai_n161_), .B(mai_mai_n84_), .C(mai_mai_n85_), .Y(mai_mai_n676_));
  NA3        m0654(.A(mai_mai_n676_), .B(mai_mai_n675_), .C(mai_mai_n673_), .Y(mai_mai_n677_));
  OAI210     m0655(.A0(mai_mai_n677_), .A1(mai_mai_n672_), .B0(i_1_), .Y(mai_mai_n678_));
  AOI210     m0656(.A0(mai_mai_n265_), .A1(mai_mai_n97_), .B0(i_1_), .Y(mai_mai_n679_));
  NO2        m0657(.A(mai_mai_n372_), .B(i_2_), .Y(mai_mai_n680_));
  NA2        m0658(.A(mai_mai_n680_), .B(mai_mai_n679_), .Y(mai_mai_n681_));
  OAI210     m0659(.A0(mai_mai_n643_), .A1(mai_mai_n447_), .B0(mai_mai_n681_), .Y(mai_mai_n682_));
  INV        m0660(.A(mai_mai_n682_), .Y(mai_mai_n683_));
  AOI210     m0661(.A0(mai_mai_n683_), .A1(mai_mai_n678_), .B0(i_13_), .Y(mai_mai_n684_));
  OR2        m0662(.A(i_11_), .B(i_7_), .Y(mai_mai_n685_));
  NA3        m0663(.A(mai_mai_n685_), .B(mai_mai_n106_), .C(mai_mai_n138_), .Y(mai_mai_n686_));
  AOI220     m0664(.A0(mai_mai_n470_), .A1(mai_mai_n161_), .B0(mai_mai_n449_), .B1(mai_mai_n138_), .Y(mai_mai_n687_));
  OAI210     m0665(.A0(mai_mai_n687_), .A1(mai_mai_n45_), .B0(mai_mai_n686_), .Y(mai_mai_n688_));
  AOI210     m0666(.A0(mai_mai_n639_), .A1(mai_mai_n55_), .B0(i_12_), .Y(mai_mai_n689_));
  INV        m0667(.A(mai_mai_n689_), .Y(mai_mai_n690_));
  NA2        m0668(.A(mai_mai_n247_), .B(mai_mai_n132_), .Y(mai_mai_n691_));
  OAI220     m0669(.A0(mai_mai_n691_), .A1(mai_mai_n41_), .B0(mai_mai_n690_), .B1(mai_mai_n92_), .Y(mai_mai_n692_));
  AOI210     m0670(.A0(mai_mai_n688_), .A1(mai_mai_n332_), .B0(mai_mai_n692_), .Y(mai_mai_n693_));
  INV        m0671(.A(mai_mai_n115_), .Y(mai_mai_n694_));
  AOI220     m0672(.A0(mai_mai_n694_), .A1(mai_mai_n72_), .B0(mai_mai_n384_), .B1(mai_mai_n640_), .Y(mai_mai_n695_));
  NO2        m0673(.A(mai_mai_n695_), .B(mai_mai_n244_), .Y(mai_mai_n696_));
  AOI210     m0674(.A0(mai_mai_n447_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n697_));
  NA2        m0675(.A(mai_mai_n128_), .B(i_13_), .Y(mai_mai_n698_));
  NO2        m0676(.A(mai_mai_n639_), .B(mai_mai_n115_), .Y(mai_mai_n699_));
  INV        m0677(.A(mai_mai_n699_), .Y(mai_mai_n700_));
  OAI220     m0678(.A0(mai_mai_n700_), .A1(mai_mai_n71_), .B0(mai_mai_n698_), .B1(mai_mai_n679_), .Y(mai_mai_n701_));
  NO3        m0679(.A(mai_mai_n71_), .B(mai_mai_n32_), .C(mai_mai_n101_), .Y(mai_mai_n702_));
  NA2        m0680(.A(mai_mai_n26_), .B(mai_mai_n195_), .Y(mai_mai_n703_));
  INV        m0681(.A(mai_mai_n703_), .Y(mai_mai_n704_));
  NO3        m0682(.A(mai_mai_n478_), .B(mai_mai_n238_), .C(mai_mai_n85_), .Y(mai_mai_n705_));
  AOI210     m0683(.A0(mai_mai_n705_), .A1(mai_mai_n704_), .B0(mai_mai_n702_), .Y(mai_mai_n706_));
  NA2        m0684(.A(mai_mai_n91_), .B(mai_mai_n102_), .Y(mai_mai_n707_));
  OAI220     m0685(.A0(mai_mai_n707_), .A1(mai_mai_n592_), .B0(mai_mai_n706_), .B1(mai_mai_n607_), .Y(mai_mai_n708_));
  NO3        m0686(.A(mai_mai_n708_), .B(mai_mai_n701_), .C(mai_mai_n696_), .Y(mai_mai_n709_));
  OR2        m0687(.A(i_11_), .B(i_6_), .Y(mai_mai_n710_));
  NA3        m0688(.A(mai_mai_n591_), .B(mai_mai_n703_), .C(i_7_), .Y(mai_mai_n711_));
  AOI210     m0689(.A0(mai_mai_n711_), .A1(mai_mai_n700_), .B0(mai_mai_n710_), .Y(mai_mai_n712_));
  NA3        m0690(.A(mai_mai_n410_), .B(mai_mai_n596_), .C(mai_mai_n97_), .Y(mai_mai_n713_));
  NA2        m0691(.A(mai_mai_n632_), .B(i_13_), .Y(mai_mai_n714_));
  NA2        m0692(.A(mai_mai_n102_), .B(mai_mai_n703_), .Y(mai_mai_n715_));
  NAi21      m0693(.An(i_11_), .B(i_12_), .Y(mai_mai_n716_));
  NOi41      m0694(.An(mai_mai_n111_), .B(mai_mai_n716_), .C(i_13_), .D(mai_mai_n85_), .Y(mai_mai_n717_));
  NO3        m0695(.A(mai_mai_n478_), .B(mai_mai_n576_), .C(mai_mai_n597_), .Y(mai_mai_n718_));
  AOI220     m0696(.A0(mai_mai_n718_), .A1(mai_mai_n312_), .B0(mai_mai_n717_), .B1(mai_mai_n715_), .Y(mai_mai_n719_));
  NA3        m0697(.A(mai_mai_n719_), .B(mai_mai_n714_), .C(mai_mai_n713_), .Y(mai_mai_n720_));
  OAI210     m0698(.A0(mai_mai_n720_), .A1(mai_mai_n712_), .B0(mai_mai_n63_), .Y(mai_mai_n721_));
  NO2        m0699(.A(i_2_), .B(i_12_), .Y(mai_mai_n722_));
  NA2        m0700(.A(mai_mai_n371_), .B(mai_mai_n722_), .Y(mai_mai_n723_));
  NO3        m0701(.A(i_9_), .B(i_3_), .C(mai_mai_n591_), .Y(mai_mai_n724_));
  NA2        m0702(.A(mai_mai_n724_), .B(mai_mai_n371_), .Y(mai_mai_n725_));
  NO2        m0703(.A(mai_mai_n129_), .B(i_2_), .Y(mai_mai_n726_));
  NA2        m0704(.A(mai_mai_n726_), .B(mai_mai_n628_), .Y(mai_mai_n727_));
  NA3        m0705(.A(mai_mai_n727_), .B(mai_mai_n725_), .C(mai_mai_n723_), .Y(mai_mai_n728_));
  NA3        m0706(.A(mai_mai_n728_), .B(mai_mai_n46_), .C(mai_mai_n226_), .Y(mai_mai_n729_));
  NA4        m0707(.A(mai_mai_n729_), .B(mai_mai_n721_), .C(mai_mai_n709_), .D(mai_mai_n693_), .Y(mai_mai_n730_));
  OR4        m0708(.A(mai_mai_n730_), .B(mai_mai_n684_), .C(mai_mai_n669_), .D(mai_mai_n610_), .Y(mai5));
  AOI210     m0709(.A0(mai_mai_n655_), .A1(mai_mai_n268_), .B0(mai_mai_n419_), .Y(mai_mai_n732_));
  AN2        m0710(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n733_));
  NA3        m0711(.A(mai_mai_n733_), .B(mai_mai_n722_), .C(mai_mai_n108_), .Y(mai_mai_n734_));
  NO2        m0712(.A(mai_mai_n592_), .B(i_11_), .Y(mai_mai_n735_));
  NA2        m0713(.A(mai_mai_n88_), .B(mai_mai_n735_), .Y(mai_mai_n736_));
  NA3        m0714(.A(mai_mai_n736_), .B(mai_mai_n734_), .C(mai_mai_n732_), .Y(mai_mai_n737_));
  NO3        m0715(.A(i_11_), .B(mai_mai_n238_), .C(i_13_), .Y(mai_mai_n738_));
  NO2        m0716(.A(mai_mai_n125_), .B(mai_mai_n23_), .Y(mai_mai_n739_));
  NA2        m0717(.A(i_12_), .B(i_8_), .Y(mai_mai_n740_));
  OAI210     m0718(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n740_), .Y(mai_mai_n741_));
  INV        m0719(.A(mai_mai_n446_), .Y(mai_mai_n742_));
  AOI220     m0720(.A0(mai_mai_n317_), .A1(mai_mai_n569_), .B0(mai_mai_n741_), .B1(mai_mai_n739_), .Y(mai_mai_n743_));
  INV        m0721(.A(mai_mai_n743_), .Y(mai_mai_n744_));
  NO2        m0722(.A(mai_mai_n744_), .B(mai_mai_n737_), .Y(mai_mai_n745_));
  INV        m0723(.A(mai_mai_n172_), .Y(mai_mai_n746_));
  INV        m0724(.A(mai_mai_n247_), .Y(mai_mai_n747_));
  OAI210     m0725(.A0(mai_mai_n680_), .A1(mai_mai_n448_), .B0(mai_mai_n111_), .Y(mai_mai_n748_));
  AOI210     m0726(.A0(mai_mai_n748_), .A1(mai_mai_n747_), .B0(mai_mai_n746_), .Y(mai_mai_n749_));
  NO2        m0727(.A(mai_mai_n456_), .B(mai_mai_n26_), .Y(mai_mai_n750_));
  NO2        m0728(.A(mai_mai_n750_), .B(mai_mai_n421_), .Y(mai_mai_n751_));
  NA2        m0729(.A(mai_mai_n751_), .B(i_2_), .Y(mai_mai_n752_));
  INV        m0730(.A(mai_mai_n752_), .Y(mai_mai_n753_));
  AOI210     m0731(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n417_), .Y(mai_mai_n754_));
  AOI210     m0732(.A0(mai_mai_n754_), .A1(mai_mai_n753_), .B0(mai_mai_n749_), .Y(mai_mai_n755_));
  NO2        m0733(.A(mai_mai_n192_), .B(mai_mai_n126_), .Y(mai_mai_n756_));
  OAI210     m0734(.A0(mai_mai_n756_), .A1(mai_mai_n739_), .B0(i_2_), .Y(mai_mai_n757_));
  INV        m0735(.A(mai_mai_n173_), .Y(mai_mai_n758_));
  NO3        m0736(.A(mai_mai_n612_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n759_));
  AOI210     m0737(.A0(mai_mai_n758_), .A1(mai_mai_n88_), .B0(mai_mai_n759_), .Y(mai_mai_n760_));
  AOI210     m0738(.A0(mai_mai_n760_), .A1(mai_mai_n757_), .B0(mai_mai_n195_), .Y(mai_mai_n761_));
  OA210      m0739(.A0(mai_mai_n613_), .A1(mai_mai_n127_), .B0(i_13_), .Y(mai_mai_n762_));
  NA2        m0740(.A(mai_mai_n201_), .B(mai_mai_n204_), .Y(mai_mai_n763_));
  NA2        m0741(.A(mai_mai_n151_), .B(mai_mai_n588_), .Y(mai_mai_n764_));
  AOI210     m0742(.A0(mai_mai_n764_), .A1(mai_mai_n763_), .B0(mai_mai_n373_), .Y(mai_mai_n765_));
  AOI210     m0743(.A0(mai_mai_n209_), .A1(mai_mai_n148_), .B0(mai_mai_n513_), .Y(mai_mai_n766_));
  NA2        m0744(.A(mai_mai_n766_), .B(mai_mai_n421_), .Y(mai_mai_n767_));
  NO2        m0745(.A(mai_mai_n102_), .B(mai_mai_n45_), .Y(mai_mai_n768_));
  INV        m0746(.A(mai_mai_n301_), .Y(mai_mai_n769_));
  NA4        m0747(.A(mai_mai_n769_), .B(mai_mai_n305_), .C(mai_mai_n125_), .D(mai_mai_n43_), .Y(mai_mai_n770_));
  OAI210     m0748(.A0(mai_mai_n770_), .A1(mai_mai_n768_), .B0(mai_mai_n767_), .Y(mai_mai_n771_));
  NO4        m0749(.A(mai_mai_n771_), .B(mai_mai_n765_), .C(mai_mai_n762_), .D(mai_mai_n761_), .Y(mai_mai_n772_));
  NA2        m0750(.A(mai_mai_n569_), .B(mai_mai_n28_), .Y(mai_mai_n773_));
  NA2        m0751(.A(mai_mai_n738_), .B(mai_mai_n275_), .Y(mai_mai_n774_));
  NA2        m0752(.A(mai_mai_n774_), .B(mai_mai_n773_), .Y(mai_mai_n775_));
  NO2        m0753(.A(mai_mai_n62_), .B(i_12_), .Y(mai_mai_n776_));
  NO2        m0754(.A(mai_mai_n776_), .B(mai_mai_n127_), .Y(mai_mai_n777_));
  NO2        m0755(.A(mai_mai_n777_), .B(mai_mai_n588_), .Y(mai_mai_n778_));
  AOI220     m0756(.A0(mai_mai_n778_), .A1(mai_mai_n36_), .B0(mai_mai_n775_), .B1(mai_mai_n47_), .Y(mai_mai_n779_));
  NA4        m0757(.A(mai_mai_n779_), .B(mai_mai_n772_), .C(mai_mai_n755_), .D(mai_mai_n745_), .Y(mai6));
  NO3        m0758(.A(i_9_), .B(mai_mai_n307_), .C(i_1_), .Y(mai_mai_n781_));
  NO2        m0759(.A(mai_mai_n187_), .B(mai_mai_n139_), .Y(mai_mai_n782_));
  OAI210     m0760(.A0(mai_mai_n782_), .A1(mai_mai_n781_), .B0(mai_mai_n726_), .Y(mai_mai_n783_));
  NA4        m0761(.A(mai_mai_n388_), .B(mai_mai_n483_), .C(mai_mai_n71_), .D(mai_mai_n101_), .Y(mai_mai_n784_));
  INV        m0762(.A(mai_mai_n784_), .Y(mai_mai_n785_));
  NO2        m0763(.A(i_11_), .B(i_9_), .Y(mai_mai_n786_));
  NO2        m0764(.A(mai_mai_n785_), .B(mai_mai_n328_), .Y(mai_mai_n787_));
  AO210      m0765(.A0(mai_mai_n787_), .A1(mai_mai_n783_), .B0(i_12_), .Y(mai_mai_n788_));
  NA2        m0766(.A(mai_mai_n374_), .B(mai_mai_n335_), .Y(mai_mai_n789_));
  NA2        m0767(.A(mai_mai_n576_), .B(mai_mai_n63_), .Y(mai_mai_n790_));
  NA2        m0768(.A(mai_mai_n671_), .B(mai_mai_n71_), .Y(mai_mai_n791_));
  BUFFER     m0769(.A(mai_mai_n618_), .Y(mai_mai_n792_));
  NA4        m0770(.A(mai_mai_n792_), .B(mai_mai_n791_), .C(mai_mai_n790_), .D(mai_mai_n789_), .Y(mai_mai_n793_));
  INV        m0771(.A(mai_mai_n198_), .Y(mai_mai_n794_));
  AOI220     m0772(.A0(mai_mai_n794_), .A1(mai_mai_n786_), .B0(mai_mai_n793_), .B1(mai_mai_n73_), .Y(mai_mai_n795_));
  INV        m0773(.A(mai_mai_n327_), .Y(mai_mai_n796_));
  NA2        m0774(.A(mai_mai_n75_), .B(mai_mai_n132_), .Y(mai_mai_n797_));
  INV        m0775(.A(mai_mai_n125_), .Y(mai_mai_n798_));
  NA2        m0776(.A(mai_mai_n798_), .B(mai_mai_n47_), .Y(mai_mai_n799_));
  AOI210     m0777(.A0(mai_mai_n799_), .A1(mai_mai_n797_), .B0(mai_mai_n796_), .Y(mai_mai_n800_));
  NO2        m0778(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n801_));
  NA3        m0779(.A(mai_mai_n801_), .B(mai_mai_n474_), .C(mai_mai_n388_), .Y(mai_mai_n802_));
  NAi32      m0780(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n803_));
  AOI210     m0781(.A0(mai_mai_n710_), .A1(mai_mai_n86_), .B0(mai_mai_n803_), .Y(mai_mai_n804_));
  OAI210     m0782(.A0(mai_mai_n670_), .A1(mai_mai_n557_), .B0(mai_mai_n556_), .Y(mai_mai_n805_));
  NAi31      m0783(.An(mai_mai_n804_), .B(mai_mai_n805_), .C(mai_mai_n802_), .Y(mai_mai_n806_));
  OR2        m0784(.A(mai_mai_n806_), .B(mai_mai_n800_), .Y(mai_mai_n807_));
  NO2        m0785(.A(mai_mai_n685_), .B(i_2_), .Y(mai_mai_n808_));
  NA2        m0786(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n809_));
  OAI210     m0787(.A0(mai_mai_n809_), .A1(mai_mai_n409_), .B0(mai_mai_n361_), .Y(mai_mai_n810_));
  NA2        m0788(.A(mai_mai_n810_), .B(mai_mai_n808_), .Y(mai_mai_n811_));
  AO210      m0789(.A0(mai_mai_n360_), .A1(mai_mai_n351_), .B0(mai_mai_n395_), .Y(mai_mai_n812_));
  NA3        m0790(.A(mai_mai_n812_), .B(mai_mai_n256_), .C(i_7_), .Y(mai_mai_n813_));
  OR2        m0791(.A(mai_mai_n613_), .B(mai_mai_n448_), .Y(mai_mai_n814_));
  NA3        m0792(.A(mai_mai_n814_), .B(mai_mai_n147_), .C(mai_mai_n69_), .Y(mai_mai_n815_));
  OR2        m0793(.A(mai_mai_n742_), .B(mai_mai_n36_), .Y(mai_mai_n816_));
  NA4        m0794(.A(mai_mai_n816_), .B(mai_mai_n815_), .C(mai_mai_n813_), .D(mai_mai_n811_), .Y(mai_mai_n817_));
  OAI210     m0795(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n86_), .Y(mai_mai_n818_));
  NA2        m0796(.A(mai_mai_n818_), .B(mai_mai_n556_), .Y(mai_mai_n819_));
  NA2        m0797(.A(mai_mai_n395_), .B(mai_mai_n70_), .Y(mai_mai_n820_));
  NA3        m0798(.A(mai_mai_n820_), .B(mai_mai_n819_), .C(mai_mai_n595_), .Y(mai_mai_n821_));
  AO210      m0799(.A0(mai_mai_n513_), .A1(mai_mai_n47_), .B0(mai_mai_n87_), .Y(mai_mai_n822_));
  NA3        m0800(.A(mai_mai_n822_), .B(mai_mai_n484_), .C(mai_mai_n219_), .Y(mai_mai_n823_));
  AOI210     m0801(.A0(mai_mai_n448_), .A1(mai_mai_n446_), .B0(mai_mai_n555_), .Y(mai_mai_n824_));
  NA2        m0802(.A(mai_mai_n112_), .B(mai_mai_n408_), .Y(mai_mai_n825_));
  NA2        m0803(.A(mai_mai_n246_), .B(mai_mai_n47_), .Y(mai_mai_n826_));
  NA3        m0804(.A(mai_mai_n825_), .B(mai_mai_n824_), .C(mai_mai_n823_), .Y(mai_mai_n827_));
  NO4        m0805(.A(mai_mai_n827_), .B(mai_mai_n821_), .C(mai_mai_n817_), .D(mai_mai_n807_), .Y(mai_mai_n828_));
  NA4        m0806(.A(mai_mai_n828_), .B(mai_mai_n795_), .C(mai_mai_n788_), .D(mai_mai_n379_), .Y(mai3));
  NA2        m0807(.A(i_6_), .B(i_7_), .Y(mai_mai_n830_));
  NO2        m0808(.A(mai_mai_n830_), .B(i_0_), .Y(mai_mai_n831_));
  NO2        m0809(.A(i_11_), .B(mai_mai_n238_), .Y(mai_mai_n832_));
  OAI210     m0810(.A0(mai_mai_n831_), .A1(mai_mai_n289_), .B0(mai_mai_n832_), .Y(mai_mai_n833_));
  NO2        m0811(.A(mai_mai_n833_), .B(mai_mai_n195_), .Y(mai_mai_n834_));
  NO3        m0812(.A(mai_mai_n452_), .B(mai_mai_n89_), .C(mai_mai_n45_), .Y(mai_mai_n835_));
  OA210      m0813(.A0(mai_mai_n835_), .A1(mai_mai_n834_), .B0(mai_mai_n175_), .Y(mai_mai_n836_));
  NA2        m0814(.A(mai_mai_n410_), .B(mai_mai_n46_), .Y(mai_mai_n837_));
  NO4        m0815(.A(mai_mai_n375_), .B(mai_mai_n382_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n838_));
  INV        m0816(.A(mai_mai_n838_), .Y(mai_mai_n839_));
  NA2        m0817(.A(mai_mai_n697_), .B(mai_mai_n663_), .Y(mai_mai_n840_));
  NA2        m0818(.A(mai_mai_n333_), .B(mai_mai_n438_), .Y(mai_mai_n841_));
  OAI220     m0819(.A0(mai_mai_n841_), .A1(mai_mai_n840_), .B0(mai_mai_n839_), .B1(mai_mai_n63_), .Y(mai_mai_n842_));
  NOi21      m0820(.An(i_5_), .B(i_9_), .Y(mai_mai_n843_));
  NA2        m0821(.A(mai_mai_n843_), .B(mai_mai_n445_), .Y(mai_mai_n844_));
  AOI210     m0822(.A0(mai_mai_n265_), .A1(mai_mai_n476_), .B0(mai_mai_n674_), .Y(mai_mai_n845_));
  NO3        m0823(.A(mai_mai_n413_), .B(mai_mai_n265_), .C(mai_mai_n73_), .Y(mai_mai_n846_));
  NO2        m0824(.A(mai_mai_n176_), .B(mai_mai_n148_), .Y(mai_mai_n847_));
  AOI210     m0825(.A0(mai_mai_n847_), .A1(mai_mai_n246_), .B0(mai_mai_n846_), .Y(mai_mai_n848_));
  OAI220     m0826(.A0(mai_mai_n848_), .A1(mai_mai_n182_), .B0(mai_mai_n845_), .B1(mai_mai_n844_), .Y(mai_mai_n849_));
  NO3        m0827(.A(mai_mai_n849_), .B(mai_mai_n842_), .C(mai_mai_n836_), .Y(mai_mai_n850_));
  NA2        m0828(.A(mai_mai_n187_), .B(mai_mai_n24_), .Y(mai_mai_n851_));
  NO2        m0829(.A(mai_mai_n661_), .B(mai_mai_n586_), .Y(mai_mai_n852_));
  NO2        m0830(.A(mai_mai_n852_), .B(mai_mai_n851_), .Y(mai_mai_n853_));
  NA2        m0831(.A(mai_mai_n312_), .B(mai_mai_n130_), .Y(mai_mai_n854_));
  NAi21      m0832(.An(mai_mai_n162_), .B(mai_mai_n438_), .Y(mai_mai_n855_));
  OAI220     m0833(.A0(mai_mai_n855_), .A1(mai_mai_n826_), .B0(mai_mai_n854_), .B1(mai_mai_n400_), .Y(mai_mai_n856_));
  NO2        m0834(.A(mai_mai_n856_), .B(mai_mai_n853_), .Y(mai_mai_n857_));
  NO2        m0835(.A(mai_mai_n388_), .B(mai_mai_n293_), .Y(mai_mai_n858_));
  NA2        m0836(.A(mai_mai_n858_), .B(mai_mai_n699_), .Y(mai_mai_n859_));
  NA2        m0837(.A(mai_mai_n566_), .B(i_0_), .Y(mai_mai_n860_));
  NO3        m0838(.A(mai_mai_n860_), .B(mai_mai_n383_), .C(mai_mai_n88_), .Y(mai_mai_n861_));
  INV        m0839(.A(mai_mai_n861_), .Y(mai_mai_n862_));
  AN2        m0840(.A(mai_mai_n96_), .B(mai_mai_n245_), .Y(mai_mai_n863_));
  NA2        m0841(.A(mai_mai_n738_), .B(mai_mai_n328_), .Y(mai_mai_n864_));
  INV        m0842(.A(mai_mai_n58_), .Y(mai_mai_n865_));
  OAI220     m0843(.A0(mai_mai_n865_), .A1(mai_mai_n864_), .B0(mai_mai_n650_), .B1(mai_mai_n531_), .Y(mai_mai_n866_));
  NA2        m0844(.A(i_0_), .B(i_10_), .Y(mai_mai_n867_));
  NA2        m0845(.A(mai_mai_n187_), .B(mai_mai_n84_), .Y(mai_mai_n868_));
  NA2        m0846(.A(mai_mai_n560_), .B(i_4_), .Y(mai_mai_n869_));
  NA2        m0847(.A(mai_mai_n190_), .B(mai_mai_n204_), .Y(mai_mai_n870_));
  OAI220     m0848(.A0(mai_mai_n870_), .A1(mai_mai_n864_), .B0(mai_mai_n869_), .B1(mai_mai_n868_), .Y(mai_mai_n871_));
  NO3        m0849(.A(mai_mai_n871_), .B(mai_mai_n866_), .C(mai_mai_n863_), .Y(mai_mai_n872_));
  NA4        m0850(.A(mai_mai_n872_), .B(mai_mai_n862_), .C(mai_mai_n859_), .D(mai_mai_n857_), .Y(mai_mai_n873_));
  NA2        m0851(.A(i_11_), .B(i_9_), .Y(mai_mai_n874_));
  NO2        m0852(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n875_));
  NA2        m0853(.A(mai_mai_n393_), .B(mai_mai_n180_), .Y(mai_mai_n876_));
  NA2        m0854(.A(mai_mai_n876_), .B(mai_mai_n160_), .Y(mai_mai_n877_));
  NO2        m0855(.A(mai_mai_n874_), .B(mai_mai_n73_), .Y(mai_mai_n878_));
  NO2        m0856(.A(mai_mai_n176_), .B(i_0_), .Y(mai_mai_n879_));
  INV        m0857(.A(mai_mai_n879_), .Y(mai_mai_n880_));
  NA2        m0858(.A(mai_mai_n474_), .B(mai_mai_n232_), .Y(mai_mai_n881_));
  NO2        m0859(.A(mai_mai_n881_), .B(mai_mai_n880_), .Y(mai_mai_n882_));
  NO2        m0860(.A(mai_mai_n882_), .B(mai_mai_n877_), .Y(mai_mai_n883_));
  NA2        m0861(.A(mai_mai_n649_), .B(mai_mai_n122_), .Y(mai_mai_n884_));
  NO2        m0862(.A(i_6_), .B(mai_mai_n884_), .Y(mai_mai_n885_));
  AOI210     m0863(.A0(mai_mai_n447_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n886_));
  NA2        m0864(.A(mai_mai_n172_), .B(mai_mai_n103_), .Y(mai_mai_n887_));
  NOi32      m0865(.An(mai_mai_n886_), .Bn(mai_mai_n190_), .C(mai_mai_n887_), .Y(mai_mai_n888_));
  NA2        m0866(.A(mai_mai_n596_), .B(mai_mai_n328_), .Y(mai_mai_n889_));
  NO2        m0867(.A(mai_mai_n889_), .B(mai_mai_n837_), .Y(mai_mai_n890_));
  NO3        m0868(.A(mai_mai_n890_), .B(mai_mai_n888_), .C(mai_mai_n885_), .Y(mai_mai_n891_));
  NOi21      m0869(.An(i_7_), .B(i_5_), .Y(mai_mai_n892_));
  NOi31      m0870(.An(mai_mai_n892_), .B(i_0_), .C(mai_mai_n716_), .Y(mai_mai_n893_));
  NA3        m0871(.A(mai_mai_n893_), .B(i_3_), .C(i_6_), .Y(mai_mai_n894_));
  BUFFER     m0872(.A(mai_mai_n894_), .Y(mai_mai_n895_));
  NO3        m0873(.A(mai_mai_n403_), .B(mai_mai_n363_), .C(mai_mai_n359_), .Y(mai_mai_n896_));
  NO2        m0874(.A(mai_mai_n259_), .B(mai_mai_n318_), .Y(mai_mai_n897_));
  INV        m0875(.A(mai_mai_n716_), .Y(mai_mai_n898_));
  AOI210     m0876(.A0(mai_mai_n898_), .A1(mai_mai_n897_), .B0(mai_mai_n896_), .Y(mai_mai_n899_));
  NA4        m0877(.A(mai_mai_n899_), .B(mai_mai_n895_), .C(mai_mai_n891_), .D(mai_mai_n883_), .Y(mai_mai_n900_));
  NO2        m0878(.A(mai_mai_n851_), .B(mai_mai_n241_), .Y(mai_mai_n901_));
  AN2        m0879(.A(mai_mai_n332_), .B(mai_mai_n328_), .Y(mai_mai_n902_));
  AN2        m0880(.A(mai_mai_n902_), .B(mai_mai_n847_), .Y(mai_mai_n903_));
  OAI210     m0881(.A0(mai_mai_n903_), .A1(mai_mai_n901_), .B0(i_10_), .Y(mai_mai_n904_));
  OA210      m0882(.A0(mai_mai_n474_), .A1(mai_mai_n224_), .B0(mai_mai_n473_), .Y(mai_mai_n905_));
  NA3        m0883(.A(mai_mai_n473_), .B(mai_mai_n410_), .C(mai_mai_n46_), .Y(mai_mai_n906_));
  OAI210     m0884(.A0(mai_mai_n855_), .A1(i_6_), .B0(mai_mai_n906_), .Y(mai_mai_n907_));
  NA2        m0885(.A(mai_mai_n878_), .B(mai_mai_n305_), .Y(mai_mai_n908_));
  NA2        m0886(.A(mai_mai_n189_), .B(mai_mai_n908_), .Y(mai_mai_n909_));
  AOI220     m0887(.A0(mai_mai_n909_), .A1(mai_mai_n474_), .B0(mai_mai_n907_), .B1(mai_mai_n73_), .Y(mai_mai_n910_));
  NO2        m0888(.A(mai_mai_n75_), .B(mai_mai_n740_), .Y(mai_mai_n911_));
  AOI220     m0889(.A0(mai_mai_n911_), .A1(i_11_), .B0(mai_mai_n175_), .B1(mai_mai_n586_), .Y(mai_mai_n912_));
  NO2        m0890(.A(mai_mai_n912_), .B(mai_mai_n48_), .Y(mai_mai_n913_));
  NO3        m0891(.A(i_5_), .B(mai_mai_n358_), .C(mai_mai_n24_), .Y(mai_mai_n914_));
  INV        m0892(.A(mai_mai_n914_), .Y(mai_mai_n915_));
  NAi21      m0893(.An(i_9_), .B(i_5_), .Y(mai_mai_n916_));
  NO2        m0894(.A(mai_mai_n590_), .B(mai_mai_n105_), .Y(mai_mai_n917_));
  NA2        m0895(.A(mai_mai_n917_), .B(i_0_), .Y(mai_mai_n918_));
  OAI220     m0896(.A0(mai_mai_n918_), .A1(mai_mai_n85_), .B0(mai_mai_n915_), .B1(mai_mai_n173_), .Y(mai_mai_n919_));
  NO2        m0897(.A(mai_mai_n919_), .B(mai_mai_n913_), .Y(mai_mai_n920_));
  NA3        m0898(.A(mai_mai_n920_), .B(mai_mai_n910_), .C(mai_mai_n904_), .Y(mai_mai_n921_));
  NO3        m0899(.A(mai_mai_n921_), .B(mai_mai_n900_), .C(mai_mai_n873_), .Y(mai_mai_n922_));
  NO2        m0900(.A(i_0_), .B(mai_mai_n716_), .Y(mai_mai_n923_));
  NA2        m0901(.A(mai_mai_n73_), .B(mai_mai_n45_), .Y(mai_mai_n924_));
  NO2        m0902(.A(mai_mai_n790_), .B(mai_mai_n887_), .Y(mai_mai_n925_));
  INV        m0903(.A(mai_mai_n925_), .Y(mai_mai_n926_));
  NA2        m0904(.A(mai_mai_n726_), .B(mai_mai_n146_), .Y(mai_mai_n927_));
  INV        m0905(.A(mai_mai_n927_), .Y(mai_mai_n928_));
  NA3        m0906(.A(mai_mai_n928_), .B(mai_mai_n663_), .C(mai_mai_n73_), .Y(mai_mai_n929_));
  NO2        m0907(.A(mai_mai_n805_), .B(mai_mai_n403_), .Y(mai_mai_n930_));
  NA2        m0908(.A(mai_mai_n246_), .B(mai_mai_n231_), .Y(mai_mai_n931_));
  AOI210     m0909(.A0(mai_mai_n931_), .A1(mai_mai_n860_), .B0(mai_mai_n153_), .Y(mai_mai_n932_));
  NO2        m0910(.A(mai_mai_n932_), .B(mai_mai_n930_), .Y(mai_mai_n933_));
  NA3        m0911(.A(mai_mai_n933_), .B(mai_mai_n929_), .C(mai_mai_n926_), .Y(mai_mai_n934_));
  NA2        m0912(.A(mai_mai_n902_), .B(mai_mai_n373_), .Y(mai_mai_n935_));
  AOI210     m0913(.A0(mai_mai_n300_), .A1(mai_mai_n162_), .B0(mai_mai_n935_), .Y(mai_mai_n936_));
  NA3        m0914(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n937_));
  NA2        m0915(.A(mai_mai_n875_), .B(mai_mai_n488_), .Y(mai_mai_n938_));
  AOI210     m0916(.A0(mai_mai_n937_), .A1(mai_mai_n162_), .B0(mai_mai_n938_), .Y(mai_mai_n939_));
  NO2        m0917(.A(mai_mai_n939_), .B(mai_mai_n936_), .Y(mai_mai_n940_));
  NO3        m0918(.A(mai_mai_n867_), .B(mai_mai_n843_), .C(mai_mai_n192_), .Y(mai_mai_n941_));
  AOI220     m0919(.A0(mai_mai_n941_), .A1(i_11_), .B0(mai_mai_n561_), .B1(mai_mai_n75_), .Y(mai_mai_n942_));
  NO3        m0920(.A(mai_mai_n210_), .B(mai_mai_n382_), .C(i_0_), .Y(mai_mai_n943_));
  OAI210     m0921(.A0(mai_mai_n943_), .A1(mai_mai_n76_), .B0(i_13_), .Y(mai_mai_n944_));
  INV        m0922(.A(mai_mai_n219_), .Y(mai_mai_n945_));
  NO2        m0923(.A(mai_mai_n524_), .B(mai_mai_n139_), .Y(mai_mai_n946_));
  NA3        m0924(.A(mai_mai_n946_), .B(i_7_), .C(mai_mai_n945_), .Y(mai_mai_n947_));
  NA4        m0925(.A(mai_mai_n947_), .B(mai_mai_n944_), .C(mai_mai_n942_), .D(mai_mai_n940_), .Y(mai_mai_n948_));
  INV        m0926(.A(mai_mai_n92_), .Y(mai_mai_n949_));
  AOI210     m0927(.A0(mai_mai_n949_), .A1(mai_mai_n923_), .B0(mai_mai_n109_), .Y(mai_mai_n950_));
  AOI220     m0928(.A0(mai_mai_n892_), .A1(mai_mai_n488_), .B0(mai_mai_n831_), .B1(mai_mai_n163_), .Y(mai_mai_n951_));
  NA2        m0929(.A(mai_mai_n351_), .B(mai_mai_n177_), .Y(mai_mai_n952_));
  OA220      m0930(.A0(mai_mai_n952_), .A1(mai_mai_n951_), .B0(mai_mai_n950_), .B1(i_5_), .Y(mai_mai_n953_));
  AOI210     m0931(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n176_), .Y(mai_mai_n954_));
  NA2        m0932(.A(mai_mai_n954_), .B(mai_mai_n905_), .Y(mai_mai_n955_));
  NO3        m0933(.A(mai_mai_n837_), .B(mai_mai_n55_), .C(mai_mai_n49_), .Y(mai_mai_n956_));
  NA2        m0934(.A(mai_mai_n493_), .B(mai_mai_n471_), .Y(mai_mai_n957_));
  NO2        m0935(.A(mai_mai_n957_), .B(mai_mai_n956_), .Y(mai_mai_n958_));
  NA3        m0936(.A(mai_mai_n388_), .B(mai_mai_n172_), .C(mai_mai_n171_), .Y(mai_mai_n959_));
  NA3        m0937(.A(mai_mai_n875_), .B(mai_mai_n289_), .C(mai_mai_n231_), .Y(mai_mai_n960_));
  NA2        m0938(.A(mai_mai_n960_), .B(mai_mai_n959_), .Y(mai_mai_n961_));
  NA3        m0939(.A(mai_mai_n388_), .B(mai_mai_n334_), .C(mai_mai_n222_), .Y(mai_mai_n962_));
  INV        m0940(.A(mai_mai_n962_), .Y(mai_mai_n963_));
  NOi31      m0941(.An(mai_mai_n387_), .B(mai_mai_n924_), .C(mai_mai_n241_), .Y(mai_mai_n964_));
  NO3        m0942(.A(mai_mai_n874_), .B(mai_mai_n219_), .C(mai_mai_n192_), .Y(mai_mai_n965_));
  NO4        m0943(.A(mai_mai_n965_), .B(mai_mai_n964_), .C(mai_mai_n963_), .D(mai_mai_n961_), .Y(mai_mai_n966_));
  NA4        m0944(.A(mai_mai_n966_), .B(mai_mai_n958_), .C(mai_mai_n955_), .D(mai_mai_n953_), .Y(mai_mai_n967_));
  NA2        m0945(.A(mai_mai_n305_), .B(i_5_), .Y(mai_mai_n968_));
  NA2        m0946(.A(mai_mai_n968_), .B(mai_mai_n244_), .Y(mai_mai_n969_));
  NO4        m0947(.A(mai_mai_n241_), .B(mai_mai_n210_), .C(i_0_), .D(i_12_), .Y(mai_mai_n970_));
  AOI220     m0948(.A0(mai_mai_n970_), .A1(mai_mai_n969_), .B0(mai_mai_n785_), .B1(mai_mai_n177_), .Y(mai_mai_n971_));
  AN2        m0949(.A(mai_mai_n867_), .B(mai_mai_n153_), .Y(mai_mai_n972_));
  NO4        m0950(.A(mai_mai_n972_), .B(i_12_), .C(mai_mai_n637_), .D(mai_mai_n132_), .Y(mai_mai_n973_));
  NA2        m0951(.A(mai_mai_n973_), .B(mai_mai_n219_), .Y(mai_mai_n974_));
  NA3        m0952(.A(mai_mai_n98_), .B(mai_mai_n565_), .C(i_11_), .Y(mai_mai_n975_));
  NO2        m0953(.A(mai_mai_n975_), .B(mai_mai_n155_), .Y(mai_mai_n976_));
  NA2        m0954(.A(mai_mai_n892_), .B(mai_mai_n470_), .Y(mai_mai_n977_));
  NA2        m0955(.A(mai_mai_n64_), .B(mai_mai_n101_), .Y(mai_mai_n978_));
  OAI220     m0956(.A0(mai_mai_n978_), .A1(mai_mai_n968_), .B0(mai_mai_n977_), .B1(mai_mai_n664_), .Y(mai_mai_n979_));
  AOI210     m0957(.A0(mai_mai_n979_), .A1(mai_mai_n879_), .B0(mai_mai_n976_), .Y(mai_mai_n980_));
  NA3        m0958(.A(mai_mai_n980_), .B(mai_mai_n974_), .C(mai_mai_n971_), .Y(mai_mai_n981_));
  NO4        m0959(.A(mai_mai_n981_), .B(mai_mai_n967_), .C(mai_mai_n948_), .D(mai_mai_n934_), .Y(mai_mai_n982_));
  OAI210     m0960(.A0(mai_mai_n808_), .A1(mai_mai_n801_), .B0(mai_mai_n37_), .Y(mai_mai_n983_));
  NA3        m0961(.A(mai_mai_n886_), .B(mai_mai_n371_), .C(i_5_), .Y(mai_mai_n984_));
  NA3        m0962(.A(mai_mai_n984_), .B(mai_mai_n983_), .C(mai_mai_n602_), .Y(mai_mai_n985_));
  NA2        m0963(.A(mai_mai_n985_), .B(mai_mai_n207_), .Y(mai_mai_n986_));
  NA2        m0964(.A(mai_mai_n188_), .B(mai_mai_n190_), .Y(mai_mai_n987_));
  AO210      m0965(.A0(i_11_), .A1(mai_mai_n33_), .B0(mai_mai_n987_), .Y(mai_mai_n988_));
  OAI210     m0966(.A0(mai_mai_n606_), .A1(mai_mai_n604_), .B0(mai_mai_n317_), .Y(mai_mai_n989_));
  NA2        m0967(.A(mai_mai_n989_), .B(mai_mai_n988_), .Y(mai_mai_n990_));
  NO2        m0968(.A(mai_mai_n461_), .B(mai_mai_n265_), .Y(mai_mai_n991_));
  NO4        m0969(.A(mai_mai_n234_), .B(mai_mai_n145_), .C(mai_mai_n667_), .D(mai_mai_n37_), .Y(mai_mai_n992_));
  NO2        m0970(.A(mai_mai_n992_), .B(mai_mai_n991_), .Y(mai_mai_n993_));
  OAI210     m0971(.A0(mai_mai_n975_), .A1(mai_mai_n148_), .B0(mai_mai_n993_), .Y(mai_mai_n994_));
  AOI210     m0972(.A0(mai_mai_n990_), .A1(mai_mai_n49_), .B0(mai_mai_n994_), .Y(mai_mai_n995_));
  AOI210     m0973(.A0(mai_mai_n995_), .A1(mai_mai_n986_), .B0(mai_mai_n73_), .Y(mai_mai_n996_));
  NO2        m0974(.A(mai_mai_n558_), .B(mai_mai_n378_), .Y(mai_mai_n997_));
  NO2        m0975(.A(mai_mai_n997_), .B(mai_mai_n746_), .Y(mai_mai_n998_));
  INV        m0976(.A(mai_mai_n76_), .Y(mai_mai_n999_));
  AOI210     m0977(.A0(mai_mai_n954_), .A1(mai_mai_n875_), .B0(mai_mai_n893_), .Y(mai_mai_n1000_));
  AOI210     m0978(.A0(mai_mai_n1000_), .A1(mai_mai_n999_), .B0(mai_mai_n667_), .Y(mai_mai_n1001_));
  NA2        m0979(.A(mai_mai_n259_), .B(mai_mai_n57_), .Y(mai_mai_n1002_));
  NA2        m0980(.A(mai_mai_n1002_), .B(mai_mai_n76_), .Y(mai_mai_n1003_));
  NO2        m0981(.A(mai_mai_n1003_), .B(mai_mai_n238_), .Y(mai_mai_n1004_));
  NA3        m0982(.A(mai_mai_n96_), .B(mai_mai_n307_), .C(mai_mai_n31_), .Y(mai_mai_n1005_));
  INV        m0983(.A(mai_mai_n1005_), .Y(mai_mai_n1006_));
  NO3        m0984(.A(mai_mai_n1006_), .B(mai_mai_n1004_), .C(mai_mai_n1001_), .Y(mai_mai_n1007_));
  OAI210     m0985(.A0(mai_mai_n267_), .A1(mai_mai_n158_), .B0(mai_mai_n88_), .Y(mai_mai_n1008_));
  NA3        m0986(.A(mai_mai_n750_), .B(mai_mai_n289_), .C(mai_mai_n80_), .Y(mai_mai_n1009_));
  AOI210     m0987(.A0(mai_mai_n1009_), .A1(mai_mai_n1008_), .B0(i_11_), .Y(mai_mai_n1010_));
  OAI210     m0988(.A0(mai_mai_n1025_), .A1(mai_mai_n886_), .B0(mai_mai_n207_), .Y(mai_mai_n1011_));
  NA2        m0989(.A(mai_mai_n164_), .B(i_5_), .Y(mai_mai_n1012_));
  AOI210     m0990(.A0(mai_mai_n1011_), .A1(mai_mai_n763_), .B0(mai_mai_n1012_), .Y(mai_mai_n1013_));
  NO4        m0991(.A(mai_mai_n916_), .B(mai_mai_n477_), .C(mai_mai_n255_), .D(mai_mai_n254_), .Y(mai_mai_n1014_));
  NO2        m0992(.A(mai_mai_n1014_), .B(mai_mai_n555_), .Y(mai_mai_n1015_));
  INV        m0993(.A(mai_mai_n364_), .Y(mai_mai_n1016_));
  AOI210     m0994(.A0(mai_mai_n1016_), .A1(mai_mai_n1015_), .B0(mai_mai_n41_), .Y(mai_mai_n1017_));
  NO3        m0995(.A(mai_mai_n1017_), .B(mai_mai_n1013_), .C(mai_mai_n1010_), .Y(mai_mai_n1018_));
  OAI210     m0996(.A0(mai_mai_n1007_), .A1(i_4_), .B0(mai_mai_n1018_), .Y(mai_mai_n1019_));
  NO3        m0997(.A(mai_mai_n1019_), .B(mai_mai_n998_), .C(mai_mai_n996_), .Y(mai_mai_n1020_));
  NA4        m0998(.A(mai_mai_n1020_), .B(mai_mai_n982_), .C(mai_mai_n922_), .D(mai_mai_n850_), .Y(mai4));
  INV        m0999(.A(i_2_), .Y(mai_mai_n1024_));
  INV        m1000(.A(i_12_), .Y(mai_mai_n1025_));
  INV        m1001(.A(i_12_), .Y(mai_mai_n1026_));
  INV        m1002(.A(mai_mai_n82_), .Y(mai_mai_n1027_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  NA2        u0029(.A(i_0_), .B(i_2_), .Y(men_men_n52_));
  NA2        u0030(.A(i_7_), .B(i_9_), .Y(men_men_n53_));
  NO2        u0031(.A(men_men_n53_), .B(men_men_n52_), .Y(men_men_n54_));
  NA3        u0032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n55_));
  NO2        u0033(.A(i_1_), .B(i_6_), .Y(men_men_n56_));
  NA2        u0034(.A(i_8_), .B(i_7_), .Y(men_men_n57_));
  INV        u0035(.A(men_men_n55_), .Y(men_men_n58_));
  NA2        u0036(.A(men_men_n58_), .B(i_12_), .Y(men_men_n59_));
  NAi21      u0037(.An(i_2_), .B(i_7_), .Y(men_men_n60_));
  INV        u0038(.A(i_1_), .Y(men_men_n61_));
  NA2        u0039(.A(men_men_n61_), .B(i_6_), .Y(men_men_n62_));
  NA3        u0040(.A(men_men_n62_), .B(men_men_n60_), .C(men_men_n31_), .Y(men_men_n63_));
  NA2        u0041(.A(i_1_), .B(i_10_), .Y(men_men_n64_));
  NO2        u0042(.A(men_men_n64_), .B(i_6_), .Y(men_men_n65_));
  NAi31      u0043(.An(men_men_n65_), .B(men_men_n63_), .C(men_men_n59_), .Y(men_men_n66_));
  NA2        u0044(.A(men_men_n51_), .B(i_2_), .Y(men_men_n67_));
  AOI210     u0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n68_));
  NA2        u0046(.A(i_1_), .B(i_6_), .Y(men_men_n69_));
  NO2        u0047(.A(men_men_n69_), .B(men_men_n25_), .Y(men_men_n70_));
  INV        u0048(.A(i_0_), .Y(men_men_n71_));
  NAi21      u0049(.An(i_5_), .B(i_10_), .Y(men_men_n72_));
  NA2        u0050(.A(i_5_), .B(i_9_), .Y(men_men_n73_));
  AOI210     u0051(.A0(men_men_n73_), .A1(men_men_n72_), .B0(men_men_n71_), .Y(men_men_n74_));
  NO2        u0052(.A(men_men_n74_), .B(men_men_n70_), .Y(men_men_n75_));
  OAI210     u0053(.A0(men_men_n68_), .A1(men_men_n67_), .B0(men_men_n75_), .Y(men_men_n76_));
  OAI210     u0054(.A0(men_men_n76_), .A1(men_men_n66_), .B0(i_0_), .Y(men_men_n77_));
  NA2        u0055(.A(i_12_), .B(i_5_), .Y(men_men_n78_));
  NA2        u0056(.A(i_2_), .B(i_8_), .Y(men_men_n79_));
  NO2        u0057(.A(i_3_), .B(i_9_), .Y(men_men_n80_));
  NO2        u0058(.A(i_3_), .B(i_7_), .Y(men_men_n81_));
  NO3        u0059(.A(men_men_n81_), .B(men_men_n80_), .C(men_men_n61_), .Y(men_men_n82_));
  INV        u0060(.A(i_6_), .Y(men_men_n83_));
  OR4        u0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n84_));
  INV        u0062(.A(men_men_n84_), .Y(men_men_n85_));
  NO2        u0063(.A(i_2_), .B(i_7_), .Y(men_men_n86_));
  NO2        u0064(.A(men_men_n85_), .B(men_men_n86_), .Y(men_men_n87_));
  NA2        u0065(.A(men_men_n82_), .B(men_men_n87_), .Y(men_men_n88_));
  NAi21      u0066(.An(i_6_), .B(i_10_), .Y(men_men_n89_));
  NA2        u0067(.A(i_6_), .B(i_9_), .Y(men_men_n90_));
  AOI210     u0068(.A0(men_men_n90_), .A1(men_men_n89_), .B0(men_men_n61_), .Y(men_men_n91_));
  NA2        u0069(.A(i_2_), .B(i_6_), .Y(men_men_n92_));
  NO3        u0070(.A(men_men_n92_), .B(men_men_n50_), .C(men_men_n25_), .Y(men_men_n93_));
  NO2        u0071(.A(men_men_n93_), .B(men_men_n91_), .Y(men_men_n94_));
  AOI210     u0072(.A0(men_men_n94_), .A1(men_men_n88_), .B0(men_men_n78_), .Y(men_men_n95_));
  AN3        u0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n96_));
  NAi21      u0074(.An(i_6_), .B(i_11_), .Y(men_men_n97_));
  NO2        u0075(.A(i_5_), .B(i_8_), .Y(men_men_n98_));
  NOi21      u0076(.An(men_men_n98_), .B(men_men_n97_), .Y(men_men_n99_));
  AOI220     u0077(.A0(men_men_n99_), .A1(men_men_n60_), .B0(men_men_n96_), .B1(men_men_n32_), .Y(men_men_n100_));
  INV        u0078(.A(i_7_), .Y(men_men_n101_));
  NA2        u0079(.A(men_men_n47_), .B(men_men_n101_), .Y(men_men_n102_));
  NO2        u0080(.A(i_0_), .B(i_5_), .Y(men_men_n103_));
  NO2        u0081(.A(men_men_n103_), .B(men_men_n83_), .Y(men_men_n104_));
  NA2        u0082(.A(i_12_), .B(i_3_), .Y(men_men_n105_));
  INV        u0083(.A(men_men_n105_), .Y(men_men_n106_));
  NA3        u0084(.A(men_men_n106_), .B(men_men_n104_), .C(men_men_n102_), .Y(men_men_n107_));
  NAi21      u0085(.An(i_7_), .B(i_11_), .Y(men_men_n108_));
  NO3        u0086(.A(men_men_n108_), .B(men_men_n89_), .C(men_men_n52_), .Y(men_men_n109_));
  AN2        u0087(.A(i_2_), .B(i_10_), .Y(men_men_n110_));
  NO2        u0088(.A(men_men_n110_), .B(i_7_), .Y(men_men_n111_));
  OR2        u0089(.A(men_men_n78_), .B(men_men_n56_), .Y(men_men_n112_));
  NO2        u0090(.A(i_8_), .B(men_men_n101_), .Y(men_men_n113_));
  NO3        u0091(.A(men_men_n113_), .B(men_men_n112_), .C(men_men_n111_), .Y(men_men_n114_));
  NA2        u0092(.A(i_12_), .B(i_7_), .Y(men_men_n115_));
  NO2        u0093(.A(men_men_n61_), .B(men_men_n26_), .Y(men_men_n116_));
  NA2        u0094(.A(men_men_n116_), .B(i_0_), .Y(men_men_n117_));
  NA2        u0095(.A(i_11_), .B(i_12_), .Y(men_men_n118_));
  OAI210     u0096(.A0(men_men_n117_), .A1(men_men_n115_), .B0(men_men_n118_), .Y(men_men_n119_));
  NO2        u0097(.A(men_men_n119_), .B(men_men_n114_), .Y(men_men_n120_));
  NAi41      u0098(.An(men_men_n109_), .B(men_men_n120_), .C(men_men_n107_), .D(men_men_n100_), .Y(men_men_n121_));
  NOi21      u0099(.An(i_1_), .B(i_5_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n122_), .B(i_11_), .Y(men_men_n123_));
  NA2        u0101(.A(men_men_n101_), .B(men_men_n37_), .Y(men_men_n124_));
  NA2        u0102(.A(i_7_), .B(men_men_n25_), .Y(men_men_n125_));
  NA2        u0103(.A(men_men_n125_), .B(men_men_n124_), .Y(men_men_n126_));
  NO2        u0104(.A(men_men_n126_), .B(men_men_n47_), .Y(men_men_n127_));
  NA2        u0105(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n128_));
  NAi21      u0106(.An(i_3_), .B(i_8_), .Y(men_men_n129_));
  NA2        u0107(.A(men_men_n129_), .B(men_men_n60_), .Y(men_men_n130_));
  NOi21      u0108(.An(men_men_n130_), .B(men_men_n128_), .Y(men_men_n131_));
  NO2        u0109(.A(i_1_), .B(men_men_n83_), .Y(men_men_n132_));
  NO2        u0110(.A(i_6_), .B(i_5_), .Y(men_men_n133_));
  NA2        u0111(.A(men_men_n133_), .B(i_3_), .Y(men_men_n134_));
  AO210      u0112(.A0(men_men_n134_), .A1(men_men_n48_), .B0(men_men_n132_), .Y(men_men_n135_));
  OAI220     u0113(.A0(men_men_n135_), .A1(men_men_n108_), .B0(men_men_n131_), .B1(men_men_n123_), .Y(men_men_n136_));
  NO3        u0114(.A(men_men_n136_), .B(men_men_n121_), .C(men_men_n95_), .Y(men_men_n137_));
  NA2        u0115(.A(men_men_n137_), .B(men_men_n77_), .Y(men2));
  NO2        u0116(.A(men_men_n61_), .B(men_men_n37_), .Y(men_men_n139_));
  NA2        u0117(.A(i_6_), .B(men_men_n25_), .Y(men_men_n140_));
  NA2        u0118(.A(men_men_n140_), .B(men_men_n139_), .Y(men_men_n141_));
  NA4        u0119(.A(men_men_n141_), .B(men_men_n75_), .C(men_men_n67_), .D(men_men_n30_), .Y(men0));
  AN2        u0120(.A(i_8_), .B(i_7_), .Y(men_men_n143_));
  NA2        u0121(.A(men_men_n143_), .B(i_6_), .Y(men_men_n144_));
  NO2        u0122(.A(i_12_), .B(i_13_), .Y(men_men_n145_));
  NAi21      u0123(.An(i_5_), .B(i_11_), .Y(men_men_n146_));
  NOi21      u0124(.An(men_men_n145_), .B(men_men_n146_), .Y(men_men_n147_));
  NO2        u0125(.A(i_0_), .B(i_1_), .Y(men_men_n148_));
  NA2        u0126(.A(i_2_), .B(i_3_), .Y(men_men_n149_));
  NO2        u0127(.A(men_men_n149_), .B(i_4_), .Y(men_men_n150_));
  NA3        u0128(.A(men_men_n150_), .B(men_men_n148_), .C(men_men_n147_), .Y(men_men_n151_));
  OR2        u0129(.A(men_men_n151_), .B(men_men_n25_), .Y(men_men_n152_));
  AN2        u0130(.A(men_men_n145_), .B(men_men_n80_), .Y(men_men_n153_));
  NO2        u0131(.A(men_men_n153_), .B(men_men_n27_), .Y(men_men_n154_));
  NA2        u0132(.A(i_1_), .B(i_5_), .Y(men_men_n155_));
  NO2        u0133(.A(men_men_n71_), .B(men_men_n47_), .Y(men_men_n156_));
  NA2        u0134(.A(men_men_n156_), .B(men_men_n36_), .Y(men_men_n157_));
  NO3        u0135(.A(men_men_n157_), .B(men_men_n155_), .C(men_men_n154_), .Y(men_men_n158_));
  OR2        u0136(.A(i_0_), .B(i_1_), .Y(men_men_n159_));
  NO3        u0137(.A(men_men_n159_), .B(men_men_n78_), .C(i_13_), .Y(men_men_n160_));
  NAi32      u0138(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n161_));
  NAi21      u0139(.An(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  NOi21      u0140(.An(i_4_), .B(i_10_), .Y(men_men_n163_));
  NA2        u0141(.A(men_men_n163_), .B(men_men_n40_), .Y(men_men_n164_));
  NO2        u0142(.A(i_3_), .B(i_5_), .Y(men_men_n165_));
  NO3        u0143(.A(men_men_n71_), .B(i_2_), .C(i_1_), .Y(men_men_n166_));
  NA2        u0144(.A(men_men_n166_), .B(men_men_n165_), .Y(men_men_n167_));
  OAI210     u0145(.A0(men_men_n167_), .A1(men_men_n164_), .B0(men_men_n162_), .Y(men_men_n168_));
  NO2        u0146(.A(men_men_n168_), .B(men_men_n158_), .Y(men_men_n169_));
  AOI210     u0147(.A0(men_men_n169_), .A1(men_men_n152_), .B0(men_men_n144_), .Y(men_men_n170_));
  NA2        u0148(.A(i_3_), .B(men_men_n49_), .Y(men_men_n171_));
  NOi21      u0149(.An(i_4_), .B(i_9_), .Y(men_men_n172_));
  NOi21      u0150(.An(i_11_), .B(i_13_), .Y(men_men_n173_));
  NA2        u0151(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  NO2        u0152(.A(i_4_), .B(i_5_), .Y(men_men_n175_));
  NAi21      u0153(.An(i_12_), .B(i_11_), .Y(men_men_n176_));
  NO2        u0154(.A(men_men_n176_), .B(i_13_), .Y(men_men_n177_));
  NA3        u0155(.A(men_men_n177_), .B(men_men_n175_), .C(men_men_n80_), .Y(men_men_n178_));
  AOI210     u0156(.A0(men_men_n178_), .A1(men_men_n174_), .B0(i_2_), .Y(men_men_n179_));
  NO2        u0157(.A(men_men_n71_), .B(men_men_n61_), .Y(men_men_n180_));
  NAi31      u0158(.An(men_men_n1101_), .B(men_men_n153_), .C(i_11_), .Y(men_men_n181_));
  NA2        u0159(.A(i_3_), .B(i_5_), .Y(men_men_n182_));
  AOI210     u0160(.A0(men_men_n174_), .A1(men_men_n181_), .B0(i_2_), .Y(men_men_n183_));
  NO2        u0161(.A(men_men_n71_), .B(i_5_), .Y(men_men_n184_));
  NO2        u0162(.A(i_13_), .B(i_10_), .Y(men_men_n185_));
  NA3        u0163(.A(men_men_n185_), .B(men_men_n184_), .C(men_men_n45_), .Y(men_men_n186_));
  NO2        u0164(.A(i_2_), .B(i_1_), .Y(men_men_n187_));
  NA2        u0165(.A(men_men_n187_), .B(i_3_), .Y(men_men_n188_));
  NAi21      u0166(.An(i_4_), .B(i_12_), .Y(men_men_n189_));
  NO4        u0167(.A(men_men_n189_), .B(men_men_n188_), .C(men_men_n186_), .D(men_men_n25_), .Y(men_men_n190_));
  NO3        u0168(.A(men_men_n190_), .B(men_men_n183_), .C(men_men_n179_), .Y(men_men_n191_));
  INV        u0169(.A(i_8_), .Y(men_men_n192_));
  NO2        u0170(.A(men_men_n192_), .B(i_7_), .Y(men_men_n193_));
  NA2        u0171(.A(men_men_n193_), .B(i_6_), .Y(men_men_n194_));
  NO3        u0172(.A(i_3_), .B(men_men_n83_), .C(men_men_n49_), .Y(men_men_n195_));
  NA2        u0173(.A(men_men_n195_), .B(men_men_n113_), .Y(men_men_n196_));
  NO3        u0174(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n197_));
  NA3        u0175(.A(men_men_n197_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n198_));
  NO3        u0176(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n199_));
  OAI210     u0177(.A0(men_men_n96_), .A1(i_12_), .B0(men_men_n199_), .Y(men_men_n200_));
  AOI210     u0178(.A0(men_men_n200_), .A1(men_men_n198_), .B0(men_men_n196_), .Y(men_men_n201_));
  NO2        u0179(.A(i_3_), .B(i_8_), .Y(men_men_n202_));
  NO3        u0180(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n203_));
  NA3        u0181(.A(men_men_n203_), .B(men_men_n202_), .C(men_men_n40_), .Y(men_men_n204_));
  NO2        u0182(.A(men_men_n103_), .B(men_men_n56_), .Y(men_men_n205_));
  NO2        u0183(.A(i_13_), .B(i_9_), .Y(men_men_n206_));
  NA3        u0184(.A(men_men_n206_), .B(i_6_), .C(men_men_n192_), .Y(men_men_n207_));
  NAi21      u0185(.An(i_12_), .B(i_3_), .Y(men_men_n208_));
  OR2        u0186(.A(men_men_n208_), .B(men_men_n207_), .Y(men_men_n209_));
  NO2        u0187(.A(men_men_n45_), .B(i_5_), .Y(men_men_n210_));
  NO3        u0188(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n211_));
  NA2        u0189(.A(men_men_n211_), .B(i_10_), .Y(men_men_n212_));
  OAI220     u0190(.A0(men_men_n212_), .A1(men_men_n209_), .B0(men_men_n103_), .B1(men_men_n204_), .Y(men_men_n213_));
  AOI210     u0191(.A0(men_men_n213_), .A1(i_7_), .B0(men_men_n201_), .Y(men_men_n214_));
  OAI220     u0192(.A0(men_men_n214_), .A1(i_4_), .B0(men_men_n194_), .B1(men_men_n191_), .Y(men_men_n215_));
  NAi21      u0193(.An(i_12_), .B(i_7_), .Y(men_men_n216_));
  NA3        u0194(.A(i_13_), .B(men_men_n192_), .C(i_10_), .Y(men_men_n217_));
  NO2        u0195(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n218_));
  NA2        u0196(.A(i_0_), .B(i_5_), .Y(men_men_n219_));
  NA2        u0197(.A(men_men_n219_), .B(men_men_n104_), .Y(men_men_n220_));
  OAI220     u0198(.A0(men_men_n220_), .A1(men_men_n188_), .B0(i_2_), .B1(men_men_n134_), .Y(men_men_n221_));
  NAi31      u0199(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n222_));
  NO2        u0200(.A(men_men_n36_), .B(i_13_), .Y(men_men_n223_));
  NO2        u0201(.A(men_men_n71_), .B(men_men_n26_), .Y(men_men_n224_));
  NO2        u0202(.A(men_men_n47_), .B(men_men_n61_), .Y(men_men_n225_));
  NA3        u0203(.A(men_men_n225_), .B(men_men_n224_), .C(men_men_n223_), .Y(men_men_n226_));
  INV        u0204(.A(i_13_), .Y(men_men_n227_));
  NO2        u0205(.A(i_12_), .B(men_men_n227_), .Y(men_men_n228_));
  NA3        u0206(.A(men_men_n228_), .B(men_men_n197_), .C(men_men_n195_), .Y(men_men_n229_));
  OAI210     u0207(.A0(men_men_n226_), .A1(men_men_n222_), .B0(men_men_n229_), .Y(men_men_n230_));
  AOI220     u0208(.A0(men_men_n230_), .A1(men_men_n143_), .B0(men_men_n221_), .B1(men_men_n218_), .Y(men_men_n231_));
  NO2        u0209(.A(i_12_), .B(men_men_n37_), .Y(men_men_n232_));
  NO2        u0210(.A(men_men_n182_), .B(i_4_), .Y(men_men_n233_));
  NA2        u0211(.A(men_men_n233_), .B(men_men_n232_), .Y(men_men_n234_));
  OR2        u0212(.A(i_8_), .B(i_7_), .Y(men_men_n235_));
  NO2        u0213(.A(men_men_n235_), .B(men_men_n83_), .Y(men_men_n236_));
  NO2        u0214(.A(men_men_n52_), .B(i_1_), .Y(men_men_n237_));
  NA2        u0215(.A(men_men_n237_), .B(men_men_n236_), .Y(men_men_n238_));
  INV        u0216(.A(i_12_), .Y(men_men_n239_));
  NO3        u0217(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n240_));
  NA2        u0218(.A(i_2_), .B(i_1_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n238_), .B(men_men_n234_), .Y(men_men_n242_));
  NO3        u0220(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n243_));
  NAi21      u0221(.An(i_4_), .B(i_3_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n244_), .B(men_men_n73_), .Y(men_men_n245_));
  NO2        u0223(.A(i_0_), .B(i_6_), .Y(men_men_n246_));
  NOi41      u0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n247_));
  NA2        u0225(.A(men_men_n247_), .B(men_men_n246_), .Y(men_men_n248_));
  NO2        u0226(.A(men_men_n241_), .B(men_men_n182_), .Y(men_men_n249_));
  NA2        u0227(.A(men_men_n242_), .B(men_men_n206_), .Y(men_men_n250_));
  NO2        u0228(.A(i_11_), .B(men_men_n227_), .Y(men_men_n251_));
  NOi21      u0229(.An(i_1_), .B(i_6_), .Y(men_men_n252_));
  NAi21      u0230(.An(i_3_), .B(i_7_), .Y(men_men_n253_));
  NA2        u0231(.A(men_men_n239_), .B(i_9_), .Y(men_men_n254_));
  OR4        u0232(.A(men_men_n254_), .B(men_men_n253_), .C(men_men_n252_), .D(men_men_n184_), .Y(men_men_n255_));
  NO2        u0233(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n256_));
  NO2        u0234(.A(i_12_), .B(i_3_), .Y(men_men_n257_));
  NA2        u0235(.A(men_men_n71_), .B(i_5_), .Y(men_men_n258_));
  NA2        u0236(.A(i_3_), .B(i_9_), .Y(men_men_n259_));
  NAi21      u0237(.An(i_7_), .B(i_10_), .Y(men_men_n260_));
  NO2        u0238(.A(men_men_n260_), .B(men_men_n259_), .Y(men_men_n261_));
  NA3        u0239(.A(men_men_n261_), .B(men_men_n258_), .C(men_men_n62_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n262_), .B(men_men_n255_), .Y(men_men_n263_));
  NA3        u0241(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n264_));
  NA2        u0242(.A(men_men_n263_), .B(men_men_n251_), .Y(men_men_n265_));
  NO2        u0243(.A(men_men_n235_), .B(men_men_n37_), .Y(men_men_n266_));
  NA2        u0244(.A(i_12_), .B(i_6_), .Y(men_men_n267_));
  OR2        u0245(.A(i_13_), .B(i_9_), .Y(men_men_n268_));
  NO3        u0246(.A(men_men_n268_), .B(men_men_n267_), .C(men_men_n49_), .Y(men_men_n269_));
  NO2        u0247(.A(men_men_n244_), .B(i_2_), .Y(men_men_n270_));
  NA3        u0248(.A(men_men_n270_), .B(men_men_n269_), .C(men_men_n45_), .Y(men_men_n271_));
  NA2        u0249(.A(men_men_n251_), .B(i_9_), .Y(men_men_n272_));
  NA2        u0250(.A(men_men_n258_), .B(men_men_n62_), .Y(men_men_n273_));
  OAI210     u0251(.A0(men_men_n273_), .A1(men_men_n272_), .B0(men_men_n271_), .Y(men_men_n274_));
  NA2        u0252(.A(men_men_n156_), .B(men_men_n61_), .Y(men_men_n275_));
  NO3        u0253(.A(i_11_), .B(men_men_n227_), .C(men_men_n25_), .Y(men_men_n276_));
  NO2        u0254(.A(men_men_n253_), .B(i_8_), .Y(men_men_n277_));
  NO2        u0255(.A(i_6_), .B(men_men_n49_), .Y(men_men_n278_));
  NA3        u0256(.A(men_men_n278_), .B(men_men_n277_), .C(men_men_n276_), .Y(men_men_n279_));
  NO3        u0257(.A(men_men_n26_), .B(men_men_n83_), .C(i_5_), .Y(men_men_n280_));
  NA3        u0258(.A(men_men_n280_), .B(men_men_n266_), .C(men_men_n228_), .Y(men_men_n281_));
  AOI210     u0259(.A0(men_men_n281_), .A1(men_men_n279_), .B0(men_men_n275_), .Y(men_men_n282_));
  AOI210     u0260(.A0(men_men_n274_), .A1(men_men_n266_), .B0(men_men_n282_), .Y(men_men_n283_));
  NA4        u0261(.A(men_men_n283_), .B(men_men_n265_), .C(men_men_n250_), .D(men_men_n231_), .Y(men_men_n284_));
  NO3        u0262(.A(i_12_), .B(men_men_n227_), .C(men_men_n37_), .Y(men_men_n285_));
  INV        u0263(.A(men_men_n285_), .Y(men_men_n286_));
  NA2        u0264(.A(i_8_), .B(men_men_n101_), .Y(men_men_n287_));
  NOi21      u0265(.An(men_men_n165_), .B(men_men_n83_), .Y(men_men_n288_));
  NO3        u0266(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n289_));
  AOI220     u0267(.A0(men_men_n289_), .A1(men_men_n195_), .B0(men_men_n288_), .B1(men_men_n237_), .Y(men_men_n290_));
  NO2        u0268(.A(men_men_n290_), .B(men_men_n287_), .Y(men_men_n291_));
  NO3        u0269(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n292_));
  NO2        u0270(.A(men_men_n241_), .B(i_0_), .Y(men_men_n293_));
  AOI220     u0271(.A0(men_men_n293_), .A1(men_men_n193_), .B0(men_men_n292_), .B1(men_men_n143_), .Y(men_men_n294_));
  NA2        u0272(.A(men_men_n278_), .B(men_men_n26_), .Y(men_men_n295_));
  NO2        u0273(.A(men_men_n295_), .B(men_men_n294_), .Y(men_men_n296_));
  NA2        u0274(.A(i_0_), .B(i_1_), .Y(men_men_n297_));
  NO2        u0275(.A(men_men_n297_), .B(i_2_), .Y(men_men_n298_));
  NO2        u0276(.A(men_men_n57_), .B(i_6_), .Y(men_men_n299_));
  NA3        u0277(.A(men_men_n299_), .B(men_men_n298_), .C(men_men_n165_), .Y(men_men_n300_));
  OAI210     u0278(.A0(men_men_n167_), .A1(men_men_n144_), .B0(men_men_n300_), .Y(men_men_n301_));
  NO3        u0279(.A(men_men_n301_), .B(men_men_n296_), .C(men_men_n291_), .Y(men_men_n302_));
  NO2        u0280(.A(i_3_), .B(i_10_), .Y(men_men_n303_));
  NA3        u0281(.A(men_men_n303_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n304_));
  NO2        u0282(.A(i_2_), .B(men_men_n101_), .Y(men_men_n305_));
  NOi21      u0283(.An(men_men_n219_), .B(men_men_n103_), .Y(men_men_n306_));
  NA3        u0284(.A(men_men_n306_), .B(i_1_), .C(men_men_n305_), .Y(men_men_n307_));
  AN2        u0285(.A(i_3_), .B(i_10_), .Y(men_men_n308_));
  NA4        u0286(.A(men_men_n308_), .B(men_men_n197_), .C(men_men_n177_), .D(men_men_n175_), .Y(men_men_n309_));
  NO2        u0287(.A(i_5_), .B(men_men_n37_), .Y(men_men_n310_));
  NO2        u0288(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n311_));
  OR2        u0289(.A(men_men_n307_), .B(men_men_n304_), .Y(men_men_n312_));
  OAI220     u0290(.A0(men_men_n312_), .A1(i_6_), .B0(men_men_n302_), .B1(men_men_n286_), .Y(men_men_n313_));
  NO4        u0291(.A(men_men_n313_), .B(men_men_n284_), .C(men_men_n215_), .D(men_men_n170_), .Y(men_men_n314_));
  NO3        u0292(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n315_));
  NO2        u0293(.A(men_men_n57_), .B(men_men_n83_), .Y(men_men_n316_));
  NA2        u0294(.A(men_men_n293_), .B(men_men_n316_), .Y(men_men_n317_));
  NO3        u0295(.A(i_6_), .B(men_men_n192_), .C(i_7_), .Y(men_men_n318_));
  NA2        u0296(.A(men_men_n318_), .B(men_men_n197_), .Y(men_men_n319_));
  AOI210     u0297(.A0(men_men_n319_), .A1(men_men_n317_), .B0(men_men_n171_), .Y(men_men_n320_));
  NO2        u0298(.A(i_2_), .B(i_3_), .Y(men_men_n321_));
  OR2        u0299(.A(i_0_), .B(i_5_), .Y(men_men_n322_));
  NA2        u0300(.A(men_men_n219_), .B(men_men_n322_), .Y(men_men_n323_));
  NA4        u0301(.A(men_men_n323_), .B(men_men_n236_), .C(men_men_n321_), .D(i_1_), .Y(men_men_n324_));
  NA3        u0302(.A(men_men_n293_), .B(men_men_n288_), .C(men_men_n113_), .Y(men_men_n325_));
  NO2        u0303(.A(men_men_n159_), .B(men_men_n47_), .Y(men_men_n326_));
  NA3        u0304(.A(men_men_n326_), .B(i_7_), .C(men_men_n165_), .Y(men_men_n327_));
  NA3        u0305(.A(men_men_n327_), .B(men_men_n325_), .C(men_men_n324_), .Y(men_men_n328_));
  OAI210     u0306(.A0(men_men_n328_), .A1(men_men_n320_), .B0(i_4_), .Y(men_men_n329_));
  NO2        u0307(.A(i_12_), .B(i_10_), .Y(men_men_n330_));
  NOi21      u0308(.An(i_5_), .B(i_0_), .Y(men_men_n331_));
  AOI210     u0309(.A0(i_2_), .A1(men_men_n49_), .B0(men_men_n101_), .Y(men_men_n332_));
  NO3        u0310(.A(men_men_n332_), .B(i_4_), .C(men_men_n129_), .Y(men_men_n333_));
  NA4        u0311(.A(men_men_n81_), .B(men_men_n36_), .C(men_men_n83_), .D(i_8_), .Y(men_men_n334_));
  NA2        u0312(.A(men_men_n333_), .B(men_men_n330_), .Y(men_men_n335_));
  NO2        u0313(.A(i_6_), .B(i_8_), .Y(men_men_n336_));
  NOi21      u0314(.An(i_0_), .B(i_2_), .Y(men_men_n337_));
  AN2        u0315(.A(men_men_n337_), .B(men_men_n336_), .Y(men_men_n338_));
  NO2        u0316(.A(i_1_), .B(i_7_), .Y(men_men_n339_));
  NA3        u0317(.A(men_men_n336_), .B(men_men_n42_), .C(i_5_), .Y(men_men_n340_));
  NA3        u0318(.A(men_men_n340_), .B(men_men_n335_), .C(men_men_n329_), .Y(men_men_n341_));
  NO2        u0319(.A(i_8_), .B(men_men_n323_), .Y(men_men_n342_));
  NOi21      u0320(.An(men_men_n155_), .B(men_men_n104_), .Y(men_men_n343_));
  NO2        u0321(.A(men_men_n343_), .B(men_men_n125_), .Y(men_men_n344_));
  OAI210     u0322(.A0(men_men_n344_), .A1(men_men_n342_), .B0(i_3_), .Y(men_men_n345_));
  INV        u0323(.A(men_men_n81_), .Y(men_men_n346_));
  NO2        u0324(.A(men_men_n297_), .B(men_men_n79_), .Y(men_men_n347_));
  NA2        u0325(.A(men_men_n347_), .B(men_men_n133_), .Y(men_men_n348_));
  NO2        u0326(.A(men_men_n92_), .B(men_men_n192_), .Y(men_men_n349_));
  NA3        u0327(.A(men_men_n306_), .B(men_men_n349_), .C(men_men_n61_), .Y(men_men_n350_));
  AOI210     u0328(.A0(men_men_n350_), .A1(men_men_n348_), .B0(men_men_n346_), .Y(men_men_n351_));
  NO2        u0329(.A(men_men_n192_), .B(i_9_), .Y(men_men_n352_));
  NA2        u0330(.A(men_men_n352_), .B(men_men_n205_), .Y(men_men_n353_));
  NO2        u0331(.A(men_men_n351_), .B(men_men_n296_), .Y(men_men_n354_));
  AOI210     u0332(.A0(men_men_n354_), .A1(men_men_n345_), .B0(men_men_n164_), .Y(men_men_n355_));
  AOI210     u0333(.A0(men_men_n341_), .A1(men_men_n315_), .B0(men_men_n355_), .Y(men_men_n356_));
  NOi32      u0334(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n357_));
  INV        u0335(.A(men_men_n357_), .Y(men_men_n358_));
  NAi21      u0336(.An(i_0_), .B(i_6_), .Y(men_men_n359_));
  NAi21      u0337(.An(i_1_), .B(i_5_), .Y(men_men_n360_));
  NA2        u0338(.A(men_men_n360_), .B(men_men_n359_), .Y(men_men_n361_));
  NA2        u0339(.A(men_men_n361_), .B(men_men_n25_), .Y(men_men_n362_));
  OAI210     u0340(.A0(men_men_n362_), .A1(men_men_n161_), .B0(men_men_n248_), .Y(men_men_n363_));
  NAi41      u0341(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n364_));
  OAI220     u0342(.A0(men_men_n364_), .A1(men_men_n360_), .B0(men_men_n222_), .B1(men_men_n161_), .Y(men_men_n365_));
  AOI210     u0343(.A0(men_men_n364_), .A1(men_men_n161_), .B0(men_men_n159_), .Y(men_men_n366_));
  NOi32      u0344(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n367_));
  NAi21      u0345(.An(i_6_), .B(i_1_), .Y(men_men_n368_));
  NA3        u0346(.A(men_men_n368_), .B(men_men_n367_), .C(men_men_n47_), .Y(men_men_n369_));
  NO2        u0347(.A(men_men_n369_), .B(i_0_), .Y(men_men_n370_));
  OR3        u0348(.A(men_men_n370_), .B(men_men_n366_), .C(men_men_n365_), .Y(men_men_n371_));
  NO2        u0349(.A(i_1_), .B(men_men_n101_), .Y(men_men_n372_));
  NAi21      u0350(.An(i_3_), .B(i_4_), .Y(men_men_n373_));
  NO2        u0351(.A(men_men_n373_), .B(i_9_), .Y(men_men_n374_));
  AN2        u0352(.A(i_6_), .B(i_7_), .Y(men_men_n375_));
  OAI210     u0353(.A0(men_men_n375_), .A1(men_men_n372_), .B0(men_men_n374_), .Y(men_men_n376_));
  NA2        u0354(.A(i_2_), .B(i_7_), .Y(men_men_n377_));
  NO2        u0355(.A(men_men_n373_), .B(i_10_), .Y(men_men_n378_));
  NA3        u0356(.A(men_men_n378_), .B(men_men_n377_), .C(men_men_n246_), .Y(men_men_n379_));
  AOI210     u0357(.A0(men_men_n379_), .A1(men_men_n376_), .B0(men_men_n184_), .Y(men_men_n380_));
  AOI210     u0358(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n381_));
  NA2        u0359(.A(men_men_n378_), .B(men_men_n339_), .Y(men_men_n382_));
  NO3        u0360(.A(men_men_n380_), .B(men_men_n371_), .C(men_men_n363_), .Y(men_men_n383_));
  NO2        u0361(.A(men_men_n383_), .B(men_men_n358_), .Y(men_men_n384_));
  NO2        u0362(.A(men_men_n57_), .B(men_men_n25_), .Y(men_men_n385_));
  AN2        u0363(.A(i_12_), .B(i_5_), .Y(men_men_n386_));
  NO2        u0364(.A(i_4_), .B(men_men_n26_), .Y(men_men_n387_));
  NA2        u0365(.A(men_men_n387_), .B(men_men_n386_), .Y(men_men_n388_));
  NO2        u0366(.A(i_11_), .B(i_6_), .Y(men_men_n389_));
  NA3        u0367(.A(men_men_n389_), .B(men_men_n326_), .C(men_men_n227_), .Y(men_men_n390_));
  NO2        u0368(.A(men_men_n390_), .B(men_men_n388_), .Y(men_men_n391_));
  NO2        u0369(.A(men_men_n244_), .B(i_5_), .Y(men_men_n392_));
  NO2        u0370(.A(i_5_), .B(i_10_), .Y(men_men_n393_));
  NA2        u0371(.A(men_men_n145_), .B(men_men_n46_), .Y(men_men_n394_));
  NO2        u0372(.A(men_men_n394_), .B(men_men_n1100_), .Y(men_men_n395_));
  OAI210     u0373(.A0(men_men_n395_), .A1(men_men_n391_), .B0(men_men_n385_), .Y(men_men_n396_));
  NO2        u0374(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n397_));
  NO2        u0375(.A(men_men_n151_), .B(men_men_n83_), .Y(men_men_n398_));
  OAI210     u0376(.A0(men_men_n398_), .A1(men_men_n391_), .B0(men_men_n397_), .Y(men_men_n399_));
  NO3        u0377(.A(men_men_n83_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n400_));
  NO2        u0378(.A(i_3_), .B(men_men_n101_), .Y(men_men_n401_));
  NA3        u0379(.A(men_men_n303_), .B(men_men_n73_), .C(men_men_n53_), .Y(men_men_n402_));
  NO2        u0380(.A(i_11_), .B(i_12_), .Y(men_men_n403_));
  NA2        u0381(.A(men_men_n403_), .B(men_men_n36_), .Y(men_men_n404_));
  NO2        u0382(.A(men_men_n402_), .B(men_men_n404_), .Y(men_men_n405_));
  NA2        u0383(.A(men_men_n393_), .B(men_men_n239_), .Y(men_men_n406_));
  NA3        u0384(.A(men_men_n113_), .B(men_men_n42_), .C(i_11_), .Y(men_men_n407_));
  NO2        u0385(.A(men_men_n407_), .B(men_men_n222_), .Y(men_men_n408_));
  NAi21      u0386(.An(i_13_), .B(i_0_), .Y(men_men_n409_));
  NO2        u0387(.A(men_men_n409_), .B(men_men_n241_), .Y(men_men_n410_));
  OAI210     u0388(.A0(men_men_n408_), .A1(men_men_n405_), .B0(men_men_n410_), .Y(men_men_n411_));
  NA3        u0389(.A(men_men_n411_), .B(men_men_n399_), .C(men_men_n396_), .Y(men_men_n412_));
  NO3        u0390(.A(i_1_), .B(i_12_), .C(men_men_n83_), .Y(men_men_n413_));
  NO2        u0391(.A(i_0_), .B(i_11_), .Y(men_men_n414_));
  AN2        u0392(.A(i_1_), .B(i_6_), .Y(men_men_n415_));
  NOi21      u0393(.An(i_2_), .B(i_12_), .Y(men_men_n416_));
  NA2        u0394(.A(men_men_n416_), .B(men_men_n415_), .Y(men_men_n417_));
  NO2        u0395(.A(men_men_n417_), .B(men_men_n1096_), .Y(men_men_n418_));
  NA2        u0396(.A(men_men_n143_), .B(i_9_), .Y(men_men_n419_));
  NO2        u0397(.A(men_men_n419_), .B(i_4_), .Y(men_men_n420_));
  NA2        u0398(.A(men_men_n418_), .B(men_men_n420_), .Y(men_men_n421_));
  NAi21      u0399(.An(i_9_), .B(i_4_), .Y(men_men_n422_));
  OR2        u0400(.A(i_13_), .B(i_10_), .Y(men_men_n423_));
  NO3        u0401(.A(men_men_n423_), .B(men_men_n118_), .C(men_men_n422_), .Y(men_men_n424_));
  NO2        u0402(.A(men_men_n174_), .B(men_men_n124_), .Y(men_men_n425_));
  BUFFER     u0403(.A(men_men_n217_), .Y(men_men_n426_));
  NO2        u0404(.A(men_men_n101_), .B(men_men_n25_), .Y(men_men_n427_));
  NA2        u0405(.A(men_men_n285_), .B(men_men_n427_), .Y(men_men_n428_));
  NA2        u0406(.A(men_men_n278_), .B(men_men_n211_), .Y(men_men_n429_));
  OAI220     u0407(.A0(men_men_n429_), .A1(men_men_n426_), .B0(men_men_n428_), .B1(men_men_n343_), .Y(men_men_n430_));
  INV        u0408(.A(men_men_n430_), .Y(men_men_n431_));
  AOI210     u0409(.A0(men_men_n431_), .A1(men_men_n421_), .B0(men_men_n26_), .Y(men_men_n432_));
  NA2        u0410(.A(men_men_n325_), .B(men_men_n324_), .Y(men_men_n433_));
  AOI220     u0411(.A0(men_men_n299_), .A1(men_men_n289_), .B0(men_men_n293_), .B1(men_men_n316_), .Y(men_men_n434_));
  NO2        u0412(.A(men_men_n434_), .B(men_men_n171_), .Y(men_men_n435_));
  NO2        u0413(.A(men_men_n182_), .B(men_men_n83_), .Y(men_men_n436_));
  AOI220     u0414(.A0(men_men_n436_), .A1(men_men_n298_), .B0(men_men_n280_), .B1(men_men_n211_), .Y(men_men_n437_));
  NO2        u0415(.A(men_men_n437_), .B(men_men_n287_), .Y(men_men_n438_));
  NO3        u0416(.A(men_men_n438_), .B(men_men_n435_), .C(men_men_n433_), .Y(men_men_n439_));
  NA2        u0417(.A(men_men_n195_), .B(men_men_n96_), .Y(men_men_n440_));
  NA3        u0418(.A(men_men_n326_), .B(men_men_n165_), .C(men_men_n83_), .Y(men_men_n441_));
  AOI210     u0419(.A0(men_men_n441_), .A1(men_men_n440_), .B0(i_8_), .Y(men_men_n442_));
  NA2        u0420(.A(men_men_n192_), .B(i_10_), .Y(men_men_n443_));
  NA3        u0421(.A(men_men_n258_), .B(men_men_n62_), .C(i_2_), .Y(men_men_n444_));
  NA2        u0422(.A(men_men_n299_), .B(men_men_n237_), .Y(men_men_n445_));
  OAI220     u0423(.A0(men_men_n445_), .A1(men_men_n182_), .B0(men_men_n444_), .B1(men_men_n443_), .Y(men_men_n446_));
  NO2        u0424(.A(i_3_), .B(men_men_n49_), .Y(men_men_n447_));
  NA3        u0425(.A(men_men_n339_), .B(men_men_n338_), .C(men_men_n447_), .Y(men_men_n448_));
  NA2        u0426(.A(men_men_n318_), .B(men_men_n323_), .Y(men_men_n449_));
  OAI210     u0427(.A0(men_men_n449_), .A1(men_men_n188_), .B0(men_men_n448_), .Y(men_men_n450_));
  NO3        u0428(.A(men_men_n450_), .B(men_men_n446_), .C(men_men_n442_), .Y(men_men_n451_));
  AOI210     u0429(.A0(men_men_n451_), .A1(men_men_n439_), .B0(men_men_n272_), .Y(men_men_n452_));
  NO4        u0430(.A(men_men_n452_), .B(men_men_n432_), .C(men_men_n412_), .D(men_men_n384_), .Y(men_men_n453_));
  NO2        u0431(.A(men_men_n61_), .B(i_4_), .Y(men_men_n454_));
  NO2        u0432(.A(men_men_n71_), .B(i_13_), .Y(men_men_n455_));
  NO2        u0433(.A(i_10_), .B(i_9_), .Y(men_men_n456_));
  NAi21      u0434(.An(i_12_), .B(i_8_), .Y(men_men_n457_));
  NO2        u0435(.A(men_men_n457_), .B(i_3_), .Y(men_men_n458_));
  NA2        u0436(.A(i_2_), .B(men_men_n104_), .Y(men_men_n459_));
  NO2        u0437(.A(men_men_n459_), .B(men_men_n204_), .Y(men_men_n460_));
  NA2        u0438(.A(men_men_n311_), .B(i_0_), .Y(men_men_n461_));
  NO3        u0439(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n462_));
  NA2        u0440(.A(men_men_n267_), .B(men_men_n97_), .Y(men_men_n463_));
  NA2        u0441(.A(men_men_n463_), .B(men_men_n462_), .Y(men_men_n464_));
  NA2        u0442(.A(i_8_), .B(i_9_), .Y(men_men_n465_));
  NA2        u0443(.A(men_men_n285_), .B(men_men_n205_), .Y(men_men_n466_));
  OAI220     u0444(.A0(men_men_n466_), .A1(men_men_n465_), .B0(men_men_n464_), .B1(men_men_n461_), .Y(men_men_n467_));
  NO3        u0445(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n468_));
  NA3        u0446(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n469_));
  NO2        u0447(.A(men_men_n467_), .B(men_men_n460_), .Y(men_men_n470_));
  NA2        u0448(.A(men_men_n298_), .B(men_men_n108_), .Y(men_men_n471_));
  OR2        u0449(.A(men_men_n471_), .B(men_men_n207_), .Y(men_men_n472_));
  BUFFER     u0450(.A(men_men_n353_), .Y(men_men_n473_));
  OA220      u0451(.A0(men_men_n473_), .A1(men_men_n164_), .B0(men_men_n472_), .B1(men_men_n234_), .Y(men_men_n474_));
  NA2        u0452(.A(men_men_n96_), .B(i_13_), .Y(men_men_n475_));
  NA2        u0453(.A(men_men_n436_), .B(men_men_n385_), .Y(men_men_n476_));
  NO2        u0454(.A(i_2_), .B(i_13_), .Y(men_men_n477_));
  NA3        u0455(.A(men_men_n477_), .B(men_men_n163_), .C(men_men_n99_), .Y(men_men_n478_));
  OAI220     u0456(.A0(men_men_n478_), .A1(men_men_n239_), .B0(men_men_n476_), .B1(men_men_n475_), .Y(men_men_n479_));
  NO3        u0457(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n480_));
  NO2        u0458(.A(i_6_), .B(i_7_), .Y(men_men_n481_));
  NO2        u0459(.A(i_11_), .B(i_1_), .Y(men_men_n482_));
  OR2        u0460(.A(i_11_), .B(i_8_), .Y(men_men_n483_));
  NOi21      u0461(.An(i_2_), .B(i_7_), .Y(men_men_n484_));
  NAi31      u0462(.An(men_men_n483_), .B(men_men_n484_), .C(men_men_n1098_), .Y(men_men_n485_));
  NO2        u0463(.A(men_men_n423_), .B(i_6_), .Y(men_men_n486_));
  NA3        u0464(.A(men_men_n486_), .B(men_men_n454_), .C(men_men_n73_), .Y(men_men_n487_));
  NO2        u0465(.A(men_men_n487_), .B(men_men_n485_), .Y(men_men_n488_));
  NO2        u0466(.A(i_3_), .B(men_men_n192_), .Y(men_men_n489_));
  NO2        u0467(.A(i_6_), .B(i_10_), .Y(men_men_n490_));
  NA4        u0468(.A(men_men_n490_), .B(men_men_n315_), .C(men_men_n489_), .D(men_men_n239_), .Y(men_men_n491_));
  NO2        u0469(.A(men_men_n491_), .B(men_men_n157_), .Y(men_men_n492_));
  NA3        u0470(.A(men_men_n247_), .B(men_men_n173_), .C(men_men_n133_), .Y(men_men_n493_));
  NA2        u0471(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n494_));
  NO2        u0472(.A(men_men_n159_), .B(i_3_), .Y(men_men_n495_));
  NA3        u0473(.A(men_men_n397_), .B(men_men_n180_), .C(men_men_n150_), .Y(men_men_n496_));
  NA2        u0474(.A(men_men_n496_), .B(men_men_n493_), .Y(men_men_n497_));
  NO4        u0475(.A(men_men_n497_), .B(men_men_n492_), .C(men_men_n488_), .D(men_men_n479_), .Y(men_men_n498_));
  NA2        u0476(.A(men_men_n468_), .B(men_men_n393_), .Y(men_men_n499_));
  NO2        u0477(.A(men_men_n499_), .B(men_men_n226_), .Y(men_men_n500_));
  NAi21      u0478(.An(men_men_n217_), .B(men_men_n403_), .Y(men_men_n501_));
  NA2        u0479(.A(men_men_n339_), .B(men_men_n219_), .Y(men_men_n502_));
  NO2        u0480(.A(men_men_n26_), .B(i_5_), .Y(men_men_n503_));
  NO2        u0481(.A(i_0_), .B(men_men_n83_), .Y(men_men_n504_));
  NA3        u0482(.A(men_men_n504_), .B(men_men_n503_), .C(men_men_n143_), .Y(men_men_n505_));
  OR3        u0483(.A(i_4_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n506_));
  OAI220     u0484(.A0(men_men_n506_), .A1(men_men_n505_), .B0(men_men_n502_), .B1(men_men_n501_), .Y(men_men_n507_));
  NA2        u0485(.A(men_men_n27_), .B(i_10_), .Y(men_men_n508_));
  NA2        u0486(.A(men_men_n315_), .B(men_men_n240_), .Y(men_men_n509_));
  OAI220     u0487(.A0(men_men_n509_), .A1(men_men_n444_), .B0(men_men_n508_), .B1(men_men_n475_), .Y(men_men_n510_));
  NO3        u0488(.A(men_men_n510_), .B(men_men_n507_), .C(men_men_n500_), .Y(men_men_n511_));
  NA4        u0489(.A(men_men_n511_), .B(men_men_n498_), .C(men_men_n474_), .D(men_men_n470_), .Y(men_men_n512_));
  NA3        u0490(.A(men_men_n308_), .B(men_men_n177_), .C(men_men_n175_), .Y(men_men_n513_));
  OAI210     u0491(.A0(men_men_n304_), .A1(men_men_n1101_), .B0(men_men_n513_), .Y(men_men_n514_));
  AN2        u0492(.A(men_men_n289_), .B(men_men_n236_), .Y(men_men_n515_));
  NA2        u0493(.A(men_men_n515_), .B(men_men_n514_), .Y(men_men_n516_));
  NA2        u0494(.A(men_men_n123_), .B(men_men_n112_), .Y(men_men_n517_));
  AO220      u0495(.A0(men_men_n517_), .A1(men_men_n462_), .B0(men_men_n424_), .B1(i_6_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n315_), .B(men_men_n166_), .Y(men_men_n519_));
  OAI210     u0497(.A0(men_men_n519_), .A1(men_men_n234_), .B0(men_men_n309_), .Y(men_men_n520_));
  AOI220     u0498(.A0(men_men_n520_), .A1(i_7_), .B0(men_men_n518_), .B1(men_men_n311_), .Y(men_men_n521_));
  NA2        u0499(.A(men_men_n386_), .B(men_men_n227_), .Y(men_men_n522_));
  NA2        u0500(.A(men_men_n357_), .B(men_men_n71_), .Y(men_men_n523_));
  NA2        u0501(.A(men_men_n375_), .B(men_men_n367_), .Y(men_men_n524_));
  AO210      u0502(.A0(men_men_n523_), .A1(men_men_n522_), .B0(men_men_n524_), .Y(men_men_n525_));
  NO2        u0503(.A(men_men_n36_), .B(i_8_), .Y(men_men_n526_));
  AOI210     u0504(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n424_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n527_), .B(men_men_n525_), .Y(men_men_n528_));
  INV        u0506(.A(men_men_n528_), .Y(men_men_n529_));
  OAI210     u0507(.A0(i_8_), .A1(i_5_), .B0(men_men_n135_), .Y(men_men_n530_));
  AOI210     u0508(.A0(men_men_n193_), .A1(i_9_), .B0(men_men_n266_), .Y(men_men_n531_));
  NO2        u0509(.A(men_men_n531_), .B(men_men_n198_), .Y(men_men_n532_));
  OR2        u0510(.A(men_men_n182_), .B(i_4_), .Y(men_men_n533_));
  INV        u0511(.A(men_men_n533_), .Y(men_men_n534_));
  AOI220     u0512(.A0(men_men_n534_), .A1(men_men_n532_), .B0(men_men_n530_), .B1(men_men_n425_), .Y(men_men_n535_));
  NA4        u0513(.A(men_men_n535_), .B(men_men_n529_), .C(men_men_n521_), .D(men_men_n516_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n392_), .B(men_men_n298_), .Y(men_men_n537_));
  OAI210     u0515(.A0(men_men_n388_), .A1(i_2_), .B0(men_men_n537_), .Y(men_men_n538_));
  NO2        u0516(.A(i_12_), .B(men_men_n192_), .Y(men_men_n539_));
  NA2        u0517(.A(men_men_n539_), .B(men_men_n227_), .Y(men_men_n540_));
  NO3        u0518(.A(i_10_), .B(men_men_n540_), .C(men_men_n471_), .Y(men_men_n541_));
  NOi31      u0519(.An(men_men_n318_), .B(men_men_n423_), .C(men_men_n38_), .Y(men_men_n542_));
  OAI210     u0520(.A0(men_men_n542_), .A1(men_men_n541_), .B0(men_men_n538_), .Y(men_men_n543_));
  NO2        u0521(.A(i_8_), .B(i_7_), .Y(men_men_n544_));
  OAI210     u0522(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n545_));
  NA2        u0523(.A(men_men_n545_), .B(men_men_n225_), .Y(men_men_n546_));
  AOI220     u0524(.A0(men_men_n326_), .A1(men_men_n40_), .B0(men_men_n237_), .B1(men_men_n206_), .Y(men_men_n547_));
  OAI220     u0525(.A0(men_men_n547_), .A1(men_men_n533_), .B0(men_men_n546_), .B1(men_men_n244_), .Y(men_men_n548_));
  NA2        u0526(.A(men_men_n45_), .B(i_10_), .Y(men_men_n549_));
  NO2        u0527(.A(men_men_n549_), .B(i_6_), .Y(men_men_n550_));
  NA3        u0528(.A(men_men_n550_), .B(men_men_n548_), .C(men_men_n544_), .Y(men_men_n551_));
  AOI220     u0529(.A0(men_men_n436_), .A1(men_men_n326_), .B0(men_men_n249_), .B1(men_men_n246_), .Y(men_men_n552_));
  OAI220     u0530(.A0(men_men_n552_), .A1(i_12_), .B0(men_men_n475_), .B1(men_men_n134_), .Y(men_men_n553_));
  NA2        u0531(.A(men_men_n553_), .B(men_men_n266_), .Y(men_men_n554_));
  NOi31      u0532(.An(men_men_n293_), .B(men_men_n304_), .C(men_men_n1101_), .Y(men_men_n555_));
  NA3        u0533(.A(men_men_n308_), .B(men_men_n175_), .C(men_men_n96_), .Y(men_men_n556_));
  NO2        u0534(.A(men_men_n223_), .B(men_men_n45_), .Y(men_men_n557_));
  NO2        u0535(.A(men_men_n159_), .B(i_5_), .Y(men_men_n558_));
  NA2        u0536(.A(men_men_n558_), .B(men_men_n321_), .Y(men_men_n559_));
  OAI210     u0537(.A0(men_men_n559_), .A1(men_men_n557_), .B0(men_men_n556_), .Y(men_men_n560_));
  OAI210     u0538(.A0(men_men_n560_), .A1(men_men_n555_), .B0(men_men_n468_), .Y(men_men_n561_));
  NA4        u0539(.A(men_men_n561_), .B(men_men_n554_), .C(men_men_n551_), .D(men_men_n543_), .Y(men_men_n562_));
  NA3        u0540(.A(men_men_n219_), .B(men_men_n69_), .C(men_men_n45_), .Y(men_men_n563_));
  NA2        u0541(.A(men_men_n285_), .B(men_men_n81_), .Y(men_men_n564_));
  AOI210     u0542(.A0(men_men_n563_), .A1(men_men_n348_), .B0(men_men_n564_), .Y(men_men_n565_));
  NA2        u0543(.A(men_men_n299_), .B(men_men_n289_), .Y(men_men_n566_));
  NO2        u0544(.A(men_men_n566_), .B(men_men_n174_), .Y(men_men_n567_));
  NA2        u0545(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n568_));
  NA2        u0546(.A(men_men_n456_), .B(men_men_n223_), .Y(men_men_n569_));
  NO2        u0547(.A(men_men_n568_), .B(men_men_n569_), .Y(men_men_n570_));
  AOI210     u0548(.A0(men_men_n368_), .A1(men_men_n47_), .B0(men_men_n372_), .Y(men_men_n571_));
  NA2        u0549(.A(i_0_), .B(men_men_n49_), .Y(men_men_n572_));
  NA3        u0550(.A(men_men_n539_), .B(men_men_n276_), .C(men_men_n572_), .Y(men_men_n573_));
  NO2        u0551(.A(men_men_n571_), .B(men_men_n573_), .Y(men_men_n574_));
  NO4        u0552(.A(men_men_n574_), .B(men_men_n570_), .C(men_men_n567_), .D(men_men_n565_), .Y(men_men_n575_));
  NO4        u0553(.A(men_men_n252_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n576_));
  NO3        u0554(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n577_));
  NO2        u0555(.A(men_men_n235_), .B(men_men_n36_), .Y(men_men_n578_));
  AN2        u0556(.A(men_men_n578_), .B(men_men_n577_), .Y(men_men_n579_));
  OA210      u0557(.A0(men_men_n579_), .A1(men_men_n576_), .B0(men_men_n357_), .Y(men_men_n580_));
  NO2        u0558(.A(men_men_n423_), .B(i_1_), .Y(men_men_n581_));
  NOi31      u0559(.An(men_men_n581_), .B(men_men_n463_), .C(men_men_n71_), .Y(men_men_n582_));
  AN4        u0560(.A(men_men_n582_), .B(men_men_n420_), .C(men_men_n503_), .D(i_2_), .Y(men_men_n583_));
  NO2        u0561(.A(men_men_n434_), .B(men_men_n178_), .Y(men_men_n584_));
  NO3        u0562(.A(men_men_n584_), .B(men_men_n583_), .C(men_men_n580_), .Y(men_men_n585_));
  NOi21      u0563(.An(i_10_), .B(i_6_), .Y(men_men_n586_));
  NO2        u0564(.A(men_men_n83_), .B(men_men_n25_), .Y(men_men_n587_));
  AOI220     u0565(.A0(men_men_n285_), .A1(men_men_n587_), .B0(men_men_n276_), .B1(men_men_n586_), .Y(men_men_n588_));
  NO2        u0566(.A(men_men_n588_), .B(men_men_n461_), .Y(men_men_n589_));
  NO2        u0567(.A(men_men_n115_), .B(men_men_n23_), .Y(men_men_n590_));
  NA2        u0568(.A(men_men_n318_), .B(men_men_n166_), .Y(men_men_n591_));
  AOI220     u0569(.A0(men_men_n591_), .A1(men_men_n445_), .B0(men_men_n174_), .B1(men_men_n181_), .Y(men_men_n592_));
  NO2        u0570(.A(men_men_n197_), .B(men_men_n37_), .Y(men_men_n593_));
  NOi31      u0571(.An(men_men_n147_), .B(men_men_n593_), .C(men_men_n334_), .Y(men_men_n594_));
  NO3        u0572(.A(men_men_n594_), .B(men_men_n592_), .C(men_men_n589_), .Y(men_men_n595_));
  NO2        u0573(.A(men_men_n523_), .B(men_men_n382_), .Y(men_men_n596_));
  INV        u0574(.A(men_men_n321_), .Y(men_men_n597_));
  NO2        u0575(.A(i_12_), .B(men_men_n83_), .Y(men_men_n598_));
  NA3        u0576(.A(men_men_n598_), .B(men_men_n276_), .C(men_men_n572_), .Y(men_men_n599_));
  NA3        u0577(.A(men_men_n389_), .B(men_men_n285_), .C(men_men_n219_), .Y(men_men_n600_));
  AOI210     u0578(.A0(men_men_n600_), .A1(men_men_n599_), .B0(men_men_n597_), .Y(men_men_n601_));
  NA2        u0579(.A(men_men_n175_), .B(i_0_), .Y(men_men_n602_));
  NO3        u0580(.A(men_men_n602_), .B(i_8_), .C(men_men_n304_), .Y(men_men_n603_));
  OR2        u0581(.A(i_2_), .B(i_5_), .Y(men_men_n604_));
  OR2        u0582(.A(men_men_n604_), .B(men_men_n415_), .Y(men_men_n605_));
  INV        u0583(.A(men_men_n197_), .Y(men_men_n606_));
  AOI210     u0584(.A0(men_men_n606_), .A1(men_men_n605_), .B0(men_men_n501_), .Y(men_men_n607_));
  NO4        u0585(.A(men_men_n607_), .B(men_men_n603_), .C(men_men_n601_), .D(men_men_n596_), .Y(men_men_n608_));
  NA4        u0586(.A(men_men_n608_), .B(men_men_n595_), .C(men_men_n585_), .D(men_men_n575_), .Y(men_men_n609_));
  NO4        u0587(.A(men_men_n609_), .B(men_men_n562_), .C(men_men_n536_), .D(men_men_n512_), .Y(men_men_n610_));
  NA4        u0588(.A(men_men_n610_), .B(men_men_n453_), .C(men_men_n356_), .D(men_men_n314_), .Y(men7));
  NO2        u0589(.A(men_men_n92_), .B(men_men_n53_), .Y(men_men_n612_));
  NO2        u0590(.A(men_men_n108_), .B(men_men_n89_), .Y(men_men_n613_));
  NA2        u0591(.A(men_men_n387_), .B(men_men_n613_), .Y(men_men_n614_));
  NA2        u0592(.A(men_men_n490_), .B(men_men_n81_), .Y(men_men_n615_));
  NA2        u0593(.A(i_11_), .B(men_men_n192_), .Y(men_men_n616_));
  NA2        u0594(.A(men_men_n145_), .B(men_men_n616_), .Y(men_men_n617_));
  OAI210     u0595(.A0(men_men_n617_), .A1(men_men_n615_), .B0(men_men_n614_), .Y(men_men_n618_));
  NA3        u0596(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n619_));
  NO2        u0597(.A(men_men_n239_), .B(i_4_), .Y(men_men_n620_));
  NA2        u0598(.A(men_men_n620_), .B(i_8_), .Y(men_men_n621_));
  NA2        u0599(.A(i_2_), .B(men_men_n83_), .Y(men_men_n622_));
  OAI210     u0600(.A0(men_men_n86_), .A1(men_men_n202_), .B0(men_men_n203_), .Y(men_men_n623_));
  NO2        u0601(.A(i_7_), .B(men_men_n37_), .Y(men_men_n624_));
  NA2        u0602(.A(i_4_), .B(i_8_), .Y(men_men_n625_));
  AOI210     u0603(.A0(men_men_n625_), .A1(men_men_n308_), .B0(men_men_n624_), .Y(men_men_n626_));
  OAI220     u0604(.A0(men_men_n626_), .A1(men_men_n622_), .B0(men_men_n623_), .B1(i_13_), .Y(men_men_n627_));
  NO3        u0605(.A(men_men_n627_), .B(men_men_n618_), .C(men_men_n612_), .Y(men_men_n628_));
  INV        u0606(.A(men_men_n163_), .Y(men_men_n629_));
  OR2        u0607(.A(i_6_), .B(i_10_), .Y(men_men_n630_));
  NO2        u0608(.A(men_men_n630_), .B(men_men_n23_), .Y(men_men_n631_));
  OR3        u0609(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n632_));
  NO3        u0610(.A(men_men_n632_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n633_));
  INV        u0611(.A(men_men_n199_), .Y(men_men_n634_));
  NO2        u0612(.A(men_men_n633_), .B(men_men_n631_), .Y(men_men_n635_));
  OA220      u0613(.A0(men_men_n635_), .A1(men_men_n597_), .B0(men_men_n629_), .B1(men_men_n268_), .Y(men_men_n636_));
  AOI210     u0614(.A0(men_men_n636_), .A1(men_men_n628_), .B0(men_men_n61_), .Y(men_men_n637_));
  NOi21      u0615(.An(i_11_), .B(i_7_), .Y(men_men_n638_));
  AO210      u0616(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n639_));
  NO2        u0617(.A(men_men_n639_), .B(men_men_n638_), .Y(men_men_n640_));
  NA2        u0618(.A(men_men_n640_), .B(men_men_n206_), .Y(men_men_n641_));
  NA3        u0619(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n642_));
  NAi31      u0620(.An(men_men_n642_), .B(men_men_n216_), .C(i_11_), .Y(men_men_n643_));
  AOI210     u0621(.A0(men_men_n643_), .A1(men_men_n641_), .B0(men_men_n61_), .Y(men_men_n644_));
  NA2        u0622(.A(men_men_n85_), .B(men_men_n61_), .Y(men_men_n645_));
  OR2        u0623(.A(men_men_n645_), .B(men_men_n41_), .Y(men_men_n646_));
  NO3        u0624(.A(men_men_n260_), .B(men_men_n208_), .C(men_men_n616_), .Y(men_men_n647_));
  OAI210     u0625(.A0(men_men_n647_), .A1(men_men_n228_), .B0(men_men_n61_), .Y(men_men_n648_));
  NA2        u0626(.A(men_men_n416_), .B(men_men_n31_), .Y(men_men_n649_));
  OR2        u0627(.A(men_men_n208_), .B(men_men_n108_), .Y(men_men_n650_));
  NA2        u0628(.A(men_men_n650_), .B(men_men_n649_), .Y(men_men_n651_));
  NO2        u0629(.A(men_men_n61_), .B(i_9_), .Y(men_men_n652_));
  NO2        u0630(.A(men_men_n652_), .B(i_4_), .Y(men_men_n653_));
  NA2        u0631(.A(men_men_n653_), .B(men_men_n651_), .Y(men_men_n654_));
  NO2        u0632(.A(i_1_), .B(i_12_), .Y(men_men_n655_));
  NA3        u0633(.A(men_men_n655_), .B(men_men_n110_), .C(men_men_n24_), .Y(men_men_n656_));
  NA4        u0634(.A(men_men_n656_), .B(men_men_n654_), .C(men_men_n648_), .D(men_men_n646_), .Y(men_men_n657_));
  OAI210     u0635(.A0(men_men_n657_), .A1(men_men_n644_), .B0(i_6_), .Y(men_men_n658_));
  NO2        u0636(.A(men_men_n642_), .B(men_men_n108_), .Y(men_men_n659_));
  NA2        u0637(.A(men_men_n659_), .B(men_men_n598_), .Y(men_men_n660_));
  NO2        u0638(.A(i_6_), .B(i_11_), .Y(men_men_n661_));
  NA2        u0639(.A(men_men_n660_), .B(men_men_n464_), .Y(men_men_n662_));
  NO4        u0640(.A(men_men_n216_), .B(men_men_n129_), .C(i_13_), .D(men_men_n83_), .Y(men_men_n663_));
  NA2        u0641(.A(men_men_n663_), .B(men_men_n652_), .Y(men_men_n664_));
  NO3        u0642(.A(men_men_n630_), .B(men_men_n235_), .C(men_men_n23_), .Y(men_men_n665_));
  AOI210     u0643(.A0(i_1_), .A1(men_men_n261_), .B0(men_men_n665_), .Y(men_men_n666_));
  OAI210     u0644(.A0(men_men_n666_), .A1(men_men_n45_), .B0(men_men_n664_), .Y(men_men_n667_));
  NA3        u0645(.A(men_men_n544_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n668_));
  NA2        u0646(.A(men_men_n139_), .B(i_9_), .Y(men_men_n669_));
  NA3        u0647(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n670_));
  NO2        u0648(.A(men_men_n47_), .B(i_1_), .Y(men_men_n671_));
  NA3        u0649(.A(men_men_n671_), .B(men_men_n267_), .C(men_men_n45_), .Y(men_men_n672_));
  OAI220     u0650(.A0(men_men_n672_), .A1(men_men_n670_), .B0(men_men_n669_), .B1(men_men_n1095_), .Y(men_men_n673_));
  NA3        u0651(.A(men_men_n652_), .B(men_men_n321_), .C(i_6_), .Y(men_men_n674_));
  NO2        u0652(.A(men_men_n674_), .B(men_men_n23_), .Y(men_men_n675_));
  AOI210     u0653(.A0(men_men_n482_), .A1(men_men_n427_), .B0(men_men_n243_), .Y(men_men_n676_));
  NO2        u0654(.A(men_men_n676_), .B(men_men_n622_), .Y(men_men_n677_));
  NAi21      u0655(.An(men_men_n668_), .B(men_men_n91_), .Y(men_men_n678_));
  NA2        u0656(.A(men_men_n671_), .B(men_men_n267_), .Y(men_men_n679_));
  NO2        u0657(.A(i_11_), .B(men_men_n37_), .Y(men_men_n680_));
  NA2        u0658(.A(men_men_n680_), .B(men_men_n24_), .Y(men_men_n681_));
  OAI210     u0659(.A0(men_men_n681_), .A1(men_men_n679_), .B0(men_men_n678_), .Y(men_men_n682_));
  OR4        u0660(.A(men_men_n682_), .B(men_men_n677_), .C(men_men_n675_), .D(men_men_n673_), .Y(men_men_n683_));
  NO3        u0661(.A(men_men_n683_), .B(men_men_n667_), .C(men_men_n662_), .Y(men_men_n684_));
  NO2        u0662(.A(men_men_n239_), .B(men_men_n101_), .Y(men_men_n685_));
  NO2        u0663(.A(men_men_n685_), .B(men_men_n638_), .Y(men_men_n686_));
  NA2        u0664(.A(men_men_n686_), .B(i_1_), .Y(men_men_n687_));
  NO2        u0665(.A(men_men_n687_), .B(men_men_n632_), .Y(men_men_n688_));
  NO2        u0666(.A(men_men_n422_), .B(men_men_n83_), .Y(men_men_n689_));
  NA2        u0667(.A(men_men_n688_), .B(men_men_n47_), .Y(men_men_n690_));
  NA2        u0668(.A(i_3_), .B(men_men_n192_), .Y(men_men_n691_));
  NO2        u0669(.A(men_men_n691_), .B(men_men_n115_), .Y(men_men_n692_));
  AN2        u0670(.A(men_men_n692_), .B(men_men_n550_), .Y(men_men_n693_));
  NO2        u0671(.A(men_men_n118_), .B(men_men_n37_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n83_), .B(i_9_), .Y(men_men_n695_));
  NO2        u0673(.A(men_men_n695_), .B(men_men_n61_), .Y(men_men_n696_));
  NA2        u0674(.A(i_1_), .B(i_3_), .Y(men_men_n697_));
  NO2        u0675(.A(men_men_n465_), .B(men_men_n92_), .Y(men_men_n698_));
  INV        u0676(.A(men_men_n698_), .Y(men_men_n699_));
  NO2        u0677(.A(men_men_n699_), .B(men_men_n697_), .Y(men_men_n700_));
  NO2        u0678(.A(men_men_n700_), .B(men_men_n693_), .Y(men_men_n701_));
  NA4        u0679(.A(men_men_n701_), .B(men_men_n690_), .C(men_men_n684_), .D(men_men_n658_), .Y(men_men_n702_));
  NO3        u0680(.A(men_men_n483_), .B(i_3_), .C(i_7_), .Y(men_men_n703_));
  NOi21      u0681(.An(men_men_n703_), .B(i_10_), .Y(men_men_n704_));
  OA210      u0682(.A0(men_men_n704_), .A1(men_men_n247_), .B0(men_men_n83_), .Y(men_men_n705_));
  NA2        u0683(.A(men_men_n375_), .B(men_men_n374_), .Y(men_men_n706_));
  NA3        u0684(.A(men_men_n490_), .B(men_men_n526_), .C(men_men_n47_), .Y(men_men_n707_));
  NO3        u0685(.A(men_men_n484_), .B(men_men_n625_), .C(men_men_n83_), .Y(men_men_n708_));
  NA2        u0686(.A(men_men_n708_), .B(men_men_n25_), .Y(men_men_n709_));
  NA3        u0687(.A(men_men_n163_), .B(men_men_n81_), .C(men_men_n83_), .Y(men_men_n710_));
  NA4        u0688(.A(men_men_n710_), .B(men_men_n709_), .C(men_men_n707_), .D(men_men_n706_), .Y(men_men_n711_));
  OAI210     u0689(.A0(men_men_n711_), .A1(men_men_n705_), .B0(i_1_), .Y(men_men_n712_));
  AOI210     u0690(.A0(men_men_n267_), .A1(men_men_n97_), .B0(i_1_), .Y(men_men_n713_));
  NO2        u0691(.A(men_men_n373_), .B(i_2_), .Y(men_men_n714_));
  NA2        u0692(.A(men_men_n714_), .B(men_men_n713_), .Y(men_men_n715_));
  OAI210     u0693(.A0(men_men_n674_), .A1(men_men_n457_), .B0(men_men_n715_), .Y(men_men_n716_));
  INV        u0694(.A(men_men_n716_), .Y(men_men_n717_));
  AOI210     u0695(.A0(men_men_n717_), .A1(men_men_n712_), .B0(i_13_), .Y(men_men_n718_));
  OR2        u0696(.A(i_11_), .B(i_7_), .Y(men_men_n719_));
  NA3        u0697(.A(men_men_n719_), .B(men_men_n106_), .C(men_men_n139_), .Y(men_men_n720_));
  AOI220     u0698(.A0(men_men_n477_), .A1(men_men_n163_), .B0(i_2_), .B1(men_men_n139_), .Y(men_men_n721_));
  OAI210     u0699(.A0(men_men_n721_), .A1(men_men_n45_), .B0(men_men_n720_), .Y(men_men_n722_));
  AOI210     u0700(.A0(men_men_n670_), .A1(men_men_n53_), .B0(i_12_), .Y(men_men_n723_));
  INV        u0701(.A(men_men_n723_), .Y(men_men_n724_));
  NO2        u0702(.A(men_men_n484_), .B(men_men_n24_), .Y(men_men_n725_));
  AOI220     u0703(.A0(men_men_n725_), .A1(men_men_n689_), .B0(men_men_n247_), .B1(men_men_n132_), .Y(men_men_n726_));
  OAI220     u0704(.A0(men_men_n726_), .A1(men_men_n41_), .B0(men_men_n724_), .B1(men_men_n92_), .Y(men_men_n727_));
  AOI210     u0705(.A0(men_men_n722_), .A1(men_men_n336_), .B0(men_men_n727_), .Y(men_men_n728_));
  AOI220     u0706(.A0(i_12_), .A1(men_men_n70_), .B0(men_men_n389_), .B1(men_men_n671_), .Y(men_men_n729_));
  NO2        u0707(.A(men_men_n729_), .B(men_men_n244_), .Y(men_men_n730_));
  AOI210     u0708(.A0(men_men_n457_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n731_));
  NOi31      u0709(.An(men_men_n731_), .B(men_men_n615_), .C(men_men_n45_), .Y(men_men_n732_));
  NA2        u0710(.A(men_men_n128_), .B(i_13_), .Y(men_men_n733_));
  NO2        u0711(.A(men_men_n670_), .B(men_men_n115_), .Y(men_men_n734_));
  INV        u0712(.A(men_men_n734_), .Y(men_men_n735_));
  OAI220     u0713(.A0(men_men_n735_), .A1(men_men_n69_), .B0(men_men_n733_), .B1(men_men_n713_), .Y(men_men_n736_));
  NO3        u0714(.A(men_men_n69_), .B(men_men_n32_), .C(men_men_n101_), .Y(men_men_n737_));
  NA2        u0715(.A(men_men_n26_), .B(men_men_n192_), .Y(men_men_n738_));
  NA2        u0716(.A(men_men_n738_), .B(i_7_), .Y(men_men_n739_));
  NO3        u0717(.A(men_men_n484_), .B(men_men_n239_), .C(men_men_n83_), .Y(men_men_n740_));
  AOI210     u0718(.A0(men_men_n740_), .A1(men_men_n739_), .B0(men_men_n737_), .Y(men_men_n741_));
  AOI220     u0719(.A0(men_men_n389_), .A1(men_men_n671_), .B0(men_men_n91_), .B1(men_men_n102_), .Y(men_men_n742_));
  OAI220     u0720(.A0(men_men_n742_), .A1(men_men_n621_), .B0(men_men_n741_), .B1(men_men_n634_), .Y(men_men_n743_));
  NO4        u0721(.A(men_men_n743_), .B(men_men_n736_), .C(men_men_n732_), .D(men_men_n730_), .Y(men_men_n744_));
  OR2        u0722(.A(i_11_), .B(i_6_), .Y(men_men_n745_));
  NA3        u0723(.A(men_men_n620_), .B(men_men_n738_), .C(i_7_), .Y(men_men_n746_));
  AOI210     u0724(.A0(men_men_n746_), .A1(men_men_n735_), .B0(men_men_n745_), .Y(men_men_n747_));
  NA3        u0725(.A(men_men_n416_), .B(men_men_n624_), .C(men_men_n97_), .Y(men_men_n748_));
  NA2        u0726(.A(men_men_n661_), .B(i_13_), .Y(men_men_n749_));
  NA2        u0727(.A(men_men_n102_), .B(men_men_n738_), .Y(men_men_n750_));
  NAi21      u0728(.An(i_11_), .B(i_12_), .Y(men_men_n751_));
  NOi41      u0729(.An(men_men_n111_), .B(men_men_n751_), .C(i_13_), .D(men_men_n83_), .Y(men_men_n752_));
  NO3        u0730(.A(men_men_n484_), .B(men_men_n598_), .C(men_men_n625_), .Y(men_men_n753_));
  AOI220     u0731(.A0(men_men_n753_), .A1(men_men_n315_), .B0(men_men_n752_), .B1(men_men_n750_), .Y(men_men_n754_));
  NA3        u0732(.A(men_men_n754_), .B(men_men_n749_), .C(men_men_n748_), .Y(men_men_n755_));
  OAI210     u0733(.A0(men_men_n755_), .A1(men_men_n747_), .B0(men_men_n61_), .Y(men_men_n756_));
  NO2        u0734(.A(i_2_), .B(i_12_), .Y(men_men_n757_));
  NA2        u0735(.A(men_men_n372_), .B(men_men_n757_), .Y(men_men_n758_));
  NA2        u0736(.A(i_8_), .B(men_men_n25_), .Y(men_men_n759_));
  NO3        u0737(.A(men_men_n759_), .B(men_men_n387_), .C(men_men_n620_), .Y(men_men_n760_));
  NA2        u0738(.A(men_men_n760_), .B(men_men_n372_), .Y(men_men_n761_));
  NO2        u0739(.A(men_men_n129_), .B(i_2_), .Y(men_men_n762_));
  NA2        u0740(.A(men_men_n762_), .B(men_men_n655_), .Y(men_men_n763_));
  NA3        u0741(.A(men_men_n763_), .B(men_men_n761_), .C(men_men_n758_), .Y(men_men_n764_));
  NA3        u0742(.A(men_men_n764_), .B(men_men_n46_), .C(men_men_n227_), .Y(men_men_n765_));
  NA4        u0743(.A(men_men_n765_), .B(men_men_n756_), .C(men_men_n744_), .D(men_men_n728_), .Y(men_men_n766_));
  OR4        u0744(.A(men_men_n766_), .B(men_men_n718_), .C(men_men_n702_), .D(men_men_n637_), .Y(men5));
  AOI210     u0745(.A0(men_men_n686_), .A1(men_men_n270_), .B0(men_men_n425_), .Y(men_men_n768_));
  AN2        u0746(.A(men_men_n24_), .B(i_10_), .Y(men_men_n769_));
  NA3        u0747(.A(men_men_n769_), .B(men_men_n757_), .C(men_men_n108_), .Y(men_men_n770_));
  NO2        u0748(.A(men_men_n621_), .B(i_11_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n86_), .B(men_men_n771_), .Y(men_men_n772_));
  NA3        u0750(.A(men_men_n772_), .B(men_men_n770_), .C(men_men_n768_), .Y(men_men_n773_));
  NO3        u0751(.A(i_11_), .B(men_men_n239_), .C(i_13_), .Y(men_men_n774_));
  NO2        u0752(.A(men_men_n125_), .B(men_men_n23_), .Y(men_men_n775_));
  NA2        u0753(.A(i_12_), .B(i_8_), .Y(men_men_n776_));
  OAI210     u0754(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n776_), .Y(men_men_n777_));
  INV        u0755(.A(men_men_n456_), .Y(men_men_n778_));
  AOI220     u0756(.A0(men_men_n321_), .A1(men_men_n590_), .B0(men_men_n777_), .B1(men_men_n775_), .Y(men_men_n779_));
  INV        u0757(.A(men_men_n779_), .Y(men_men_n780_));
  NO2        u0758(.A(men_men_n780_), .B(men_men_n773_), .Y(men_men_n781_));
  INV        u0759(.A(men_men_n173_), .Y(men_men_n782_));
  INV        u0760(.A(men_men_n247_), .Y(men_men_n783_));
  OAI210     u0761(.A0(men_men_n714_), .A1(men_men_n458_), .B0(men_men_n111_), .Y(men_men_n784_));
  AOI210     u0762(.A0(men_men_n784_), .A1(men_men_n783_), .B0(men_men_n782_), .Y(men_men_n785_));
  NO2        u0763(.A(men_men_n465_), .B(men_men_n26_), .Y(men_men_n786_));
  NO2        u0764(.A(men_men_n786_), .B(men_men_n427_), .Y(men_men_n787_));
  NA2        u0765(.A(men_men_n787_), .B(i_2_), .Y(men_men_n788_));
  INV        u0766(.A(men_men_n788_), .Y(men_men_n789_));
  AOI210     u0767(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n423_), .Y(men_men_n790_));
  AOI210     u0768(.A0(men_men_n790_), .A1(men_men_n789_), .B0(men_men_n785_), .Y(men_men_n791_));
  NO2        u0769(.A(men_men_n189_), .B(men_men_n126_), .Y(men_men_n792_));
  OAI210     u0770(.A0(men_men_n792_), .A1(men_men_n775_), .B0(i_2_), .Y(men_men_n793_));
  NO2        u0771(.A(men_men_n793_), .B(men_men_n192_), .Y(men_men_n794_));
  OA210      u0772(.A0(men_men_n640_), .A1(men_men_n127_), .B0(i_13_), .Y(men_men_n795_));
  NA2        u0773(.A(men_men_n199_), .B(men_men_n202_), .Y(men_men_n796_));
  NA2        u0774(.A(men_men_n153_), .B(men_men_n616_), .Y(men_men_n797_));
  AOI210     u0775(.A0(men_men_n797_), .A1(men_men_n796_), .B0(men_men_n377_), .Y(men_men_n798_));
  AOI210     u0776(.A0(men_men_n208_), .A1(men_men_n149_), .B0(men_men_n526_), .Y(men_men_n799_));
  NA2        u0777(.A(men_men_n799_), .B(men_men_n427_), .Y(men_men_n800_));
  NO2        u0778(.A(men_men_n102_), .B(men_men_n45_), .Y(men_men_n801_));
  INV        u0779(.A(men_men_n305_), .Y(men_men_n802_));
  NA4        u0780(.A(men_men_n802_), .B(men_men_n308_), .C(men_men_n125_), .D(men_men_n43_), .Y(men_men_n803_));
  OAI210     u0781(.A0(men_men_n803_), .A1(men_men_n801_), .B0(men_men_n800_), .Y(men_men_n804_));
  NO4        u0782(.A(men_men_n804_), .B(men_men_n798_), .C(men_men_n795_), .D(men_men_n794_), .Y(men_men_n805_));
  NA2        u0783(.A(men_men_n590_), .B(men_men_n28_), .Y(men_men_n806_));
  NA2        u0784(.A(men_men_n774_), .B(men_men_n277_), .Y(men_men_n807_));
  NA2        u0785(.A(men_men_n807_), .B(men_men_n806_), .Y(men_men_n808_));
  NO2        u0786(.A(men_men_n60_), .B(i_12_), .Y(men_men_n809_));
  NO2        u0787(.A(men_men_n809_), .B(men_men_n127_), .Y(men_men_n810_));
  NO2        u0788(.A(men_men_n810_), .B(men_men_n616_), .Y(men_men_n811_));
  AOI220     u0789(.A0(men_men_n811_), .A1(men_men_n36_), .B0(men_men_n808_), .B1(men_men_n47_), .Y(men_men_n812_));
  NA4        u0790(.A(men_men_n812_), .B(men_men_n805_), .C(men_men_n791_), .D(men_men_n781_), .Y(men6));
  NO3        u0791(.A(men_men_n256_), .B(men_men_n310_), .C(i_1_), .Y(men_men_n814_));
  NO2        u0792(.A(men_men_n184_), .B(men_men_n140_), .Y(men_men_n815_));
  OAI210     u0793(.A0(men_men_n815_), .A1(men_men_n814_), .B0(men_men_n762_), .Y(men_men_n816_));
  NA3        u0794(.A(men_men_n393_), .B(men_men_n489_), .C(men_men_n69_), .Y(men_men_n817_));
  INV        u0795(.A(men_men_n817_), .Y(men_men_n818_));
  NO2        u0796(.A(men_men_n222_), .B(men_men_n494_), .Y(men_men_n819_));
  NO2        u0797(.A(i_11_), .B(i_9_), .Y(men_men_n820_));
  NO2        u0798(.A(men_men_n818_), .B(men_men_n331_), .Y(men_men_n821_));
  AO210      u0799(.A0(men_men_n821_), .A1(men_men_n816_), .B0(i_12_), .Y(men_men_n822_));
  NA2        u0800(.A(men_men_n378_), .B(men_men_n339_), .Y(men_men_n823_));
  NA2        u0801(.A(men_men_n598_), .B(men_men_n61_), .Y(men_men_n824_));
  NA2        u0802(.A(men_men_n704_), .B(men_men_n69_), .Y(men_men_n825_));
  NA4        u0803(.A(men_men_n645_), .B(men_men_n825_), .C(men_men_n824_), .D(men_men_n823_), .Y(men_men_n826_));
  INV        u0804(.A(men_men_n196_), .Y(men_men_n827_));
  AOI220     u0805(.A0(men_men_n827_), .A1(men_men_n820_), .B0(men_men_n826_), .B1(men_men_n71_), .Y(men_men_n828_));
  INV        u0806(.A(men_men_n330_), .Y(men_men_n829_));
  NA2        u0807(.A(men_men_n73_), .B(men_men_n132_), .Y(men_men_n830_));
  NO2        u0808(.A(men_men_n830_), .B(men_men_n829_), .Y(men_men_n831_));
  NO3        u0809(.A(men_men_n252_), .B(men_men_n133_), .C(i_9_), .Y(men_men_n832_));
  NA2        u0810(.A(men_men_n832_), .B(men_men_n809_), .Y(men_men_n833_));
  AOI210     u0811(.A0(men_men_n833_), .A1(men_men_n524_), .B0(men_men_n184_), .Y(men_men_n834_));
  NO2        u0812(.A(men_men_n32_), .B(i_11_), .Y(men_men_n835_));
  NA3        u0813(.A(men_men_n835_), .B(men_men_n481_), .C(men_men_n393_), .Y(men_men_n836_));
  NAi32      u0814(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n837_));
  AOI210     u0815(.A0(men_men_n745_), .A1(men_men_n84_), .B0(men_men_n837_), .Y(men_men_n838_));
  OAI210     u0816(.A0(men_men_n703_), .A1(men_men_n578_), .B0(men_men_n577_), .Y(men_men_n839_));
  NAi31      u0817(.An(men_men_n838_), .B(men_men_n839_), .C(men_men_n836_), .Y(men_men_n840_));
  OR3        u0818(.A(men_men_n840_), .B(men_men_n834_), .C(men_men_n831_), .Y(men_men_n841_));
  NO2        u0819(.A(men_men_n719_), .B(i_2_), .Y(men_men_n842_));
  NA2        u0820(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n843_));
  OAI210     u0821(.A0(men_men_n843_), .A1(men_men_n415_), .B0(men_men_n362_), .Y(men_men_n844_));
  NA2        u0822(.A(men_men_n844_), .B(men_men_n842_), .Y(men_men_n845_));
  AO220      u0823(.A0(men_men_n361_), .A1(men_men_n352_), .B0(men_men_n400_), .B1(men_men_n616_), .Y(men_men_n846_));
  NA3        u0824(.A(men_men_n846_), .B(men_men_n257_), .C(i_7_), .Y(men_men_n847_));
  OR2        u0825(.A(men_men_n640_), .B(men_men_n458_), .Y(men_men_n848_));
  NA3        u0826(.A(men_men_n848_), .B(men_men_n148_), .C(men_men_n67_), .Y(men_men_n849_));
  AO210      u0827(.A0(men_men_n499_), .A1(men_men_n778_), .B0(men_men_n36_), .Y(men_men_n850_));
  NA4        u0828(.A(men_men_n850_), .B(men_men_n849_), .C(men_men_n847_), .D(men_men_n845_), .Y(men_men_n851_));
  OAI210     u0829(.A0(i_6_), .A1(i_11_), .B0(men_men_n84_), .Y(men_men_n852_));
  AOI220     u0830(.A0(men_men_n852_), .A1(men_men_n577_), .B0(men_men_n819_), .B1(men_men_n739_), .Y(men_men_n853_));
  NA3        u0831(.A(men_men_n377_), .B(men_men_n240_), .C(men_men_n148_), .Y(men_men_n854_));
  NA2        u0832(.A(men_men_n400_), .B(men_men_n68_), .Y(men_men_n855_));
  NA4        u0833(.A(men_men_n855_), .B(men_men_n854_), .C(men_men_n853_), .D(men_men_n623_), .Y(men_men_n856_));
  AO210      u0834(.A0(men_men_n526_), .A1(men_men_n47_), .B0(men_men_n85_), .Y(men_men_n857_));
  NA3        u0835(.A(men_men_n857_), .B(men_men_n490_), .C(men_men_n219_), .Y(men_men_n858_));
  AOI210     u0836(.A0(men_men_n458_), .A1(men_men_n456_), .B0(men_men_n576_), .Y(men_men_n859_));
  NO2        u0837(.A(men_men_n630_), .B(men_men_n102_), .Y(men_men_n860_));
  OAI210     u0838(.A0(men_men_n860_), .A1(men_men_n112_), .B0(men_men_n414_), .Y(men_men_n861_));
  NA2        u0839(.A(men_men_n246_), .B(men_men_n47_), .Y(men_men_n862_));
  INV        u0840(.A(men_men_n605_), .Y(men_men_n863_));
  NA3        u0841(.A(men_men_n863_), .B(men_men_n330_), .C(i_7_), .Y(men_men_n864_));
  NA4        u0842(.A(men_men_n864_), .B(men_men_n861_), .C(men_men_n859_), .D(men_men_n858_), .Y(men_men_n865_));
  NO4        u0843(.A(men_men_n865_), .B(men_men_n856_), .C(men_men_n851_), .D(men_men_n841_), .Y(men_men_n866_));
  NA4        u0844(.A(men_men_n866_), .B(men_men_n828_), .C(men_men_n822_), .D(men_men_n383_), .Y(men3));
  NA2        u0845(.A(i_12_), .B(i_10_), .Y(men_men_n868_));
  NA2        u0846(.A(i_6_), .B(i_7_), .Y(men_men_n869_));
  NO2        u0847(.A(men_men_n869_), .B(i_0_), .Y(men_men_n870_));
  NO2        u0848(.A(i_11_), .B(men_men_n239_), .Y(men_men_n871_));
  OAI210     u0849(.A0(men_men_n870_), .A1(men_men_n293_), .B0(men_men_n871_), .Y(men_men_n872_));
  NO2        u0850(.A(men_men_n872_), .B(men_men_n192_), .Y(men_men_n873_));
  NO3        u0851(.A(men_men_n461_), .B(men_men_n89_), .C(men_men_n45_), .Y(men_men_n874_));
  OA210      u0852(.A0(men_men_n874_), .A1(men_men_n873_), .B0(men_men_n175_), .Y(men_men_n875_));
  NA3        u0853(.A(men_men_n854_), .B(men_men_n623_), .C(men_men_n376_), .Y(men_men_n876_));
  NA2        u0854(.A(men_men_n876_), .B(men_men_n40_), .Y(men_men_n877_));
  NO3        u0855(.A(men_men_n650_), .B(men_men_n465_), .C(men_men_n132_), .Y(men_men_n878_));
  NA2        u0856(.A(men_men_n416_), .B(men_men_n46_), .Y(men_men_n879_));
  AN2        u0857(.A(men_men_n463_), .B(men_men_n54_), .Y(men_men_n880_));
  NO2        u0858(.A(men_men_n880_), .B(men_men_n878_), .Y(men_men_n881_));
  AOI210     u0859(.A0(men_men_n881_), .A1(men_men_n877_), .B0(men_men_n49_), .Y(men_men_n882_));
  NO4        u0860(.A(men_men_n381_), .B(men_men_n386_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n883_));
  NA2        u0861(.A(men_men_n184_), .B(men_men_n586_), .Y(men_men_n884_));
  NOi21      u0862(.An(men_men_n884_), .B(men_men_n883_), .Y(men_men_n885_));
  NA2        u0863(.A(men_men_n731_), .B(men_men_n695_), .Y(men_men_n886_));
  NA2        u0864(.A(men_men_n337_), .B(men_men_n447_), .Y(men_men_n887_));
  OAI220     u0865(.A0(men_men_n887_), .A1(men_men_n886_), .B0(men_men_n885_), .B1(men_men_n61_), .Y(men_men_n888_));
  NOi21      u0866(.An(i_5_), .B(i_9_), .Y(men_men_n889_));
  NA2        u0867(.A(men_men_n889_), .B(men_men_n455_), .Y(men_men_n890_));
  AOI210     u0868(.A0(men_men_n267_), .A1(men_men_n482_), .B0(men_men_n708_), .Y(men_men_n891_));
  NO3        u0869(.A(men_men_n419_), .B(men_men_n267_), .C(men_men_n71_), .Y(men_men_n892_));
  INV        u0870(.A(men_men_n892_), .Y(men_men_n893_));
  OAI220     u0871(.A0(men_men_n893_), .A1(men_men_n1101_), .B0(men_men_n891_), .B1(men_men_n890_), .Y(men_men_n894_));
  NO4        u0872(.A(men_men_n894_), .B(men_men_n888_), .C(men_men_n882_), .D(men_men_n875_), .Y(men_men_n895_));
  NA2        u0873(.A(men_men_n184_), .B(men_men_n24_), .Y(men_men_n896_));
  NO2        u0874(.A(men_men_n694_), .B(men_men_n613_), .Y(men_men_n897_));
  NO2        u0875(.A(men_men_n897_), .B(men_men_n896_), .Y(men_men_n898_));
  NA2        u0876(.A(men_men_n315_), .B(men_men_n130_), .Y(men_men_n899_));
  NAi21      u0877(.An(men_men_n164_), .B(men_men_n447_), .Y(men_men_n900_));
  OAI220     u0878(.A0(men_men_n900_), .A1(men_men_n862_), .B0(men_men_n899_), .B1(men_men_n406_), .Y(men_men_n901_));
  NO2        u0879(.A(men_men_n901_), .B(men_men_n898_), .Y(men_men_n902_));
  NO2        u0880(.A(men_men_n393_), .B(men_men_n297_), .Y(men_men_n903_));
  NA2        u0881(.A(men_men_n903_), .B(men_men_n734_), .Y(men_men_n904_));
  NA2        u0882(.A(men_men_n587_), .B(i_0_), .Y(men_men_n905_));
  NO3        u0883(.A(men_men_n905_), .B(men_men_n388_), .C(men_men_n86_), .Y(men_men_n906_));
  NO4        u0884(.A(men_men_n604_), .B(men_men_n216_), .C(men_men_n423_), .D(men_men_n415_), .Y(men_men_n907_));
  AOI210     u0885(.A0(men_men_n907_), .A1(i_11_), .B0(men_men_n906_), .Y(men_men_n908_));
  INV        u0886(.A(men_men_n481_), .Y(men_men_n909_));
  AN2        u0887(.A(men_men_n96_), .B(men_men_n245_), .Y(men_men_n910_));
  NA2        u0888(.A(men_men_n774_), .B(men_men_n331_), .Y(men_men_n911_));
  AOI210     u0889(.A0(men_men_n490_), .A1(men_men_n86_), .B0(men_men_n56_), .Y(men_men_n912_));
  OAI220     u0890(.A0(men_men_n912_), .A1(men_men_n911_), .B0(men_men_n681_), .B1(men_men_n546_), .Y(men_men_n913_));
  NO2        u0891(.A(men_men_n254_), .B(men_men_n155_), .Y(men_men_n914_));
  NA2        u0892(.A(i_0_), .B(i_10_), .Y(men_men_n915_));
  NO4        u0893(.A(men_men_n115_), .B(men_men_n56_), .C(men_men_n691_), .D(i_5_), .Y(men_men_n916_));
  AO220      u0894(.A0(men_men_n916_), .A1(men_men_n1097_), .B0(men_men_n914_), .B1(i_6_), .Y(men_men_n917_));
  AOI220     u0895(.A0(men_men_n337_), .A1(men_men_n98_), .B0(men_men_n184_), .B1(men_men_n81_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n581_), .B(i_4_), .Y(men_men_n919_));
  NA2        u0897(.A(men_men_n187_), .B(men_men_n202_), .Y(men_men_n920_));
  OAI220     u0898(.A0(men_men_n920_), .A1(men_men_n911_), .B0(men_men_n919_), .B1(men_men_n918_), .Y(men_men_n921_));
  NO4        u0899(.A(men_men_n921_), .B(men_men_n917_), .C(men_men_n913_), .D(men_men_n910_), .Y(men_men_n922_));
  NA4        u0900(.A(men_men_n922_), .B(men_men_n908_), .C(men_men_n904_), .D(men_men_n902_), .Y(men_men_n923_));
  NO2        u0901(.A(men_men_n103_), .B(men_men_n37_), .Y(men_men_n924_));
  NA2        u0902(.A(i_11_), .B(i_9_), .Y(men_men_n925_));
  NO3        u0903(.A(i_12_), .B(men_men_n925_), .C(men_men_n622_), .Y(men_men_n926_));
  AO220      u0904(.A0(men_men_n926_), .A1(men_men_n924_), .B0(men_men_n269_), .B1(men_men_n85_), .Y(men_men_n927_));
  NO2        u0905(.A(men_men_n49_), .B(i_7_), .Y(men_men_n928_));
  NA2        u0906(.A(men_men_n397_), .B(men_men_n180_), .Y(men_men_n929_));
  NA2        u0907(.A(men_men_n929_), .B(men_men_n162_), .Y(men_men_n930_));
  NO2        u0908(.A(men_men_n925_), .B(men_men_n71_), .Y(men_men_n931_));
  NO2        u0909(.A(men_men_n176_), .B(i_0_), .Y(men_men_n932_));
  INV        u0910(.A(men_men_n932_), .Y(men_men_n933_));
  NA2        u0911(.A(men_men_n481_), .B(men_men_n233_), .Y(men_men_n934_));
  AOI210     u0912(.A0(men_men_n375_), .A1(men_men_n42_), .B0(men_men_n413_), .Y(men_men_n935_));
  OAI220     u0913(.A0(men_men_n935_), .A1(men_men_n890_), .B0(men_men_n934_), .B1(men_men_n933_), .Y(men_men_n936_));
  NO3        u0914(.A(men_men_n936_), .B(men_men_n930_), .C(men_men_n927_), .Y(men_men_n937_));
  NA2        u0915(.A(men_men_n680_), .B(men_men_n122_), .Y(men_men_n938_));
  NO2        u0916(.A(i_6_), .B(men_men_n938_), .Y(men_men_n939_));
  AOI210     u0917(.A0(men_men_n457_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n940_));
  NA2        u0918(.A(men_men_n173_), .B(men_men_n103_), .Y(men_men_n941_));
  NOi32      u0919(.An(men_men_n940_), .Bn(men_men_n187_), .C(men_men_n941_), .Y(men_men_n942_));
  NO2        u0920(.A(men_men_n1099_), .B(men_men_n879_), .Y(men_men_n943_));
  NO3        u0921(.A(men_men_n943_), .B(men_men_n942_), .C(men_men_n939_), .Y(men_men_n944_));
  NOi21      u0922(.An(i_7_), .B(i_5_), .Y(men_men_n945_));
  NOi31      u0923(.An(men_men_n945_), .B(i_0_), .C(men_men_n751_), .Y(men_men_n946_));
  NA3        u0924(.A(men_men_n946_), .B(men_men_n387_), .C(i_6_), .Y(men_men_n947_));
  OA210      u0925(.A0(men_men_n941_), .A1(men_men_n524_), .B0(men_men_n947_), .Y(men_men_n948_));
  NO3        u0926(.A(men_men_n409_), .B(men_men_n364_), .C(men_men_n360_), .Y(men_men_n949_));
  NO2        u0927(.A(men_men_n264_), .B(men_men_n322_), .Y(men_men_n950_));
  NO2        u0928(.A(men_men_n751_), .B(men_men_n259_), .Y(men_men_n951_));
  AOI210     u0929(.A0(men_men_n951_), .A1(men_men_n950_), .B0(men_men_n949_), .Y(men_men_n952_));
  NA4        u0930(.A(men_men_n952_), .B(men_men_n948_), .C(men_men_n944_), .D(men_men_n937_), .Y(men_men_n953_));
  NO2        u0931(.A(men_men_n896_), .B(men_men_n241_), .Y(men_men_n954_));
  AN2        u0932(.A(men_men_n336_), .B(men_men_n331_), .Y(men_men_n955_));
  NA2        u0933(.A(men_men_n954_), .B(i_10_), .Y(men_men_n956_));
  INV        u0934(.A(men_men_n868_), .Y(men_men_n957_));
  OA210      u0935(.A0(men_men_n481_), .A1(men_men_n225_), .B0(men_men_n480_), .Y(men_men_n958_));
  NA2        u0936(.A(men_men_n957_), .B(men_men_n931_), .Y(men_men_n959_));
  NO2        u0937(.A(men_men_n900_), .B(men_men_n909_), .Y(men_men_n960_));
  NO2        u0938(.A(men_men_n257_), .B(men_men_n47_), .Y(men_men_n961_));
  NA2        u0939(.A(men_men_n931_), .B(men_men_n308_), .Y(men_men_n962_));
  OAI210     u0940(.A0(men_men_n961_), .A1(men_men_n186_), .B0(men_men_n962_), .Y(men_men_n963_));
  AOI220     u0941(.A0(men_men_n963_), .A1(men_men_n481_), .B0(men_men_n960_), .B1(men_men_n71_), .Y(men_men_n964_));
  NA2        u0942(.A(men_men_n92_), .B(men_men_n45_), .Y(men_men_n965_));
  NO2        u0943(.A(men_men_n73_), .B(men_men_n776_), .Y(men_men_n966_));
  AOI220     u0944(.A0(men_men_n966_), .A1(men_men_n965_), .B0(men_men_n175_), .B1(men_men_n613_), .Y(men_men_n967_));
  NO2        u0945(.A(men_men_n967_), .B(men_men_n48_), .Y(men_men_n968_));
  NO3        u0946(.A(men_men_n604_), .B(men_men_n359_), .C(men_men_n24_), .Y(men_men_n969_));
  AOI210     u0947(.A0(men_men_n725_), .A1(men_men_n558_), .B0(men_men_n969_), .Y(men_men_n970_));
  NAi21      u0948(.An(i_9_), .B(i_5_), .Y(men_men_n971_));
  NO2        u0949(.A(men_men_n971_), .B(men_men_n409_), .Y(men_men_n972_));
  NO2        u0950(.A(men_men_n619_), .B(men_men_n105_), .Y(men_men_n973_));
  AOI220     u0951(.A0(men_men_n973_), .A1(i_0_), .B0(men_men_n972_), .B1(men_men_n640_), .Y(men_men_n974_));
  OAI220     u0952(.A0(men_men_n974_), .A1(men_men_n83_), .B0(men_men_n970_), .B1(men_men_n174_), .Y(men_men_n975_));
  NO3        u0953(.A(men_men_n975_), .B(men_men_n968_), .C(men_men_n528_), .Y(men_men_n976_));
  NA4        u0954(.A(men_men_n976_), .B(men_men_n964_), .C(men_men_n959_), .D(men_men_n956_), .Y(men_men_n977_));
  NO3        u0955(.A(men_men_n977_), .B(men_men_n953_), .C(men_men_n923_), .Y(men_men_n978_));
  NO2        u0956(.A(i_0_), .B(men_men_n751_), .Y(men_men_n979_));
  NA2        u0957(.A(men_men_n71_), .B(men_men_n45_), .Y(men_men_n980_));
  NA2        u0958(.A(men_men_n915_), .B(men_men_n980_), .Y(men_men_n981_));
  NO3        u0959(.A(men_men_n105_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n982_));
  AO220      u0960(.A0(men_men_n982_), .A1(men_men_n981_), .B0(men_men_n979_), .B1(men_men_n175_), .Y(men_men_n983_));
  AOI210     u0961(.A0(men_men_n824_), .A1(men_men_n706_), .B0(men_men_n941_), .Y(men_men_n984_));
  AOI210     u0962(.A0(men_men_n983_), .A1(men_men_n349_), .B0(men_men_n984_), .Y(men_men_n985_));
  NA2        u0963(.A(men_men_n762_), .B(men_men_n147_), .Y(men_men_n986_));
  INV        u0964(.A(men_men_n986_), .Y(men_men_n987_));
  NA3        u0965(.A(men_men_n987_), .B(men_men_n695_), .C(men_men_n71_), .Y(men_men_n988_));
  NO2        u0966(.A(men_men_n839_), .B(men_men_n409_), .Y(men_men_n989_));
  NA3        u0967(.A(men_men_n870_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n990_));
  NA2        u0968(.A(men_men_n871_), .B(i_9_), .Y(men_men_n991_));
  AOI210     u0969(.A0(men_men_n990_), .A1(men_men_n505_), .B0(men_men_n991_), .Y(men_men_n992_));
  OAI210     u0970(.A0(men_men_n246_), .A1(i_9_), .B0(men_men_n232_), .Y(men_men_n993_));
  AOI210     u0971(.A0(men_men_n993_), .A1(men_men_n905_), .B0(men_men_n155_), .Y(men_men_n994_));
  NO3        u0972(.A(men_men_n994_), .B(men_men_n992_), .C(men_men_n989_), .Y(men_men_n995_));
  NA3        u0973(.A(men_men_n995_), .B(men_men_n988_), .C(men_men_n985_), .Y(men_men_n996_));
  NA2        u0974(.A(men_men_n955_), .B(men_men_n377_), .Y(men_men_n997_));
  AOI210     u0975(.A0(men_men_n304_), .A1(men_men_n164_), .B0(men_men_n997_), .Y(men_men_n998_));
  NA3        u0976(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n999_));
  NA2        u0977(.A(men_men_n928_), .B(men_men_n495_), .Y(men_men_n1000_));
  AOI210     u0978(.A0(men_men_n999_), .A1(men_men_n164_), .B0(men_men_n1000_), .Y(men_men_n1001_));
  NO2        u0979(.A(men_men_n1001_), .B(men_men_n998_), .Y(men_men_n1002_));
  NA2        u0980(.A(men_men_n582_), .B(men_men_n73_), .Y(men_men_n1003_));
  NO3        u0981(.A(men_men_n210_), .B(men_men_n386_), .C(i_0_), .Y(men_men_n1004_));
  OAI210     u0982(.A0(men_men_n1004_), .A1(men_men_n74_), .B0(i_13_), .Y(men_men_n1005_));
  INV        u0983(.A(men_men_n219_), .Y(men_men_n1006_));
  OAI220     u0984(.A0(men_men_n540_), .A1(men_men_n140_), .B0(i_12_), .B1(men_men_n634_), .Y(men_men_n1007_));
  NA3        u0985(.A(men_men_n1007_), .B(men_men_n401_), .C(men_men_n1006_), .Y(men_men_n1008_));
  NA4        u0986(.A(men_men_n1008_), .B(men_men_n1005_), .C(men_men_n1003_), .D(men_men_n1002_), .Y(men_men_n1009_));
  NO2        u0987(.A(men_men_n244_), .B(men_men_n92_), .Y(men_men_n1010_));
  AOI210     u0988(.A0(men_men_n1010_), .A1(men_men_n979_), .B0(men_men_n109_), .Y(men_men_n1011_));
  AOI220     u0989(.A0(men_men_n945_), .A1(men_men_n495_), .B0(men_men_n870_), .B1(men_men_n165_), .Y(men_men_n1012_));
  NA2        u0990(.A(men_men_n352_), .B(men_men_n177_), .Y(men_men_n1013_));
  OA220      u0991(.A0(men_men_n1013_), .A1(men_men_n1012_), .B0(men_men_n1011_), .B1(i_5_), .Y(men_men_n1014_));
  AOI210     u0992(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n176_), .Y(men_men_n1015_));
  NA2        u0993(.A(men_men_n1015_), .B(men_men_n958_), .Y(men_men_n1016_));
  NA3        u0994(.A(men_men_n631_), .B(men_men_n184_), .C(men_men_n81_), .Y(men_men_n1017_));
  NA2        u0995(.A(men_men_n1017_), .B(men_men_n556_), .Y(men_men_n1018_));
  NA2        u0996(.A(men_men_n493_), .B(men_men_n478_), .Y(men_men_n1019_));
  NO2        u0997(.A(men_men_n1019_), .B(men_men_n1018_), .Y(men_men_n1020_));
  NA3        u0998(.A(men_men_n928_), .B(men_men_n293_), .C(men_men_n232_), .Y(men_men_n1021_));
  INV        u0999(.A(men_men_n1021_), .Y(men_men_n1022_));
  NA3        u1000(.A(men_men_n393_), .B(men_men_n338_), .C(men_men_n223_), .Y(men_men_n1023_));
  INV        u1001(.A(men_men_n1023_), .Y(men_men_n1024_));
  NOi31      u1002(.An(men_men_n392_), .B(men_men_n980_), .C(men_men_n241_), .Y(men_men_n1025_));
  NO3        u1003(.A(men_men_n1025_), .B(men_men_n1024_), .C(men_men_n1022_), .Y(men_men_n1026_));
  NA4        u1004(.A(men_men_n1026_), .B(men_men_n1020_), .C(men_men_n1016_), .D(men_men_n1014_), .Y(men_men_n1027_));
  INV        u1005(.A(men_men_n633_), .Y(men_men_n1028_));
  NO3        u1006(.A(men_men_n1028_), .B(men_men_n572_), .C(men_men_n346_), .Y(men_men_n1029_));
  INV        u1007(.A(men_men_n1029_), .Y(men_men_n1030_));
  NA3        u1008(.A(men_men_n308_), .B(i_5_), .C(men_men_n192_), .Y(men_men_n1031_));
  NAi31      u1009(.An(men_men_n243_), .B(men_men_n1031_), .C(men_men_n244_), .Y(men_men_n1032_));
  NO4        u1010(.A(men_men_n241_), .B(men_men_n210_), .C(i_0_), .D(i_12_), .Y(men_men_n1033_));
  AOI220     u1011(.A0(men_men_n1033_), .A1(men_men_n1032_), .B0(men_men_n818_), .B1(men_men_n177_), .Y(men_men_n1034_));
  AN2        u1012(.A(men_men_n915_), .B(men_men_n155_), .Y(men_men_n1035_));
  NO4        u1013(.A(men_men_n1035_), .B(i_12_), .C(men_men_n668_), .D(men_men_n132_), .Y(men_men_n1036_));
  NA2        u1014(.A(men_men_n1036_), .B(men_men_n219_), .Y(men_men_n1037_));
  NA3        u1015(.A(men_men_n98_), .B(men_men_n586_), .C(i_11_), .Y(men_men_n1038_));
  NO2        u1016(.A(men_men_n1038_), .B(men_men_n157_), .Y(men_men_n1039_));
  NA2        u1017(.A(men_men_n945_), .B(men_men_n477_), .Y(men_men_n1040_));
  OAI220     u1018(.A0(i_7_), .A1(men_men_n1031_), .B0(men_men_n1040_), .B1(men_men_n696_), .Y(men_men_n1041_));
  AOI210     u1019(.A0(men_men_n1041_), .A1(men_men_n932_), .B0(men_men_n1039_), .Y(men_men_n1042_));
  NA4        u1020(.A(men_men_n1042_), .B(men_men_n1037_), .C(men_men_n1034_), .D(men_men_n1030_), .Y(men_men_n1043_));
  NO4        u1021(.A(men_men_n1043_), .B(men_men_n1027_), .C(men_men_n1009_), .D(men_men_n996_), .Y(men_men_n1044_));
  NA2        u1022(.A(men_men_n835_), .B(men_men_n37_), .Y(men_men_n1045_));
  NA3        u1023(.A(men_men_n940_), .B(men_men_n372_), .C(i_5_), .Y(men_men_n1046_));
  NA3        u1024(.A(men_men_n1046_), .B(men_men_n1045_), .C(men_men_n629_), .Y(men_men_n1047_));
  NA2        u1025(.A(men_men_n1047_), .B(men_men_n206_), .Y(men_men_n1048_));
  AN2        u1026(.A(men_men_n719_), .B(men_men_n373_), .Y(men_men_n1049_));
  NA2        u1027(.A(men_men_n185_), .B(men_men_n187_), .Y(men_men_n1050_));
  AO210      u1028(.A0(men_men_n1049_), .A1(men_men_n33_), .B0(men_men_n1050_), .Y(men_men_n1051_));
  OAI210     u1029(.A0(men_men_n633_), .A1(men_men_n631_), .B0(men_men_n321_), .Y(men_men_n1052_));
  NAi31      u1030(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1053_));
  AOI210     u1031(.A0(men_men_n118_), .A1(men_men_n68_), .B0(men_men_n1053_), .Y(men_men_n1054_));
  NO2        u1032(.A(men_men_n1054_), .B(men_men_n665_), .Y(men_men_n1055_));
  NA3        u1033(.A(men_men_n1055_), .B(men_men_n1052_), .C(men_men_n1051_), .Y(men_men_n1056_));
  NO2        u1034(.A(men_men_n469_), .B(men_men_n267_), .Y(men_men_n1057_));
  NO4        u1035(.A(men_men_n235_), .B(men_men_n146_), .C(men_men_n697_), .D(men_men_n37_), .Y(men_men_n1058_));
  NO3        u1036(.A(men_men_n1058_), .B(men_men_n1057_), .C(men_men_n907_), .Y(men_men_n1059_));
  OAI210     u1037(.A0(men_men_n1038_), .A1(men_men_n149_), .B0(men_men_n1059_), .Y(men_men_n1060_));
  AOI210     u1038(.A0(men_men_n1056_), .A1(men_men_n49_), .B0(men_men_n1060_), .Y(men_men_n1061_));
  AOI210     u1039(.A0(men_men_n1061_), .A1(men_men_n1048_), .B0(men_men_n71_), .Y(men_men_n1062_));
  INV        u1040(.A(men_men_n579_), .Y(men_men_n1063_));
  NO2        u1041(.A(men_men_n1063_), .B(men_men_n782_), .Y(men_men_n1064_));
  OAI210     u1042(.A0(men_men_n78_), .A1(men_men_n53_), .B0(men_men_n108_), .Y(men_men_n1065_));
  NA2        u1043(.A(men_men_n1065_), .B(men_men_n74_), .Y(men_men_n1066_));
  AOI210     u1044(.A0(men_men_n1015_), .A1(men_men_n928_), .B0(men_men_n946_), .Y(men_men_n1067_));
  AOI210     u1045(.A0(men_men_n1067_), .A1(men_men_n1066_), .B0(men_men_n697_), .Y(men_men_n1068_));
  NA2        u1046(.A(men_men_n264_), .B(men_men_n55_), .Y(men_men_n1069_));
  AOI220     u1047(.A0(men_men_n1069_), .A1(men_men_n74_), .B0(men_men_n347_), .B1(men_men_n256_), .Y(men_men_n1070_));
  NO2        u1048(.A(men_men_n1070_), .B(men_men_n239_), .Y(men_men_n1071_));
  NA3        u1049(.A(men_men_n96_), .B(men_men_n310_), .C(men_men_n31_), .Y(men_men_n1072_));
  INV        u1050(.A(men_men_n1072_), .Y(men_men_n1073_));
  NO3        u1051(.A(men_men_n1073_), .B(men_men_n1071_), .C(men_men_n1068_), .Y(men_men_n1074_));
  OAI210     u1052(.A0(men_men_n269_), .A1(men_men_n160_), .B0(men_men_n86_), .Y(men_men_n1075_));
  NA3        u1053(.A(men_men_n786_), .B(men_men_n293_), .C(men_men_n78_), .Y(men_men_n1076_));
  AOI210     u1054(.A0(men_men_n1076_), .A1(men_men_n1075_), .B0(i_11_), .Y(men_men_n1077_));
  NA2        u1055(.A(men_men_n625_), .B(men_men_n216_), .Y(men_men_n1078_));
  OAI210     u1056(.A0(men_men_n1078_), .A1(men_men_n940_), .B0(men_men_n206_), .Y(men_men_n1079_));
  NA2        u1057(.A(men_men_n166_), .B(i_5_), .Y(men_men_n1080_));
  AOI210     u1058(.A0(men_men_n1079_), .A1(men_men_n796_), .B0(men_men_n1080_), .Y(men_men_n1081_));
  NO3        u1059(.A(men_men_n57_), .B(men_men_n56_), .C(i_4_), .Y(men_men_n1082_));
  OAI210     u1060(.A0(men_men_n950_), .A1(men_men_n310_), .B0(men_men_n1082_), .Y(men_men_n1083_));
  NO2        u1061(.A(men_men_n1083_), .B(men_men_n751_), .Y(men_men_n1084_));
  NO4        u1062(.A(men_men_n971_), .B(men_men_n483_), .C(men_men_n253_), .D(men_men_n252_), .Y(men_men_n1085_));
  NO2        u1063(.A(men_men_n1085_), .B(men_men_n576_), .Y(men_men_n1086_));
  INV        u1064(.A(men_men_n365_), .Y(men_men_n1087_));
  AOI210     u1065(.A0(men_men_n1087_), .A1(men_men_n1086_), .B0(men_men_n41_), .Y(men_men_n1088_));
  NO4        u1066(.A(men_men_n1088_), .B(men_men_n1084_), .C(men_men_n1081_), .D(men_men_n1077_), .Y(men_men_n1089_));
  OAI210     u1067(.A0(men_men_n1074_), .A1(i_4_), .B0(men_men_n1089_), .Y(men_men_n1090_));
  NO3        u1068(.A(men_men_n1090_), .B(men_men_n1064_), .C(men_men_n1062_), .Y(men_men_n1091_));
  NA4        u1069(.A(men_men_n1091_), .B(men_men_n1044_), .C(men_men_n978_), .D(men_men_n895_), .Y(men4));
  INV        u1070(.A(i_2_), .Y(men_men_n1095_));
  INV        u1071(.A(i_5_), .Y(men_men_n1096_));
  INV        u1072(.A(men_men_n915_), .Y(men_men_n1097_));
  INV        u1073(.A(i_3_), .Y(men_men_n1098_));
  INV        u1074(.A(men_men_n331_), .Y(men_men_n1099_));
  INV        u1075(.A(men_men_n393_), .Y(men_men_n1100_));
  INV        u1076(.A(i_5_), .Y(men_men_n1101_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule