// Benchmark "top" written by ABC on Thu Jun 20 14:00:11 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n42_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n112_, new_new_n113_, new_new_n115_, new_new_n116_,
    new_new_n117_, new_new_n118_, new_new_n119_, new_new_n120_,
    new_new_n121_, new_new_n122_, new_new_n123_, new_new_n124_,
    new_new_n125_, new_new_n126_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n283_, new_new_n284_, new_new_n285_,
    new_new_n286_, new_new_n287_, new_new_n288_, new_new_n289_,
    new_new_n290_, new_new_n291_, new_new_n292_, new_new_n293_,
    new_new_n294_, new_new_n295_, new_new_n296_, new_new_n297_,
    new_new_n298_, new_new_n299_, new_new_n300_, new_new_n301_,
    new_new_n302_, new_new_n303_, new_new_n304_, new_new_n305_,
    new_new_n306_, new_new_n307_, new_new_n308_, new_new_n309_,
    new_new_n310_, new_new_n311_, new_new_n312_, new_new_n313_,
    new_new_n314_, new_new_n315_, new_new_n316_, new_new_n317_,
    new_new_n318_, new_new_n319_, new_new_n320_, new_new_n321_,
    new_new_n322_, new_new_n323_, new_new_n324_, new_new_n325_,
    new_new_n326_, new_new_n327_, new_new_n328_, new_new_n329_,
    new_new_n330_, new_new_n331_, new_new_n332_, new_new_n333_,
    new_new_n334_, new_new_n335_, new_new_n336_, new_new_n337_,
    new_new_n338_, new_new_n339_, new_new_n340_, new_new_n341_,
    new_new_n342_, new_new_n343_, new_new_n344_, new_new_n345_,
    new_new_n346_, new_new_n347_, new_new_n348_, new_new_n349_,
    new_new_n350_, new_new_n351_, new_new_n352_, new_new_n353_,
    new_new_n354_, new_new_n355_, new_new_n356_, new_new_n357_,
    new_new_n358_, new_new_n359_, new_new_n360_, new_new_n361_,
    new_new_n362_, new_new_n363_, new_new_n364_, new_new_n365_,
    new_new_n366_, new_new_n367_, new_new_n368_, new_new_n369_,
    new_new_n370_, new_new_n371_, new_new_n372_, new_new_n374_,
    new_new_n375_, new_new_n376_, new_new_n377_, new_new_n378_,
    new_new_n379_, new_new_n380_, new_new_n381_, new_new_n382_,
    new_new_n383_, new_new_n384_, new_new_n385_, new_new_n386_,
    new_new_n387_, new_new_n388_, new_new_n389_, new_new_n390_,
    new_new_n391_, new_new_n392_, new_new_n393_, new_new_n394_,
    new_new_n395_, new_new_n396_, new_new_n397_, new_new_n398_,
    new_new_n399_, new_new_n400_, new_new_n401_, new_new_n403_,
    new_new_n404_, new_new_n405_, new_new_n406_, new_new_n407_,
    new_new_n408_, new_new_n409_, new_new_n410_, new_new_n411_,
    new_new_n412_, new_new_n413_, new_new_n414_, new_new_n415_,
    new_new_n416_, new_new_n417_, new_new_n418_, new_new_n419_,
    new_new_n420_, new_new_n421_, new_new_n422_, new_new_n423_,
    new_new_n424_, new_new_n425_, new_new_n426_, new_new_n427_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n514_, new_new_n515_,
    new_new_n516_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  BUFFER     g008(.A(i_11_), .Y(new_new_n31_));
  BUFFER     g009(.A(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n35_), .Y(ori1));
  INV        g019(.A(i_11_), .Y(new_new_n42_));
  NO2        g020(.A(new_new_n42_), .B(i_6_), .Y(new_new_n43_));
  INV        g021(.A(i_2_), .Y(new_new_n44_));
  INV        g022(.A(i_5_), .Y(new_new_n45_));
  NO2        g023(.A(i_7_), .B(i_10_), .Y(new_new_n46_));
  AOI210     g024(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n46_), .Y(new_new_n47_));
  NA2        g025(.A(i_0_), .B(i_2_), .Y(new_new_n48_));
  NA2        g026(.A(i_7_), .B(i_9_), .Y(new_new_n49_));
  NO2        g027(.A(new_new_n49_), .B(new_new_n48_), .Y(new_new_n50_));
  NA2        g028(.A(i_2_), .B(new_new_n43_), .Y(new_new_n51_));
  NO2        g029(.A(i_1_), .B(i_6_), .Y(new_new_n52_));
  NA2        g030(.A(i_8_), .B(i_7_), .Y(new_new_n53_));
  NAi21      g031(.An(i_2_), .B(i_7_), .Y(new_new_n54_));
  INV        g032(.A(i_1_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n55_), .B(i_6_), .Y(new_new_n56_));
  NA3        g034(.A(new_new_n56_), .B(new_new_n54_), .C(new_new_n31_), .Y(new_new_n57_));
  NA2        g035(.A(i_1_), .B(i_10_), .Y(new_new_n58_));
  NO2        g036(.A(new_new_n58_), .B(i_6_), .Y(new_new_n59_));
  NAi21      g037(.An(new_new_n59_), .B(new_new_n57_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n47_), .B(i_2_), .Y(new_new_n61_));
  AOI210     g039(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_6_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(new_new_n25_), .Y(new_new_n64_));
  INV        g042(.A(i_0_), .Y(new_new_n65_));
  NA2        g043(.A(i_5_), .B(i_9_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(new_new_n65_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(new_new_n64_), .Y(new_new_n68_));
  OAI210     g046(.A0(new_new_n62_), .A1(new_new_n61_), .B0(new_new_n68_), .Y(new_new_n69_));
  OAI210     g047(.A0(new_new_n69_), .A1(new_new_n60_), .B0(i_0_), .Y(new_new_n70_));
  NA2        g048(.A(i_12_), .B(i_5_), .Y(new_new_n71_));
  NO2        g049(.A(i_3_), .B(i_7_), .Y(new_new_n72_));
  INV        g050(.A(i_6_), .Y(new_new_n73_));
  NO2        g051(.A(i_2_), .B(i_7_), .Y(new_new_n74_));
  INV        g052(.A(new_new_n74_), .Y(new_new_n75_));
  NA2        g053(.A(i_1_), .B(new_new_n75_), .Y(new_new_n76_));
  NAi21      g054(.An(i_6_), .B(i_10_), .Y(new_new_n77_));
  NA2        g055(.A(i_6_), .B(i_9_), .Y(new_new_n78_));
  AOI210     g056(.A0(new_new_n78_), .A1(new_new_n77_), .B0(new_new_n55_), .Y(new_new_n79_));
  NA2        g057(.A(i_2_), .B(i_6_), .Y(new_new_n80_));
  INV        g058(.A(new_new_n79_), .Y(new_new_n81_));
  AOI210     g059(.A0(new_new_n81_), .A1(new_new_n76_), .B0(new_new_n71_), .Y(new_new_n82_));
  AN3        g060(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n83_));
  NAi21      g061(.An(i_6_), .B(i_11_), .Y(new_new_n84_));
  INV        g062(.A(i_7_), .Y(new_new_n85_));
  NA2        g063(.A(new_new_n44_), .B(new_new_n85_), .Y(new_new_n86_));
  NO2        g064(.A(i_0_), .B(i_5_), .Y(new_new_n87_));
  NO2        g065(.A(new_new_n87_), .B(new_new_n73_), .Y(new_new_n88_));
  NA2        g066(.A(i_12_), .B(i_3_), .Y(new_new_n89_));
  NA3        g067(.A(i_12_), .B(new_new_n88_), .C(new_new_n86_), .Y(new_new_n90_));
  NAi21      g068(.An(i_7_), .B(i_11_), .Y(new_new_n91_));
  AN2        g069(.A(i_2_), .B(i_10_), .Y(new_new_n92_));
  NO2        g070(.A(new_new_n92_), .B(i_7_), .Y(new_new_n93_));
  BUFFER     g071(.A(new_new_n71_), .Y(new_new_n94_));
  NA2        g072(.A(i_12_), .B(i_7_), .Y(new_new_n95_));
  NO2        g073(.A(new_new_n55_), .B(new_new_n26_), .Y(new_new_n96_));
  NA2        g074(.A(i_11_), .B(i_12_), .Y(new_new_n97_));
  NA2        g075(.A(new_new_n97_), .B(new_new_n90_), .Y(new_new_n98_));
  BUFFER     g076(.A(i_1_), .Y(new_new_n99_));
  NA2        g077(.A(new_new_n99_), .B(i_11_), .Y(new_new_n100_));
  NA2        g078(.A(new_new_n85_), .B(new_new_n37_), .Y(new_new_n101_));
  NA2        g079(.A(i_7_), .B(new_new_n25_), .Y(new_new_n102_));
  NA2        g080(.A(new_new_n102_), .B(new_new_n101_), .Y(new_new_n103_));
  NO2        g081(.A(new_new_n103_), .B(new_new_n44_), .Y(new_new_n104_));
  NA2        g082(.A(new_new_n78_), .B(new_new_n77_), .Y(new_new_n105_));
  NAi21      g083(.An(i_3_), .B(i_8_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n105_), .B(new_new_n104_), .Y(new_new_n107_));
  NO2        g085(.A(i_6_), .B(i_5_), .Y(new_new_n108_));
  NO2        g086(.A(new_new_n107_), .B(new_new_n100_), .Y(new_new_n109_));
  NO3        g087(.A(new_new_n109_), .B(new_new_n98_), .C(new_new_n82_), .Y(new_new_n110_));
  NA3        g088(.A(new_new_n110_), .B(new_new_n70_), .C(new_new_n51_), .Y(ori2));
  NO2        g089(.A(new_new_n55_), .B(new_new_n37_), .Y(new_new_n112_));
  INV        g090(.A(new_new_n112_), .Y(new_new_n113_));
  NA4        g091(.A(new_new_n113_), .B(new_new_n68_), .C(new_new_n61_), .D(new_new_n30_), .Y(ori0));
  NO2        g092(.A(i_12_), .B(i_13_), .Y(new_new_n115_));
  NAi21      g093(.An(i_5_), .B(i_11_), .Y(new_new_n116_));
  NO2        g094(.A(i_0_), .B(i_1_), .Y(new_new_n117_));
  NA2        g095(.A(i_1_), .B(i_5_), .Y(new_new_n118_));
  OR2        g096(.A(i_0_), .B(i_1_), .Y(new_new_n119_));
  NOi21      g097(.An(i_4_), .B(i_10_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(new_new_n40_), .Y(new_new_n121_));
  NOi21      g099(.An(i_4_), .B(i_9_), .Y(new_new_n122_));
  NOi21      g100(.An(i_11_), .B(i_13_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n122_), .Y(new_new_n124_));
  NO2        g102(.A(new_new_n65_), .B(i_5_), .Y(new_new_n125_));
  NO2        g103(.A(i_2_), .B(i_1_), .Y(new_new_n126_));
  NAi21      g104(.An(i_4_), .B(i_12_), .Y(new_new_n127_));
  INV        g105(.A(i_8_), .Y(new_new_n128_));
  NO2        g106(.A(i_3_), .B(i_8_), .Y(new_new_n129_));
  NO3        g107(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n130_));
  NO2        g108(.A(new_new_n87_), .B(new_new_n52_), .Y(new_new_n131_));
  NO2        g109(.A(i_13_), .B(i_9_), .Y(new_new_n132_));
  NAi21      g110(.An(i_12_), .B(i_3_), .Y(new_new_n133_));
  NO2        g111(.A(new_new_n42_), .B(i_5_), .Y(new_new_n134_));
  NA3        g112(.A(i_13_), .B(new_new_n128_), .C(i_10_), .Y(new_new_n135_));
  NA2        g113(.A(i_0_), .B(i_5_), .Y(new_new_n136_));
  NAi31      g114(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n137_));
  NO2        g115(.A(new_new_n65_), .B(new_new_n26_), .Y(new_new_n138_));
  NO2        g116(.A(new_new_n44_), .B(new_new_n55_), .Y(new_new_n139_));
  INV        g117(.A(i_13_), .Y(new_new_n140_));
  NO2        g118(.A(i_12_), .B(new_new_n140_), .Y(new_new_n141_));
  OR2        g119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  INV        g120(.A(i_12_), .Y(new_new_n143_));
  NO2        g121(.A(new_new_n42_), .B(new_new_n143_), .Y(new_new_n144_));
  NO3        g122(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n145_));
  NA2        g123(.A(i_2_), .B(i_1_), .Y(new_new_n146_));
  NAi21      g124(.An(i_4_), .B(i_3_), .Y(new_new_n147_));
  NO2        g125(.A(i_0_), .B(i_6_), .Y(new_new_n148_));
  NOi41      g126(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n149_));
  NO2        g127(.A(i_11_), .B(new_new_n140_), .Y(new_new_n150_));
  NOi21      g128(.An(i_1_), .B(i_6_), .Y(new_new_n151_));
  NAi21      g129(.An(i_3_), .B(i_7_), .Y(new_new_n152_));
  NA2        g130(.A(new_new_n143_), .B(i_9_), .Y(new_new_n153_));
  OR4        g131(.A(new_new_n153_), .B(new_new_n152_), .C(new_new_n151_), .D(new_new_n125_), .Y(new_new_n154_));
  NA2        g132(.A(new_new_n65_), .B(i_5_), .Y(new_new_n155_));
  NA2        g133(.A(i_3_), .B(i_9_), .Y(new_new_n156_));
  NAi21      g134(.An(i_7_), .B(i_10_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n157_), .B(new_new_n156_), .Y(new_new_n158_));
  NA3        g136(.A(new_new_n158_), .B(new_new_n155_), .C(new_new_n56_), .Y(new_new_n159_));
  NA2        g137(.A(new_new_n159_), .B(new_new_n154_), .Y(new_new_n160_));
  NA2        g138(.A(new_new_n160_), .B(new_new_n150_), .Y(new_new_n161_));
  NA2        g139(.A(i_12_), .B(i_6_), .Y(new_new_n162_));
  OR2        g140(.A(i_13_), .B(i_9_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n147_), .B(i_2_), .Y(new_new_n164_));
  NA2        g142(.A(new_new_n150_), .B(i_9_), .Y(new_new_n165_));
  NO3        g143(.A(i_11_), .B(new_new_n140_), .C(new_new_n25_), .Y(new_new_n166_));
  NO3        g144(.A(i_12_), .B(new_new_n140_), .C(new_new_n37_), .Y(new_new_n167_));
  AN2        g145(.A(i_3_), .B(i_10_), .Y(new_new_n168_));
  NO2        g146(.A(i_5_), .B(new_new_n37_), .Y(new_new_n169_));
  NO3        g147(.A(new_new_n42_), .B(i_13_), .C(i_9_), .Y(new_new_n170_));
  NO2        g148(.A(i_2_), .B(i_3_), .Y(new_new_n171_));
  NO2        g149(.A(i_12_), .B(i_10_), .Y(new_new_n172_));
  NOi21      g150(.An(i_5_), .B(i_0_), .Y(new_new_n173_));
  NO2        g151(.A(i_1_), .B(i_7_), .Y(new_new_n174_));
  NOi21      g152(.An(new_new_n118_), .B(new_new_n88_), .Y(new_new_n175_));
  NO2        g153(.A(new_new_n175_), .B(new_new_n102_), .Y(new_new_n176_));
  NA2        g154(.A(new_new_n176_), .B(i_3_), .Y(new_new_n177_));
  NO2        g155(.A(new_new_n128_), .B(i_9_), .Y(new_new_n178_));
  NA2        g156(.A(new_new_n178_), .B(new_new_n131_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n179_), .B(new_new_n44_), .Y(new_new_n180_));
  INV        g158(.A(new_new_n180_), .Y(new_new_n181_));
  AOI210     g159(.A0(new_new_n181_), .A1(new_new_n177_), .B0(new_new_n121_), .Y(new_new_n182_));
  INV        g160(.A(new_new_n182_), .Y(new_new_n183_));
  NOi32      g161(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n184_));
  INV        g162(.A(new_new_n184_), .Y(new_new_n185_));
  NOi32      g163(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n186_));
  NAi21      g164(.An(i_6_), .B(i_1_), .Y(new_new_n187_));
  NA3        g165(.A(new_new_n187_), .B(new_new_n186_), .C(new_new_n44_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n188_), .B(i_0_), .Y(new_new_n189_));
  NO2        g167(.A(i_1_), .B(new_new_n85_), .Y(new_new_n190_));
  NAi21      g168(.An(i_3_), .B(i_4_), .Y(new_new_n191_));
  NO2        g169(.A(new_new_n191_), .B(i_9_), .Y(new_new_n192_));
  AN2        g170(.A(i_6_), .B(i_7_), .Y(new_new_n193_));
  OAI210     g171(.A0(new_new_n193_), .A1(new_new_n190_), .B0(new_new_n192_), .Y(new_new_n194_));
  NA2        g172(.A(i_2_), .B(i_7_), .Y(new_new_n195_));
  NO2        g173(.A(new_new_n191_), .B(i_10_), .Y(new_new_n196_));
  NA3        g174(.A(new_new_n196_), .B(new_new_n195_), .C(new_new_n148_), .Y(new_new_n197_));
  AOI210     g175(.A0(new_new_n197_), .A1(new_new_n194_), .B0(new_new_n125_), .Y(new_new_n198_));
  AOI210     g176(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n199_));
  OAI210     g177(.A0(new_new_n199_), .A1(new_new_n126_), .B0(new_new_n196_), .Y(new_new_n200_));
  AOI220     g178(.A0(new_new_n196_), .A1(new_new_n174_), .B0(new_new_n145_), .B1(new_new_n126_), .Y(new_new_n201_));
  AOI210     g179(.A0(new_new_n201_), .A1(new_new_n200_), .B0(i_5_), .Y(new_new_n202_));
  NO3        g180(.A(new_new_n202_), .B(new_new_n198_), .C(new_new_n189_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n203_), .B(new_new_n185_), .Y(new_new_n204_));
  AN2        g182(.A(i_12_), .B(i_5_), .Y(new_new_n205_));
  NO2        g183(.A(i_5_), .B(i_10_), .Y(new_new_n206_));
  NO3        g184(.A(new_new_n73_), .B(new_new_n45_), .C(i_9_), .Y(new_new_n207_));
  NO2        g185(.A(i_11_), .B(i_12_), .Y(new_new_n208_));
  NAi21      g186(.An(i_13_), .B(i_0_), .Y(new_new_n209_));
  NO3        g187(.A(i_1_), .B(i_12_), .C(new_new_n73_), .Y(new_new_n210_));
  NO2        g188(.A(i_0_), .B(i_11_), .Y(new_new_n211_));
  AN2        g189(.A(i_1_), .B(i_6_), .Y(new_new_n212_));
  NAi21      g190(.An(i_9_), .B(i_4_), .Y(new_new_n213_));
  OR2        g191(.A(i_13_), .B(i_10_), .Y(new_new_n214_));
  NO3        g192(.A(new_new_n214_), .B(new_new_n97_), .C(new_new_n213_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n216_));
  NA2        g194(.A(new_new_n167_), .B(new_new_n216_), .Y(new_new_n217_));
  NO2        g195(.A(new_new_n217_), .B(new_new_n175_), .Y(new_new_n218_));
  NA2        g196(.A(new_new_n128_), .B(i_10_), .Y(new_new_n219_));
  NA3        g197(.A(new_new_n155_), .B(new_new_n56_), .C(i_2_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n221_));
  INV        g199(.A(new_new_n221_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n222_), .B(new_new_n165_), .Y(new_new_n223_));
  NO3        g201(.A(new_new_n223_), .B(new_new_n218_), .C(new_new_n204_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n65_), .B(i_13_), .Y(new_new_n225_));
  NO2        g203(.A(i_10_), .B(i_9_), .Y(new_new_n226_));
  NAi21      g204(.An(i_12_), .B(i_8_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(i_3_), .Y(new_new_n228_));
  NA2        g206(.A(new_new_n162_), .B(new_new_n84_), .Y(new_new_n229_));
  NA2        g207(.A(i_8_), .B(i_9_), .Y(new_new_n230_));
  NA2        g208(.A(new_new_n167_), .B(new_new_n131_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n231_), .B(new_new_n230_), .Y(new_new_n232_));
  NA3        g210(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n233_));
  NA4        g211(.A(new_new_n116_), .B(new_new_n96_), .C(new_new_n71_), .D(new_new_n23_), .Y(new_new_n234_));
  NO2        g212(.A(new_new_n234_), .B(new_new_n233_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n235_), .B(new_new_n232_), .Y(new_new_n236_));
  NA2        g214(.A(new_new_n83_), .B(i_13_), .Y(new_new_n237_));
  NO3        g215(.A(i_4_), .B(new_new_n45_), .C(i_8_), .Y(new_new_n238_));
  NO2        g216(.A(i_6_), .B(i_7_), .Y(new_new_n239_));
  NO2        g217(.A(i_11_), .B(i_1_), .Y(new_new_n240_));
  NOi21      g218(.An(i_2_), .B(i_7_), .Y(new_new_n241_));
  NO2        g219(.A(i_6_), .B(i_10_), .Y(new_new_n242_));
  NA3        g220(.A(new_new_n149_), .B(new_new_n123_), .C(new_new_n108_), .Y(new_new_n243_));
  NA2        g221(.A(new_new_n44_), .B(new_new_n42_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n119_), .B(i_3_), .Y(new_new_n245_));
  NAi31      g223(.An(new_new_n244_), .B(new_new_n245_), .C(new_new_n141_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n246_), .B(new_new_n243_), .Y(new_new_n247_));
  INV        g225(.A(new_new_n247_), .Y(new_new_n248_));
  NAi21      g226(.An(new_new_n135_), .B(new_new_n208_), .Y(new_new_n249_));
  NA2        g227(.A(new_new_n27_), .B(i_10_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n170_), .B(new_new_n145_), .Y(new_new_n251_));
  OAI220     g229(.A0(new_new_n251_), .A1(new_new_n220_), .B0(new_new_n250_), .B1(new_new_n237_), .Y(new_new_n252_));
  INV        g230(.A(new_new_n252_), .Y(new_new_n253_));
  NA3        g231(.A(new_new_n253_), .B(new_new_n248_), .C(new_new_n236_), .Y(new_new_n254_));
  NA2        g232(.A(new_new_n205_), .B(new_new_n140_), .Y(new_new_n255_));
  NA2        g233(.A(new_new_n193_), .B(new_new_n186_), .Y(new_new_n256_));
  OR2        g234(.A(new_new_n255_), .B(new_new_n256_), .Y(new_new_n257_));
  AOI210     g235(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n215_), .Y(new_new_n258_));
  NA2        g236(.A(new_new_n258_), .B(new_new_n257_), .Y(new_new_n259_));
  NO2        g237(.A(i_12_), .B(new_new_n128_), .Y(new_new_n260_));
  NA2        g238(.A(new_new_n42_), .B(i_10_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n119_), .B(i_5_), .Y(new_new_n262_));
  NA3        g240(.A(new_new_n136_), .B(new_new_n63_), .C(new_new_n42_), .Y(new_new_n263_));
  NA2        g241(.A(new_new_n167_), .B(new_new_n72_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n263_), .B(new_new_n264_), .Y(new_new_n265_));
  NA2        g243(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n266_));
  NA2        g244(.A(new_new_n226_), .B(i_4_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n266_), .B(new_new_n267_), .Y(new_new_n268_));
  AOI210     g246(.A0(new_new_n187_), .A1(new_new_n44_), .B0(new_new_n190_), .Y(new_new_n269_));
  NA2        g247(.A(i_0_), .B(new_new_n45_), .Y(new_new_n270_));
  NA3        g248(.A(new_new_n260_), .B(new_new_n166_), .C(new_new_n270_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n269_), .B(new_new_n271_), .Y(new_new_n272_));
  NO3        g250(.A(new_new_n272_), .B(new_new_n268_), .C(new_new_n265_), .Y(new_new_n273_));
  NOi21      g251(.An(i_10_), .B(i_6_), .Y(new_new_n274_));
  OR2        g252(.A(i_2_), .B(i_5_), .Y(new_new_n275_));
  OR2        g253(.A(new_new_n275_), .B(new_new_n212_), .Y(new_new_n276_));
  INV        g254(.A(new_new_n148_), .Y(new_new_n277_));
  AOI210     g255(.A0(new_new_n277_), .A1(new_new_n276_), .B0(new_new_n249_), .Y(new_new_n278_));
  INV        g256(.A(new_new_n278_), .Y(new_new_n279_));
  NA2        g257(.A(new_new_n279_), .B(new_new_n273_), .Y(new_new_n280_));
  NO3        g258(.A(new_new_n280_), .B(new_new_n259_), .C(new_new_n254_), .Y(new_new_n281_));
  NA4        g259(.A(new_new_n281_), .B(new_new_n224_), .C(new_new_n183_), .D(new_new_n161_), .Y(ori7));
  NO2        g260(.A(new_new_n80_), .B(new_new_n49_), .Y(new_new_n283_));
  NA2        g261(.A(new_new_n242_), .B(new_new_n72_), .Y(new_new_n284_));
  INV        g262(.A(i_11_), .Y(new_new_n285_));
  INV        g263(.A(new_new_n115_), .Y(new_new_n286_));
  NO2        g264(.A(new_new_n286_), .B(new_new_n284_), .Y(new_new_n287_));
  NA3        g265(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n288_));
  NA2        g266(.A(i_12_), .B(i_8_), .Y(new_new_n289_));
  NO2        g267(.A(new_new_n89_), .B(new_new_n288_), .Y(new_new_n290_));
  NA2        g268(.A(i_2_), .B(new_new_n73_), .Y(new_new_n291_));
  OAI210     g269(.A0(new_new_n74_), .A1(new_new_n129_), .B0(new_new_n130_), .Y(new_new_n292_));
  NA2        g270(.A(i_4_), .B(i_8_), .Y(new_new_n293_));
  INV        g271(.A(new_new_n168_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n294_), .B(new_new_n291_), .Y(new_new_n295_));
  NO4        g273(.A(new_new_n295_), .B(new_new_n290_), .C(new_new_n287_), .D(new_new_n283_), .Y(new_new_n296_));
  AOI210     g274(.A0(new_new_n106_), .A1(new_new_n54_), .B0(i_10_), .Y(new_new_n297_));
  AOI210     g275(.A0(new_new_n297_), .A1(new_new_n143_), .B0(new_new_n120_), .Y(new_new_n298_));
  OR2        g276(.A(i_6_), .B(i_10_), .Y(new_new_n299_));
  OR3        g277(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n300_));
  OR2        g278(.A(new_new_n298_), .B(new_new_n163_), .Y(new_new_n301_));
  AOI210     g279(.A0(new_new_n301_), .A1(new_new_n296_), .B0(new_new_n55_), .Y(new_new_n302_));
  NOi21      g280(.An(i_11_), .B(i_7_), .Y(new_new_n303_));
  AO210      g281(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n304_), .B(new_new_n303_), .Y(new_new_n305_));
  NA2        g283(.A(new_new_n305_), .B(new_new_n132_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n306_), .B(new_new_n55_), .Y(new_new_n307_));
  OR2        g285(.A(new_new_n133_), .B(new_new_n91_), .Y(new_new_n308_));
  NO2        g286(.A(i_1_), .B(i_12_), .Y(new_new_n309_));
  NA3        g287(.A(new_new_n309_), .B(new_new_n92_), .C(new_new_n24_), .Y(new_new_n310_));
  BUFFER     g288(.A(new_new_n310_), .Y(new_new_n311_));
  NA2        g289(.A(new_new_n311_), .B(new_new_n308_), .Y(new_new_n312_));
  OAI210     g290(.A0(new_new_n312_), .A1(new_new_n307_), .B0(i_6_), .Y(new_new_n313_));
  NO3        g291(.A(new_new_n299_), .B(new_new_n142_), .C(new_new_n23_), .Y(new_new_n314_));
  AOI210     g292(.A0(i_1_), .A1(new_new_n158_), .B0(new_new_n314_), .Y(new_new_n315_));
  NO2        g293(.A(new_new_n315_), .B(new_new_n42_), .Y(new_new_n316_));
  NO2        g294(.A(new_new_n44_), .B(i_1_), .Y(new_new_n317_));
  NA3        g295(.A(new_new_n317_), .B(new_new_n162_), .C(new_new_n42_), .Y(new_new_n318_));
  NO2        g296(.A(new_new_n515_), .B(new_new_n316_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n143_), .B(new_new_n85_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n320_), .B(new_new_n303_), .Y(new_new_n321_));
  NA2        g299(.A(new_new_n321_), .B(i_1_), .Y(new_new_n322_));
  NO2        g300(.A(new_new_n322_), .B(new_new_n300_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n213_), .B(new_new_n73_), .Y(new_new_n324_));
  NA2        g302(.A(new_new_n323_), .B(new_new_n44_), .Y(new_new_n325_));
  NA2        g303(.A(i_3_), .B(new_new_n128_), .Y(new_new_n326_));
  NO2        g304(.A(new_new_n142_), .B(new_new_n42_), .Y(new_new_n327_));
  NO3        g305(.A(new_new_n327_), .B(i_2_), .C(new_new_n144_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n329_), .B(i_6_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n73_), .B(i_9_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n331_), .B(new_new_n55_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n332_), .B(new_new_n309_), .Y(new_new_n333_));
  NO4        g311(.A(new_new_n333_), .B(new_new_n330_), .C(new_new_n328_), .D(i_4_), .Y(new_new_n334_));
  NA2        g312(.A(i_1_), .B(i_3_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n230_), .B(new_new_n80_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n327_), .B(new_new_n336_), .Y(new_new_n337_));
  NO2        g315(.A(new_new_n337_), .B(new_new_n335_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n338_), .B(new_new_n334_), .Y(new_new_n339_));
  NA4        g317(.A(new_new_n339_), .B(new_new_n325_), .C(new_new_n319_), .D(new_new_n313_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n193_), .B(new_new_n192_), .Y(new_new_n341_));
  AOI210     g319(.A0(new_new_n162_), .A1(new_new_n84_), .B0(i_1_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n191_), .B(i_2_), .Y(new_new_n343_));
  NA2        g321(.A(new_new_n343_), .B(new_new_n342_), .Y(new_new_n344_));
  AOI210     g322(.A0(new_new_n344_), .A1(new_new_n341_), .B0(i_13_), .Y(new_new_n345_));
  OR2        g323(.A(i_11_), .B(i_7_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n241_), .B(new_new_n24_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n347_), .B(new_new_n324_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(i_13_), .Y(new_new_n349_));
  INV        g327(.A(new_new_n349_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n284_), .B(new_new_n42_), .Y(new_new_n351_));
  NA2        g329(.A(new_new_n105_), .B(i_13_), .Y(new_new_n352_));
  NO2        g330(.A(new_new_n352_), .B(new_new_n342_), .Y(new_new_n353_));
  INV        g331(.A(i_7_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n79_), .B(new_new_n86_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n355_), .B(new_new_n289_), .Y(new_new_n356_));
  NO3        g334(.A(new_new_n356_), .B(new_new_n353_), .C(new_new_n351_), .Y(new_new_n357_));
  OR2        g335(.A(i_11_), .B(i_6_), .Y(new_new_n358_));
  NA2        g336(.A(i_12_), .B(i_7_), .Y(new_new_n359_));
  NO2        g337(.A(new_new_n359_), .B(new_new_n358_), .Y(new_new_n360_));
  NAi21      g338(.An(i_11_), .B(i_12_), .Y(new_new_n361_));
  NOi41      g339(.An(new_new_n93_), .B(new_new_n361_), .C(i_13_), .D(new_new_n73_), .Y(new_new_n362_));
  NO2        g340(.A(i_6_), .B(new_new_n293_), .Y(new_new_n363_));
  AOI210     g341(.A0(new_new_n363_), .A1(new_new_n170_), .B0(new_new_n362_), .Y(new_new_n364_));
  INV        g342(.A(new_new_n364_), .Y(new_new_n365_));
  OAI210     g343(.A0(new_new_n365_), .A1(new_new_n360_), .B0(new_new_n55_), .Y(new_new_n366_));
  NO2        g344(.A(i_2_), .B(i_12_), .Y(new_new_n367_));
  NA2        g345(.A(new_new_n190_), .B(new_new_n367_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n192_), .B(new_new_n190_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n369_), .B(new_new_n368_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n370_), .B(new_new_n43_), .Y(new_new_n371_));
  NA4        g349(.A(new_new_n371_), .B(new_new_n366_), .C(new_new_n357_), .D(new_new_n350_), .Y(new_new_n372_));
  OR4        g350(.A(new_new_n372_), .B(new_new_n345_), .C(new_new_n340_), .D(new_new_n302_), .Y(ori5));
  NA2        g351(.A(new_new_n321_), .B(new_new_n164_), .Y(new_new_n374_));
  AN2        g352(.A(new_new_n24_), .B(i_10_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n375_), .B(new_new_n367_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n289_), .B(i_11_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n74_), .B(new_new_n377_), .Y(new_new_n378_));
  NA3        g356(.A(new_new_n378_), .B(new_new_n376_), .C(new_new_n374_), .Y(new_new_n379_));
  NO3        g357(.A(i_11_), .B(new_new_n143_), .C(i_13_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n102_), .B(new_new_n23_), .Y(new_new_n381_));
  NA2        g359(.A(i_12_), .B(new_new_n381_), .Y(new_new_n382_));
  INV        g360(.A(new_new_n382_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n383_), .B(new_new_n379_), .Y(new_new_n384_));
  INV        g362(.A(new_new_n123_), .Y(new_new_n385_));
  INV        g363(.A(new_new_n149_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n343_), .B(new_new_n228_), .Y(new_new_n387_));
  AOI210     g365(.A0(new_new_n387_), .A1(new_new_n386_), .B0(new_new_n385_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n230_), .B(new_new_n26_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n389_), .B(new_new_n216_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n124_), .B(new_new_n128_), .Y(new_new_n391_));
  OA210      g369(.A0(new_new_n305_), .A1(new_new_n104_), .B0(i_13_), .Y(new_new_n392_));
  NO2        g370(.A(new_new_n133_), .B(new_new_n514_), .Y(new_new_n393_));
  NA2        g371(.A(new_new_n393_), .B(new_new_n216_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n85_), .B(new_new_n168_), .Y(new_new_n395_));
  OAI210     g373(.A0(new_new_n395_), .A1(i_11_), .B0(new_new_n394_), .Y(new_new_n396_));
  NO3        g374(.A(new_new_n396_), .B(new_new_n392_), .C(new_new_n391_), .Y(new_new_n397_));
  NO2        g375(.A(new_new_n54_), .B(i_12_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n104_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n399_), .B(new_new_n285_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n400_), .B(new_new_n36_), .Y(new_new_n401_));
  NA4        g379(.A(new_new_n401_), .B(new_new_n397_), .C(new_new_n516_), .D(new_new_n384_), .Y(ori6));
  NO2        g380(.A(new_new_n137_), .B(new_new_n244_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n151_), .B(i_9_), .Y(new_new_n404_));
  NA2        g382(.A(new_new_n404_), .B(new_new_n398_), .Y(new_new_n405_));
  AOI210     g383(.A0(new_new_n405_), .A1(new_new_n256_), .B0(new_new_n125_), .Y(new_new_n406_));
  NAi32      g384(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n358_), .B(new_new_n407_), .Y(new_new_n408_));
  OR2        g386(.A(new_new_n408_), .B(new_new_n406_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n346_), .B(i_2_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n45_), .B(new_new_n37_), .Y(new_new_n411_));
  INV        g389(.A(new_new_n411_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n412_), .B(new_new_n410_), .Y(new_new_n413_));
  BUFFER     g391(.A(new_new_n305_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n414_), .B(new_new_n117_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n415_), .B(new_new_n413_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n403_), .B(new_new_n354_), .Y(new_new_n417_));
  NA3        g395(.A(new_new_n195_), .B(new_new_n145_), .C(new_new_n117_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n207_), .B(new_new_n62_), .Y(new_new_n419_));
  NA4        g397(.A(new_new_n419_), .B(new_new_n418_), .C(new_new_n417_), .D(new_new_n292_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n228_), .B(new_new_n226_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n299_), .B(new_new_n86_), .Y(new_new_n422_));
  OAI210     g400(.A0(new_new_n422_), .A1(new_new_n94_), .B0(new_new_n211_), .Y(new_new_n423_));
  INV        g401(.A(new_new_n276_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n424_), .B(new_new_n172_), .Y(new_new_n425_));
  NA3        g403(.A(new_new_n425_), .B(new_new_n423_), .C(new_new_n421_), .Y(new_new_n426_));
  NO4        g404(.A(new_new_n426_), .B(new_new_n420_), .C(new_new_n416_), .D(new_new_n409_), .Y(new_new_n427_));
  NA2        g405(.A(new_new_n427_), .B(new_new_n203_), .Y(ori3));
  NA2        g406(.A(i_12_), .B(i_10_), .Y(new_new_n429_));
  NO2        g407(.A(i_11_), .B(new_new_n143_), .Y(new_new_n430_));
  NA3        g408(.A(new_new_n418_), .B(new_new_n292_), .C(new_new_n194_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n431_), .B(new_new_n40_), .Y(new_new_n432_));
  NOi21      g410(.An(new_new_n83_), .B(new_new_n390_), .Y(new_new_n433_));
  NO2        g411(.A(new_new_n308_), .B(new_new_n230_), .Y(new_new_n434_));
  AN2        g412(.A(new_new_n229_), .B(new_new_n50_), .Y(new_new_n435_));
  NO3        g413(.A(new_new_n435_), .B(new_new_n434_), .C(new_new_n433_), .Y(new_new_n436_));
  AOI210     g414(.A0(new_new_n436_), .A1(new_new_n432_), .B0(new_new_n45_), .Y(new_new_n437_));
  NO4        g415(.A(new_new_n199_), .B(new_new_n205_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n125_), .B(new_new_n274_), .Y(new_new_n439_));
  NOi21      g417(.An(new_new_n439_), .B(new_new_n438_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n440_), .B(new_new_n55_), .Y(new_new_n441_));
  NOi21      g419(.An(i_5_), .B(i_9_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n442_), .B(new_new_n225_), .Y(new_new_n443_));
  BUFFER     g421(.A(new_new_n162_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n444_), .B(new_new_n240_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n445_), .B(new_new_n443_), .Y(new_new_n446_));
  NO3        g424(.A(new_new_n446_), .B(new_new_n441_), .C(new_new_n437_), .Y(new_new_n447_));
  NO4        g425(.A(new_new_n275_), .B(i_12_), .C(new_new_n214_), .D(new_new_n212_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n448_), .B(i_11_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n380_), .B(new_new_n173_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n74_), .B(new_new_n52_), .Y(new_new_n451_));
  NO2        g429(.A(new_new_n451_), .B(new_new_n450_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n153_), .B(new_new_n118_), .Y(new_new_n453_));
  INV        g431(.A(new_new_n261_), .Y(new_new_n454_));
  NO4        g432(.A(new_new_n95_), .B(new_new_n52_), .C(new_new_n326_), .D(i_5_), .Y(new_new_n455_));
  AO220      g433(.A0(new_new_n455_), .A1(new_new_n454_), .B0(new_new_n453_), .B1(i_6_), .Y(new_new_n456_));
  NO2        g434(.A(new_new_n456_), .B(new_new_n452_), .Y(new_new_n457_));
  NA2        g435(.A(new_new_n457_), .B(new_new_n449_), .Y(new_new_n458_));
  NO2        g436(.A(new_new_n87_), .B(new_new_n37_), .Y(new_new_n459_));
  NA2        g437(.A(i_11_), .B(i_9_), .Y(new_new_n460_));
  NO3        g438(.A(i_12_), .B(new_new_n460_), .C(new_new_n291_), .Y(new_new_n461_));
  AN2        g439(.A(new_new_n461_), .B(new_new_n459_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n460_), .B(new_new_n65_), .Y(new_new_n463_));
  INV        g441(.A(new_new_n210_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n464_), .B(new_new_n443_), .Y(new_new_n465_));
  NO2        g443(.A(new_new_n465_), .B(new_new_n462_), .Y(new_new_n466_));
  INV        g444(.A(new_new_n466_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n429_), .B(new_new_n171_), .Y(new_new_n468_));
  OA210      g446(.A0(new_new_n239_), .A1(new_new_n139_), .B0(new_new_n238_), .Y(new_new_n469_));
  OAI210     g447(.A0(new_new_n469_), .A1(new_new_n468_), .B0(new_new_n463_), .Y(new_new_n470_));
  NA2        g448(.A(new_new_n347_), .B(new_new_n262_), .Y(new_new_n471_));
  NAi21      g449(.An(i_9_), .B(i_5_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n472_), .B(new_new_n209_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n473_), .B(new_new_n305_), .Y(new_new_n474_));
  OAI220     g452(.A0(new_new_n474_), .A1(new_new_n73_), .B0(new_new_n471_), .B1(new_new_n124_), .Y(new_new_n475_));
  NO2        g453(.A(new_new_n475_), .B(new_new_n259_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n476_), .B(new_new_n470_), .Y(new_new_n477_));
  NO3        g455(.A(new_new_n477_), .B(new_new_n467_), .C(new_new_n458_), .Y(new_new_n478_));
  NO3        g456(.A(new_new_n134_), .B(new_new_n205_), .C(i_0_), .Y(new_new_n479_));
  OAI210     g457(.A0(new_new_n479_), .A1(new_new_n67_), .B0(i_13_), .Y(new_new_n480_));
  INV        g458(.A(new_new_n480_), .Y(new_new_n481_));
  NO2        g459(.A(i_0_), .B(i_12_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n482_), .B(new_new_n469_), .Y(new_new_n483_));
  NA3        g461(.A(new_new_n206_), .B(new_new_n123_), .C(new_new_n122_), .Y(new_new_n484_));
  INV        g462(.A(new_new_n484_), .Y(new_new_n485_));
  NO3        g463(.A(new_new_n460_), .B(new_new_n136_), .C(new_new_n127_), .Y(new_new_n486_));
  NO2        g464(.A(new_new_n486_), .B(new_new_n485_), .Y(new_new_n487_));
  NA3        g465(.A(new_new_n487_), .B(new_new_n243_), .C(new_new_n483_), .Y(new_new_n488_));
  NO2        g466(.A(new_new_n73_), .B(i_5_), .Y(new_new_n489_));
  NA3        g467(.A(new_new_n430_), .B(new_new_n92_), .C(new_new_n102_), .Y(new_new_n490_));
  INV        g468(.A(new_new_n490_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n491_), .B(new_new_n489_), .Y(new_new_n492_));
  NAi21      g470(.An(i_10_), .B(new_new_n147_), .Y(new_new_n493_));
  NO4        g471(.A(new_new_n146_), .B(new_new_n134_), .C(i_0_), .D(i_12_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n494_), .B(new_new_n493_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n495_), .B(new_new_n492_), .Y(new_new_n496_));
  NO3        g474(.A(new_new_n496_), .B(new_new_n488_), .C(new_new_n481_), .Y(new_new_n497_));
  NA2        g475(.A(new_new_n410_), .B(new_new_n37_), .Y(new_new_n498_));
  NA2        g476(.A(new_new_n498_), .B(new_new_n298_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n499_), .B(new_new_n132_), .Y(new_new_n500_));
  NAi31      g478(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n501_));
  NO2        g479(.A(new_new_n62_), .B(new_new_n501_), .Y(new_new_n502_));
  AOI210     g480(.A0(new_new_n502_), .A1(new_new_n45_), .B0(new_new_n448_), .Y(new_new_n503_));
  AOI210     g481(.A0(new_new_n503_), .A1(new_new_n500_), .B0(new_new_n65_), .Y(new_new_n504_));
  INV        g482(.A(new_new_n202_), .Y(new_new_n505_));
  NO2        g483(.A(new_new_n505_), .B(new_new_n385_), .Y(new_new_n506_));
  NO3        g484(.A(new_new_n53_), .B(new_new_n52_), .C(i_4_), .Y(new_new_n507_));
  NA2        g485(.A(new_new_n169_), .B(new_new_n507_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n508_), .B(new_new_n361_), .Y(new_new_n509_));
  NO3        g487(.A(new_new_n509_), .B(new_new_n506_), .C(new_new_n504_), .Y(new_new_n510_));
  NA4        g488(.A(new_new_n510_), .B(new_new_n497_), .C(new_new_n478_), .D(new_new_n447_), .Y(ori4));
  INV        g489(.A(i_8_), .Y(new_new_n514_));
  INV        g490(.A(new_new_n318_), .Y(new_new_n515_));
  INV        g491(.A(new_new_n388_), .Y(new_new_n516_));
endmodule


