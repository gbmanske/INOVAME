library verilog;
use verilog.vl_types.all;
entity primeiro_vlg_vec_tst is
end primeiro_vlg_vec_tst;
