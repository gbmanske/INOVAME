// Benchmark "top" written by ABC on Fri Jun 21 17:49:26 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n138_, new_new_n139_,
    new_new_n140_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n657_, new_new_n658_,
    new_new_n659_, new_new_n660_, new_new_n661_, new_new_n662_,
    new_new_n663_, new_new_n664_, new_new_n665_, new_new_n666_,
    new_new_n667_, new_new_n668_, new_new_n669_, new_new_n670_,
    new_new_n671_, new_new_n672_, new_new_n673_, new_new_n674_,
    new_new_n675_, new_new_n676_, new_new_n677_, new_new_n678_,
    new_new_n679_, new_new_n680_, new_new_n681_, new_new_n682_,
    new_new_n683_, new_new_n684_, new_new_n685_, new_new_n686_,
    new_new_n687_, new_new_n688_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n706_, new_new_n707_,
    new_new_n708_, new_new_n709_, new_new_n710_, new_new_n711_,
    new_new_n712_, new_new_n713_, new_new_n714_, new_new_n715_,
    new_new_n716_, new_new_n717_, new_new_n718_, new_new_n719_,
    new_new_n720_, new_new_n721_, new_new_n722_, new_new_n723_,
    new_new_n724_, new_new_n725_, new_new_n726_, new_new_n727_,
    new_new_n728_, new_new_n729_, new_new_n730_, new_new_n731_,
    new_new_n732_, new_new_n733_, new_new_n734_, new_new_n735_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n924_, new_new_n925_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  NO2        g036(.A(new_new_n58_), .B(new_new_n57_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g039(.A(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NA3        g041(.A(new_new_n63_), .B(new_new_n61_), .C(new_new_n31_), .Y(new_new_n64_));
  NA2        g042(.A(i_1_), .B(i_10_), .Y(new_new_n65_));
  NO2        g043(.A(new_new_n65_), .B(i_6_), .Y(new_new_n66_));
  NAi31      g044(.An(new_new_n66_), .B(new_new_n64_), .C(new_new_n60_), .Y(new_new_n67_));
  NA2        g045(.A(new_new_n50_), .B(i_2_), .Y(new_new_n68_));
  AOI210     g046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n69_));
  NA2        g047(.A(i_1_), .B(i_6_), .Y(new_new_n70_));
  NO2        g048(.A(new_new_n70_), .B(new_new_n25_), .Y(new_new_n71_));
  INV        g049(.A(i_0_), .Y(new_new_n72_));
  NAi21      g050(.An(i_5_), .B(i_10_), .Y(new_new_n73_));
  NA2        g051(.A(i_5_), .B(i_9_), .Y(new_new_n74_));
  AOI210     g052(.A0(new_new_n74_), .A1(new_new_n73_), .B0(new_new_n72_), .Y(new_new_n75_));
  NO2        g053(.A(new_new_n75_), .B(new_new_n71_), .Y(new_new_n76_));
  OAI210     g054(.A0(new_new_n69_), .A1(new_new_n68_), .B0(new_new_n76_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n77_), .A1(new_new_n67_), .B0(i_0_), .Y(new_new_n78_));
  NA2        g056(.A(i_12_), .B(i_5_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_9_), .Y(new_new_n80_));
  NO2        g058(.A(i_3_), .B(i_7_), .Y(new_new_n81_));
  NO3        g059(.A(new_new_n81_), .B(new_new_n80_), .C(new_new_n62_), .Y(new_new_n82_));
  INV        g060(.A(i_6_), .Y(new_new_n83_));
  OR4        g061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n84_));
  INV        g062(.A(new_new_n84_), .Y(new_new_n85_));
  NO2        g063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  NO2        g064(.A(new_new_n85_), .B(new_new_n86_), .Y(new_new_n87_));
  NA2        g065(.A(new_new_n82_), .B(new_new_n87_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n62_), .Y(new_new_n91_));
  NA2        g069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  NO3        g070(.A(new_new_n92_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n93_));
  NO2        g071(.A(new_new_n93_), .B(new_new_n91_), .Y(new_new_n94_));
  AOI210     g072(.A0(new_new_n94_), .A1(new_new_n88_), .B0(new_new_n79_), .Y(new_new_n95_));
  AN3        g073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NO2        g075(.A(i_5_), .B(i_8_), .Y(new_new_n98_));
  NOi21      g076(.An(new_new_n98_), .B(new_new_n97_), .Y(new_new_n99_));
  AOI220     g077(.A0(new_new_n99_), .A1(new_new_n61_), .B0(new_new_n96_), .B1(new_new_n32_), .Y(new_new_n100_));
  INV        g078(.A(i_7_), .Y(new_new_n101_));
  NA2        g079(.A(new_new_n46_), .B(new_new_n101_), .Y(new_new_n102_));
  NO2        g080(.A(i_0_), .B(i_5_), .Y(new_new_n103_));
  NO2        g081(.A(new_new_n103_), .B(new_new_n83_), .Y(new_new_n104_));
  NA2        g082(.A(i_12_), .B(i_3_), .Y(new_new_n105_));
  INV        g083(.A(new_new_n105_), .Y(new_new_n106_));
  NA3        g084(.A(new_new_n106_), .B(new_new_n104_), .C(new_new_n102_), .Y(new_new_n107_));
  NAi21      g085(.An(i_7_), .B(i_11_), .Y(new_new_n108_));
  AN2        g086(.A(i_2_), .B(i_10_), .Y(new_new_n109_));
  NO2        g087(.A(new_new_n109_), .B(i_7_), .Y(new_new_n110_));
  OR2        g088(.A(new_new_n79_), .B(new_new_n57_), .Y(new_new_n111_));
  NO2        g089(.A(i_8_), .B(new_new_n101_), .Y(new_new_n112_));
  NO3        g090(.A(new_new_n112_), .B(new_new_n111_), .C(new_new_n110_), .Y(new_new_n113_));
  NA2        g091(.A(i_12_), .B(i_7_), .Y(new_new_n114_));
  NO2        g092(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n115_));
  NA2        g093(.A(new_new_n115_), .B(i_0_), .Y(new_new_n116_));
  NA2        g094(.A(i_11_), .B(i_12_), .Y(new_new_n117_));
  OAI210     g095(.A0(new_new_n116_), .A1(new_new_n114_), .B0(new_new_n117_), .Y(new_new_n118_));
  NO2        g096(.A(new_new_n118_), .B(new_new_n113_), .Y(new_new_n119_));
  NA3        g097(.A(new_new_n119_), .B(new_new_n107_), .C(new_new_n100_), .Y(new_new_n120_));
  NOi21      g098(.An(i_1_), .B(i_5_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n121_), .B(i_11_), .Y(new_new_n122_));
  NA2        g100(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n123_));
  NA2        g101(.A(i_7_), .B(new_new_n25_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(new_new_n123_), .Y(new_new_n125_));
  NO2        g103(.A(new_new_n125_), .B(new_new_n46_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n127_));
  NAi21      g105(.An(i_3_), .B(i_8_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(new_new_n61_), .Y(new_new_n129_));
  NOi31      g107(.An(new_new_n129_), .B(new_new_n127_), .C(new_new_n126_), .Y(new_new_n130_));
  NO2        g108(.A(i_1_), .B(new_new_n83_), .Y(new_new_n131_));
  NO2        g109(.A(i_6_), .B(i_5_), .Y(new_new_n132_));
  NA2        g110(.A(new_new_n132_), .B(i_3_), .Y(new_new_n133_));
  AO210      g111(.A0(new_new_n133_), .A1(new_new_n47_), .B0(new_new_n131_), .Y(new_new_n134_));
  OAI220     g112(.A0(new_new_n134_), .A1(new_new_n108_), .B0(new_new_n130_), .B1(new_new_n122_), .Y(new_new_n135_));
  NO3        g113(.A(new_new_n135_), .B(new_new_n120_), .C(new_new_n95_), .Y(new_new_n136_));
  NA3        g114(.A(new_new_n136_), .B(new_new_n78_), .C(new_new_n56_), .Y(ori2));
  NO2        g115(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n138_));
  INV        g116(.A(i_6_), .Y(new_new_n139_));
  NA2        g117(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n140_));
  NA4        g118(.A(new_new_n140_), .B(new_new_n76_), .C(new_new_n68_), .D(new_new_n30_), .Y(ori0));
  AN2        g119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  NA2        g120(.A(new_new_n142_), .B(i_6_), .Y(new_new_n143_));
  NO2        g121(.A(i_12_), .B(i_13_), .Y(new_new_n144_));
  NAi21      g122(.An(i_5_), .B(i_11_), .Y(new_new_n145_));
  NOi21      g123(.An(new_new_n144_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NA2        g125(.A(i_2_), .B(i_3_), .Y(new_new_n148_));
  NO2        g126(.A(new_new_n148_), .B(i_4_), .Y(new_new_n149_));
  NA3        g127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  AN2        g128(.A(new_new_n144_), .B(new_new_n80_), .Y(new_new_n151_));
  NA2        g129(.A(i_1_), .B(i_5_), .Y(new_new_n152_));
  NO2        g130(.A(new_new_n72_), .B(new_new_n46_), .Y(new_new_n153_));
  NA2        g131(.A(new_new_n153_), .B(new_new_n36_), .Y(new_new_n154_));
  OR2        g132(.A(i_0_), .B(i_1_), .Y(new_new_n155_));
  NO3        g133(.A(new_new_n155_), .B(new_new_n79_), .C(i_13_), .Y(new_new_n156_));
  NAi32      g134(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n157_));
  NAi21      g135(.An(new_new_n157_), .B(new_new_n156_), .Y(new_new_n158_));
  NOi21      g136(.An(i_4_), .B(i_10_), .Y(new_new_n159_));
  NA2        g137(.A(new_new_n159_), .B(new_new_n40_), .Y(new_new_n160_));
  NO2        g138(.A(i_3_), .B(i_5_), .Y(new_new_n161_));
  NO3        g139(.A(new_new_n72_), .B(i_2_), .C(i_1_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  OAI210     g141(.A0(new_new_n163_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n164_));
  INV        g142(.A(new_new_n164_), .Y(new_new_n165_));
  NO2        g143(.A(new_new_n165_), .B(new_new_n143_), .Y(new_new_n166_));
  NOi21      g144(.An(i_4_), .B(i_9_), .Y(new_new_n167_));
  NOi21      g145(.An(i_11_), .B(i_13_), .Y(new_new_n168_));
  NA2        g146(.A(new_new_n168_), .B(new_new_n167_), .Y(new_new_n169_));
  NO2        g147(.A(i_4_), .B(i_5_), .Y(new_new_n170_));
  NAi21      g148(.An(i_12_), .B(i_11_), .Y(new_new_n171_));
  NO2        g149(.A(new_new_n171_), .B(i_13_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n72_), .B(new_new_n62_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(new_new_n46_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n36_), .B(i_5_), .Y(new_new_n175_));
  NAi31      g153(.An(new_new_n175_), .B(new_new_n151_), .C(i_11_), .Y(new_new_n176_));
  NA2        g154(.A(i_3_), .B(i_5_), .Y(new_new_n177_));
  OR2        g155(.A(new_new_n177_), .B(new_new_n169_), .Y(new_new_n178_));
  AOI210     g156(.A0(new_new_n178_), .A1(new_new_n176_), .B0(new_new_n174_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n72_), .B(i_5_), .Y(new_new_n180_));
  NO2        g158(.A(i_13_), .B(i_10_), .Y(new_new_n181_));
  NA3        g159(.A(new_new_n181_), .B(new_new_n180_), .C(new_new_n44_), .Y(new_new_n182_));
  NO2        g160(.A(i_2_), .B(i_1_), .Y(new_new_n183_));
  NAi21      g161(.An(i_4_), .B(i_12_), .Y(new_new_n184_));
  INV        g162(.A(new_new_n179_), .Y(new_new_n185_));
  INV        g163(.A(i_8_), .Y(new_new_n186_));
  NO2        g164(.A(new_new_n186_), .B(i_7_), .Y(new_new_n187_));
  NA2        g165(.A(new_new_n187_), .B(i_6_), .Y(new_new_n188_));
  NO3        g166(.A(i_3_), .B(new_new_n83_), .C(new_new_n48_), .Y(new_new_n189_));
  NO3        g167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n190_));
  NO3        g168(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n191_));
  NO2        g169(.A(i_3_), .B(i_8_), .Y(new_new_n192_));
  NO3        g170(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n193_));
  NA3        g171(.A(new_new_n193_), .B(new_new_n192_), .C(new_new_n40_), .Y(new_new_n194_));
  NO2        g172(.A(new_new_n103_), .B(new_new_n57_), .Y(new_new_n195_));
  INV        g173(.A(new_new_n195_), .Y(new_new_n196_));
  NO2        g174(.A(i_13_), .B(i_9_), .Y(new_new_n197_));
  NAi21      g175(.An(i_12_), .B(i_3_), .Y(new_new_n198_));
  NO2        g176(.A(new_new_n44_), .B(i_5_), .Y(new_new_n199_));
  NO3        g177(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n196_), .B(new_new_n194_), .Y(new_new_n201_));
  NA2        g179(.A(new_new_n201_), .B(i_7_), .Y(new_new_n202_));
  OAI220     g180(.A0(new_new_n202_), .A1(i_4_), .B0(new_new_n188_), .B1(new_new_n185_), .Y(new_new_n203_));
  NAi21      g181(.An(i_12_), .B(i_7_), .Y(new_new_n204_));
  NA3        g182(.A(i_13_), .B(new_new_n186_), .C(i_10_), .Y(new_new_n205_));
  NA2        g183(.A(i_0_), .B(i_5_), .Y(new_new_n206_));
  NAi31      g184(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n207_));
  NO2        g185(.A(new_new_n36_), .B(i_13_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n72_), .B(new_new_n26_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n46_), .B(new_new_n62_), .Y(new_new_n210_));
  NA3        g188(.A(new_new_n210_), .B(new_new_n209_), .C(new_new_n208_), .Y(new_new_n211_));
  INV        g189(.A(i_13_), .Y(new_new_n212_));
  NO2        g190(.A(i_12_), .B(new_new_n212_), .Y(new_new_n213_));
  NA3        g191(.A(new_new_n213_), .B(new_new_n190_), .C(new_new_n189_), .Y(new_new_n214_));
  OAI210     g192(.A0(new_new_n211_), .A1(new_new_n207_), .B0(new_new_n214_), .Y(new_new_n215_));
  NA2        g193(.A(new_new_n215_), .B(new_new_n142_), .Y(new_new_n216_));
  NO2        g194(.A(i_12_), .B(new_new_n37_), .Y(new_new_n217_));
  OR2        g195(.A(i_8_), .B(i_7_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n53_), .B(i_1_), .Y(new_new_n219_));
  INV        g197(.A(i_12_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n44_), .B(new_new_n220_), .Y(new_new_n221_));
  NO3        g199(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n222_));
  NA2        g200(.A(i_2_), .B(i_1_), .Y(new_new_n223_));
  NO3        g201(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n224_));
  NAi21      g202(.An(i_4_), .B(i_3_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n225_), .B(new_new_n74_), .Y(new_new_n226_));
  NO2        g204(.A(i_0_), .B(i_6_), .Y(new_new_n227_));
  NOi41      g205(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n223_), .B(new_new_n177_), .Y(new_new_n229_));
  NO2        g207(.A(i_11_), .B(new_new_n212_), .Y(new_new_n230_));
  NOi21      g208(.An(i_1_), .B(i_6_), .Y(new_new_n231_));
  NAi21      g209(.An(i_3_), .B(i_7_), .Y(new_new_n232_));
  NA2        g210(.A(new_new_n220_), .B(i_9_), .Y(new_new_n233_));
  NA2        g211(.A(new_new_n72_), .B(i_5_), .Y(new_new_n234_));
  NAi21      g212(.An(i_7_), .B(i_10_), .Y(new_new_n235_));
  INV        g213(.A(new_new_n143_), .Y(new_new_n236_));
  NA2        g214(.A(new_new_n220_), .B(i_13_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n237_), .B(new_new_n74_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n238_), .B(new_new_n236_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n218_), .B(new_new_n37_), .Y(new_new_n240_));
  NA2        g218(.A(i_12_), .B(i_6_), .Y(new_new_n241_));
  OR2        g219(.A(i_13_), .B(i_9_), .Y(new_new_n242_));
  NO3        g220(.A(new_new_n242_), .B(new_new_n241_), .C(new_new_n48_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n225_), .B(i_2_), .Y(new_new_n244_));
  NA3        g222(.A(new_new_n244_), .B(new_new_n243_), .C(new_new_n44_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n230_), .B(i_9_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n234_), .B(new_new_n63_), .Y(new_new_n247_));
  OAI210     g225(.A0(new_new_n247_), .A1(new_new_n246_), .B0(new_new_n245_), .Y(new_new_n248_));
  NA2        g226(.A(new_new_n153_), .B(new_new_n62_), .Y(new_new_n249_));
  NO3        g227(.A(i_11_), .B(new_new_n212_), .C(new_new_n25_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n232_), .B(i_8_), .Y(new_new_n251_));
  NO2        g229(.A(i_6_), .B(new_new_n48_), .Y(new_new_n252_));
  NA3        g230(.A(new_new_n252_), .B(new_new_n251_), .C(new_new_n250_), .Y(new_new_n253_));
  NO3        g231(.A(new_new_n26_), .B(new_new_n83_), .C(i_5_), .Y(new_new_n254_));
  NA3        g232(.A(new_new_n254_), .B(new_new_n240_), .C(new_new_n213_), .Y(new_new_n255_));
  AOI210     g233(.A0(new_new_n255_), .A1(new_new_n253_), .B0(new_new_n249_), .Y(new_new_n256_));
  AOI210     g234(.A0(new_new_n248_), .A1(new_new_n240_), .B0(new_new_n256_), .Y(new_new_n257_));
  NA3        g235(.A(new_new_n257_), .B(new_new_n239_), .C(new_new_n216_), .Y(new_new_n258_));
  NO3        g236(.A(i_12_), .B(new_new_n212_), .C(new_new_n37_), .Y(new_new_n259_));
  INV        g237(.A(new_new_n259_), .Y(new_new_n260_));
  NA2        g238(.A(i_8_), .B(new_new_n101_), .Y(new_new_n261_));
  NO3        g239(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n262_));
  AOI220     g240(.A0(new_new_n262_), .A1(new_new_n189_), .B0(new_new_n161_), .B1(new_new_n219_), .Y(new_new_n263_));
  NO2        g241(.A(new_new_n263_), .B(new_new_n261_), .Y(new_new_n264_));
  NO3        g242(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n265_));
  NO2        g243(.A(new_new_n223_), .B(i_0_), .Y(new_new_n266_));
  AOI220     g244(.A0(new_new_n266_), .A1(new_new_n187_), .B0(new_new_n265_), .B1(new_new_n142_), .Y(new_new_n267_));
  NA2        g245(.A(new_new_n252_), .B(new_new_n26_), .Y(new_new_n268_));
  NO2        g246(.A(new_new_n268_), .B(new_new_n267_), .Y(new_new_n269_));
  NA2        g247(.A(i_0_), .B(i_1_), .Y(new_new_n270_));
  NO2        g248(.A(new_new_n270_), .B(i_2_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n58_), .B(i_6_), .Y(new_new_n272_));
  NO2        g250(.A(new_new_n163_), .B(new_new_n143_), .Y(new_new_n273_));
  NO3        g251(.A(new_new_n273_), .B(new_new_n269_), .C(new_new_n264_), .Y(new_new_n274_));
  NO2        g252(.A(i_3_), .B(i_10_), .Y(new_new_n275_));
  NO2        g253(.A(i_2_), .B(new_new_n101_), .Y(new_new_n276_));
  NA2        g254(.A(i_1_), .B(new_new_n36_), .Y(new_new_n277_));
  AN2        g255(.A(i_3_), .B(i_10_), .Y(new_new_n278_));
  NO2        g256(.A(i_5_), .B(new_new_n37_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n274_), .B(new_new_n260_), .Y(new_new_n281_));
  NO4        g259(.A(new_new_n281_), .B(new_new_n258_), .C(new_new_n203_), .D(new_new_n166_), .Y(new_new_n282_));
  NO3        g260(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n58_), .B(new_new_n83_), .Y(new_new_n284_));
  NA2        g262(.A(new_new_n266_), .B(new_new_n284_), .Y(new_new_n285_));
  NO3        g263(.A(i_6_), .B(new_new_n186_), .C(i_7_), .Y(new_new_n286_));
  NA2        g264(.A(new_new_n286_), .B(new_new_n190_), .Y(new_new_n287_));
  AOI210     g265(.A0(new_new_n287_), .A1(new_new_n285_), .B0(i_5_), .Y(new_new_n288_));
  NO2        g266(.A(i_2_), .B(i_3_), .Y(new_new_n289_));
  OR2        g267(.A(i_0_), .B(i_5_), .Y(new_new_n290_));
  NA3        g268(.A(new_new_n266_), .B(new_new_n161_), .C(new_new_n112_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n155_), .B(new_new_n46_), .Y(new_new_n292_));
  INV        g270(.A(new_new_n291_), .Y(new_new_n293_));
  OAI210     g271(.A0(new_new_n293_), .A1(new_new_n288_), .B0(i_4_), .Y(new_new_n294_));
  NO2        g272(.A(i_12_), .B(i_10_), .Y(new_new_n295_));
  NOi21      g273(.An(i_5_), .B(i_0_), .Y(new_new_n296_));
  NO2        g274(.A(i_2_), .B(new_new_n101_), .Y(new_new_n297_));
  NO4        g275(.A(new_new_n297_), .B(new_new_n277_), .C(new_new_n296_), .D(new_new_n128_), .Y(new_new_n298_));
  NA4        g276(.A(new_new_n81_), .B(new_new_n36_), .C(new_new_n83_), .D(i_8_), .Y(new_new_n299_));
  NA2        g277(.A(new_new_n298_), .B(new_new_n295_), .Y(new_new_n300_));
  NO2        g278(.A(i_6_), .B(i_8_), .Y(new_new_n301_));
  NOi21      g279(.An(i_0_), .B(i_2_), .Y(new_new_n302_));
  AN2        g280(.A(new_new_n302_), .B(new_new_n301_), .Y(new_new_n303_));
  NO2        g281(.A(i_1_), .B(i_7_), .Y(new_new_n304_));
  NA2        g282(.A(new_new_n300_), .B(new_new_n294_), .Y(new_new_n305_));
  NOi21      g283(.An(new_new_n152_), .B(new_new_n104_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n306_), .B(new_new_n124_), .Y(new_new_n307_));
  NA2        g285(.A(new_new_n307_), .B(i_3_), .Y(new_new_n308_));
  INV        g286(.A(new_new_n92_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n186_), .B(i_9_), .Y(new_new_n310_));
  NA2        g288(.A(new_new_n310_), .B(new_new_n195_), .Y(new_new_n311_));
  NO2        g289(.A(new_new_n311_), .B(new_new_n46_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n312_), .B(new_new_n269_), .Y(new_new_n313_));
  AOI210     g291(.A0(new_new_n313_), .A1(new_new_n308_), .B0(new_new_n160_), .Y(new_new_n314_));
  AOI210     g292(.A0(new_new_n305_), .A1(new_new_n283_), .B0(new_new_n314_), .Y(new_new_n315_));
  NOi32      g293(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n316_));
  INV        g294(.A(new_new_n316_), .Y(new_new_n317_));
  NO2        g295(.A(new_new_n207_), .B(new_new_n157_), .Y(new_new_n318_));
  NO2        g296(.A(new_new_n157_), .B(new_new_n155_), .Y(new_new_n319_));
  NOi32      g297(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n320_));
  NAi21      g298(.An(i_6_), .B(i_1_), .Y(new_new_n321_));
  NA3        g299(.A(new_new_n321_), .B(new_new_n320_), .C(new_new_n46_), .Y(new_new_n322_));
  NO2        g300(.A(new_new_n322_), .B(i_0_), .Y(new_new_n323_));
  OR3        g301(.A(new_new_n323_), .B(new_new_n319_), .C(new_new_n318_), .Y(new_new_n324_));
  NO2        g302(.A(i_1_), .B(new_new_n101_), .Y(new_new_n325_));
  NAi21      g303(.An(i_3_), .B(i_4_), .Y(new_new_n326_));
  NO2        g304(.A(new_new_n326_), .B(i_9_), .Y(new_new_n327_));
  AN2        g305(.A(i_6_), .B(i_7_), .Y(new_new_n328_));
  OAI210     g306(.A0(new_new_n328_), .A1(new_new_n325_), .B0(new_new_n327_), .Y(new_new_n329_));
  NA2        g307(.A(i_2_), .B(i_7_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n326_), .B(i_10_), .Y(new_new_n331_));
  NA3        g309(.A(new_new_n331_), .B(new_new_n330_), .C(new_new_n227_), .Y(new_new_n332_));
  AOI210     g310(.A0(new_new_n332_), .A1(new_new_n329_), .B0(new_new_n180_), .Y(new_new_n333_));
  AOI210     g311(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n334_));
  OAI210     g312(.A0(new_new_n334_), .A1(new_new_n183_), .B0(new_new_n331_), .Y(new_new_n335_));
  AOI220     g313(.A0(new_new_n331_), .A1(new_new_n304_), .B0(new_new_n222_), .B1(new_new_n183_), .Y(new_new_n336_));
  AOI210     g314(.A0(new_new_n336_), .A1(new_new_n335_), .B0(i_5_), .Y(new_new_n337_));
  NO3        g315(.A(new_new_n337_), .B(new_new_n333_), .C(new_new_n324_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n338_), .B(new_new_n317_), .Y(new_new_n339_));
  NO2        g317(.A(new_new_n58_), .B(new_new_n25_), .Y(new_new_n340_));
  AN2        g318(.A(i_12_), .B(i_5_), .Y(new_new_n341_));
  NO2        g319(.A(i_4_), .B(new_new_n26_), .Y(new_new_n342_));
  NA2        g320(.A(new_new_n342_), .B(new_new_n341_), .Y(new_new_n343_));
  NO2        g321(.A(i_11_), .B(i_6_), .Y(new_new_n344_));
  NA3        g322(.A(new_new_n344_), .B(new_new_n292_), .C(new_new_n212_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n345_), .B(new_new_n343_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n225_), .B(i_5_), .Y(new_new_n347_));
  NO2        g325(.A(i_5_), .B(i_10_), .Y(new_new_n348_));
  AOI220     g326(.A0(new_new_n348_), .A1(new_new_n244_), .B0(new_new_n347_), .B1(new_new_n190_), .Y(new_new_n349_));
  NA2        g327(.A(new_new_n144_), .B(new_new_n45_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n350_), .B(new_new_n349_), .Y(new_new_n351_));
  OAI210     g329(.A0(new_new_n351_), .A1(new_new_n346_), .B0(new_new_n340_), .Y(new_new_n352_));
  NO2        g330(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n150_), .B(new_new_n83_), .Y(new_new_n354_));
  OAI210     g332(.A0(new_new_n354_), .A1(new_new_n346_), .B0(new_new_n353_), .Y(new_new_n355_));
  NO3        g333(.A(new_new_n83_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n356_));
  NA3        g334(.A(new_new_n275_), .B(new_new_n74_), .C(new_new_n54_), .Y(new_new_n357_));
  NO2        g335(.A(i_11_), .B(i_12_), .Y(new_new_n358_));
  NA2        g336(.A(new_new_n358_), .B(new_new_n36_), .Y(new_new_n359_));
  NO2        g337(.A(new_new_n357_), .B(new_new_n359_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n348_), .B(new_new_n220_), .Y(new_new_n361_));
  NAi21      g339(.An(i_13_), .B(i_0_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n362_), .B(new_new_n223_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n360_), .B(new_new_n363_), .Y(new_new_n364_));
  NA3        g342(.A(new_new_n364_), .B(new_new_n355_), .C(new_new_n352_), .Y(new_new_n365_));
  NA2        g343(.A(new_new_n44_), .B(new_new_n212_), .Y(new_new_n366_));
  NO2        g344(.A(i_0_), .B(i_11_), .Y(new_new_n367_));
  AN2        g345(.A(i_1_), .B(i_6_), .Y(new_new_n368_));
  NOi21      g346(.An(i_2_), .B(i_12_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n142_), .B(i_9_), .Y(new_new_n370_));
  NO2        g348(.A(new_new_n370_), .B(i_4_), .Y(new_new_n371_));
  NAi21      g349(.An(i_9_), .B(i_4_), .Y(new_new_n372_));
  OR2        g350(.A(i_13_), .B(i_10_), .Y(new_new_n373_));
  NO3        g351(.A(new_new_n373_), .B(new_new_n117_), .C(new_new_n372_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n169_), .B(new_new_n123_), .Y(new_new_n375_));
  NO2        g353(.A(new_new_n101_), .B(new_new_n25_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n259_), .B(new_new_n376_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n377_), .B(new_new_n306_), .Y(new_new_n378_));
  INV        g356(.A(new_new_n378_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(new_new_n26_), .Y(new_new_n380_));
  INV        g358(.A(new_new_n291_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n177_), .B(new_new_n83_), .Y(new_new_n382_));
  AOI220     g360(.A0(new_new_n382_), .A1(new_new_n271_), .B0(new_new_n254_), .B1(new_new_n200_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n383_), .B(new_new_n261_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n384_), .B(new_new_n381_), .Y(new_new_n385_));
  NA2        g363(.A(new_new_n189_), .B(new_new_n96_), .Y(new_new_n386_));
  NA3        g364(.A(new_new_n292_), .B(new_new_n161_), .C(new_new_n83_), .Y(new_new_n387_));
  AOI210     g365(.A0(new_new_n387_), .A1(new_new_n386_), .B0(i_8_), .Y(new_new_n388_));
  NA3        g366(.A(new_new_n234_), .B(new_new_n63_), .C(i_2_), .Y(new_new_n389_));
  NA2        g367(.A(new_new_n272_), .B(new_new_n219_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n390_), .B(new_new_n177_), .Y(new_new_n391_));
  NO2        g369(.A(i_3_), .B(new_new_n48_), .Y(new_new_n392_));
  NA3        g370(.A(new_new_n304_), .B(new_new_n303_), .C(new_new_n392_), .Y(new_new_n393_));
  INV        g371(.A(new_new_n393_), .Y(new_new_n394_));
  NO3        g372(.A(new_new_n394_), .B(new_new_n391_), .C(new_new_n388_), .Y(new_new_n395_));
  AOI210     g373(.A0(new_new_n395_), .A1(new_new_n385_), .B0(new_new_n246_), .Y(new_new_n396_));
  NO4        g374(.A(new_new_n396_), .B(new_new_n380_), .C(new_new_n365_), .D(new_new_n339_), .Y(new_new_n397_));
  NO2        g375(.A(new_new_n72_), .B(i_13_), .Y(new_new_n398_));
  NO2        g376(.A(i_10_), .B(i_9_), .Y(new_new_n399_));
  NAi21      g377(.An(i_12_), .B(i_8_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n400_), .B(i_3_), .Y(new_new_n401_));
  NO2        g379(.A(new_new_n46_), .B(i_4_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n402_), .B(new_new_n104_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n403_), .B(new_new_n194_), .Y(new_new_n404_));
  NA2        g382(.A(new_new_n280_), .B(i_0_), .Y(new_new_n405_));
  NO3        g383(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n241_), .B(new_new_n97_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n407_), .B(new_new_n406_), .Y(new_new_n408_));
  NA2        g386(.A(i_8_), .B(i_9_), .Y(new_new_n409_));
  AOI210     g387(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n410_));
  OR2        g388(.A(new_new_n410_), .B(new_new_n409_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n259_), .B(new_new_n195_), .Y(new_new_n412_));
  OAI220     g390(.A0(new_new_n412_), .A1(new_new_n411_), .B0(new_new_n408_), .B1(new_new_n405_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n230_), .B(new_new_n279_), .Y(new_new_n414_));
  NO3        g392(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n415_));
  INV        g393(.A(new_new_n415_), .Y(new_new_n416_));
  NA3        g394(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n417_));
  NA4        g395(.A(new_new_n145_), .B(new_new_n115_), .C(new_new_n79_), .D(new_new_n23_), .Y(new_new_n418_));
  OAI220     g396(.A0(new_new_n418_), .A1(new_new_n417_), .B0(new_new_n416_), .B1(new_new_n414_), .Y(new_new_n419_));
  NO3        g397(.A(new_new_n419_), .B(new_new_n413_), .C(new_new_n404_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n96_), .B(i_13_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n382_), .B(new_new_n340_), .Y(new_new_n422_));
  NO2        g400(.A(i_2_), .B(i_13_), .Y(new_new_n423_));
  NO2        g401(.A(new_new_n422_), .B(new_new_n421_), .Y(new_new_n424_));
  NO3        g402(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n425_));
  NO2        g403(.A(i_6_), .B(i_7_), .Y(new_new_n426_));
  NO2        g404(.A(i_11_), .B(i_1_), .Y(new_new_n427_));
  NOi21      g405(.An(i_2_), .B(i_7_), .Y(new_new_n428_));
  NO2        g406(.A(i_3_), .B(new_new_n186_), .Y(new_new_n429_));
  NO2        g407(.A(i_6_), .B(i_10_), .Y(new_new_n430_));
  NA3        g408(.A(new_new_n228_), .B(new_new_n168_), .C(new_new_n132_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n155_), .B(i_3_), .Y(new_new_n433_));
  NAi31      g411(.An(new_new_n432_), .B(new_new_n433_), .C(new_new_n213_), .Y(new_new_n434_));
  NA3        g412(.A(new_new_n353_), .B(new_new_n173_), .C(new_new_n149_), .Y(new_new_n435_));
  NA3        g413(.A(new_new_n435_), .B(new_new_n434_), .C(new_new_n431_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n436_), .B(new_new_n424_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n406_), .B(new_new_n341_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n415_), .B(new_new_n348_), .Y(new_new_n439_));
  NO2        g417(.A(new_new_n439_), .B(new_new_n211_), .Y(new_new_n440_));
  NAi21      g418(.An(new_new_n205_), .B(new_new_n358_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n304_), .B(new_new_n206_), .Y(new_new_n442_));
  NO2        g420(.A(new_new_n442_), .B(new_new_n441_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n27_), .B(i_10_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n283_), .B(new_new_n222_), .Y(new_new_n445_));
  OAI220     g423(.A0(new_new_n445_), .A1(new_new_n389_), .B0(new_new_n444_), .B1(new_new_n421_), .Y(new_new_n446_));
  NO3        g424(.A(new_new_n446_), .B(new_new_n443_), .C(new_new_n440_), .Y(new_new_n447_));
  NA3        g425(.A(new_new_n447_), .B(new_new_n437_), .C(new_new_n420_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n122_), .B(new_new_n111_), .Y(new_new_n449_));
  AN2        g427(.A(new_new_n449_), .B(new_new_n406_), .Y(new_new_n450_));
  NA2        g428(.A(new_new_n450_), .B(new_new_n280_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n341_), .B(new_new_n212_), .Y(new_new_n452_));
  NA2        g430(.A(new_new_n316_), .B(new_new_n72_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n328_), .B(new_new_n320_), .Y(new_new_n454_));
  OR2        g432(.A(new_new_n452_), .B(new_new_n454_), .Y(new_new_n455_));
  NO2        g433(.A(new_new_n36_), .B(i_8_), .Y(new_new_n456_));
  AOI210     g434(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n374_), .Y(new_new_n457_));
  NA2        g435(.A(new_new_n457_), .B(new_new_n455_), .Y(new_new_n458_));
  INV        g436(.A(new_new_n458_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n234_), .B(new_new_n63_), .Y(new_new_n460_));
  OAI210     g438(.A0(i_8_), .A1(new_new_n460_), .B0(new_new_n134_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n461_), .B(new_new_n375_), .Y(new_new_n462_));
  NA3        g440(.A(new_new_n462_), .B(new_new_n459_), .C(new_new_n451_), .Y(new_new_n463_));
  NO2        g441(.A(i_12_), .B(new_new_n186_), .Y(new_new_n464_));
  NO2        g442(.A(i_8_), .B(i_7_), .Y(new_new_n465_));
  OAI210     g443(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n466_), .B(new_new_n210_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n467_), .B(new_new_n225_), .Y(new_new_n468_));
  NA2        g446(.A(new_new_n44_), .B(i_10_), .Y(new_new_n469_));
  NO2        g447(.A(new_new_n469_), .B(i_6_), .Y(new_new_n470_));
  NA3        g448(.A(new_new_n470_), .B(new_new_n468_), .C(new_new_n465_), .Y(new_new_n471_));
  AOI220     g449(.A0(new_new_n382_), .A1(new_new_n292_), .B0(new_new_n229_), .B1(new_new_n227_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n472_), .B(new_new_n237_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n473_), .B(new_new_n240_), .Y(new_new_n474_));
  NA3        g452(.A(new_new_n278_), .B(new_new_n170_), .C(new_new_n96_), .Y(new_new_n475_));
  NO2        g453(.A(new_new_n208_), .B(new_new_n44_), .Y(new_new_n476_));
  NO2        g454(.A(new_new_n155_), .B(i_5_), .Y(new_new_n477_));
  NA3        g455(.A(new_new_n477_), .B(new_new_n366_), .C(new_new_n289_), .Y(new_new_n478_));
  OAI210     g456(.A0(new_new_n478_), .A1(new_new_n476_), .B0(new_new_n475_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n479_), .B(new_new_n415_), .Y(new_new_n480_));
  NA3        g458(.A(new_new_n480_), .B(new_new_n474_), .C(new_new_n471_), .Y(new_new_n481_));
  AOI210     g459(.A0(new_new_n321_), .A1(new_new_n46_), .B0(new_new_n325_), .Y(new_new_n482_));
  NA2        g460(.A(i_0_), .B(new_new_n48_), .Y(new_new_n483_));
  NA3        g461(.A(new_new_n464_), .B(new_new_n250_), .C(new_new_n483_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n482_), .B(new_new_n484_), .Y(new_new_n485_));
  INV        g463(.A(new_new_n485_), .Y(new_new_n486_));
  NO3        g464(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n487_));
  NO2        g465(.A(new_new_n218_), .B(new_new_n36_), .Y(new_new_n488_));
  NO2        g466(.A(new_new_n373_), .B(i_1_), .Y(new_new_n489_));
  NOi31      g467(.An(new_new_n489_), .B(new_new_n407_), .C(new_new_n72_), .Y(new_new_n490_));
  AN4        g468(.A(new_new_n490_), .B(new_new_n371_), .C(i_3_), .D(i_2_), .Y(new_new_n491_));
  INV        g469(.A(new_new_n491_), .Y(new_new_n492_));
  NOi21      g470(.An(i_10_), .B(i_6_), .Y(new_new_n493_));
  NO2        g471(.A(new_new_n83_), .B(new_new_n25_), .Y(new_new_n494_));
  AOI220     g472(.A0(new_new_n259_), .A1(new_new_n494_), .B0(new_new_n250_), .B1(new_new_n493_), .Y(new_new_n495_));
  NO2        g473(.A(new_new_n495_), .B(new_new_n405_), .Y(new_new_n496_));
  NO2        g474(.A(new_new_n114_), .B(new_new_n23_), .Y(new_new_n497_));
  NA2        g475(.A(new_new_n286_), .B(new_new_n162_), .Y(new_new_n498_));
  AOI220     g476(.A0(new_new_n498_), .A1(new_new_n390_), .B0(new_new_n178_), .B1(new_new_n176_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n190_), .B(new_new_n37_), .Y(new_new_n500_));
  NOi31      g478(.An(new_new_n146_), .B(new_new_n500_), .C(new_new_n299_), .Y(new_new_n501_));
  NO3        g479(.A(new_new_n501_), .B(new_new_n499_), .C(new_new_n496_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n453_), .B(new_new_n336_), .Y(new_new_n503_));
  INV        g481(.A(new_new_n289_), .Y(new_new_n504_));
  NO2        g482(.A(i_12_), .B(new_new_n83_), .Y(new_new_n505_));
  NA3        g483(.A(new_new_n505_), .B(new_new_n250_), .C(new_new_n483_), .Y(new_new_n506_));
  NA3        g484(.A(new_new_n344_), .B(new_new_n259_), .C(new_new_n206_), .Y(new_new_n507_));
  AOI210     g485(.A0(new_new_n507_), .A1(new_new_n506_), .B0(new_new_n504_), .Y(new_new_n508_));
  OR2        g486(.A(i_2_), .B(i_5_), .Y(new_new_n509_));
  OR2        g487(.A(new_new_n509_), .B(new_new_n368_), .Y(new_new_n510_));
  NA2        g488(.A(new_new_n330_), .B(new_new_n227_), .Y(new_new_n511_));
  AOI210     g489(.A0(new_new_n511_), .A1(new_new_n510_), .B0(new_new_n441_), .Y(new_new_n512_));
  NO3        g490(.A(new_new_n512_), .B(new_new_n508_), .C(new_new_n503_), .Y(new_new_n513_));
  NA4        g491(.A(new_new_n513_), .B(new_new_n502_), .C(new_new_n492_), .D(new_new_n486_), .Y(new_new_n514_));
  NO4        g492(.A(new_new_n514_), .B(new_new_n481_), .C(new_new_n463_), .D(new_new_n448_), .Y(new_new_n515_));
  NA4        g493(.A(new_new_n515_), .B(new_new_n397_), .C(new_new_n315_), .D(new_new_n282_), .Y(ori7));
  NO2        g494(.A(new_new_n92_), .B(new_new_n54_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n108_), .B(new_new_n89_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n342_), .B(new_new_n518_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n430_), .B(new_new_n81_), .Y(new_new_n520_));
  NA2        g498(.A(i_11_), .B(new_new_n186_), .Y(new_new_n521_));
  INV        g499(.A(new_new_n519_), .Y(new_new_n522_));
  NA3        g500(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n523_));
  NO2        g501(.A(new_new_n220_), .B(i_4_), .Y(new_new_n524_));
  NA2        g502(.A(new_new_n524_), .B(i_8_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n105_), .B(new_new_n523_), .Y(new_new_n526_));
  NA2        g504(.A(i_2_), .B(new_new_n83_), .Y(new_new_n527_));
  OAI210     g505(.A0(new_new_n86_), .A1(new_new_n192_), .B0(new_new_n193_), .Y(new_new_n528_));
  NO2        g506(.A(i_7_), .B(new_new_n37_), .Y(new_new_n529_));
  NA2        g507(.A(i_4_), .B(i_8_), .Y(new_new_n530_));
  AOI210     g508(.A0(new_new_n530_), .A1(new_new_n278_), .B0(new_new_n529_), .Y(new_new_n531_));
  OAI220     g509(.A0(new_new_n531_), .A1(new_new_n527_), .B0(new_new_n528_), .B1(i_13_), .Y(new_new_n532_));
  NO4        g510(.A(new_new_n532_), .B(new_new_n526_), .C(new_new_n522_), .D(new_new_n517_), .Y(new_new_n533_));
  AOI210     g511(.A0(new_new_n128_), .A1(new_new_n61_), .B0(i_10_), .Y(new_new_n534_));
  AOI210     g512(.A0(new_new_n534_), .A1(new_new_n220_), .B0(new_new_n159_), .Y(new_new_n535_));
  OR2        g513(.A(i_6_), .B(i_10_), .Y(new_new_n536_));
  OR3        g514(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n537_));
  INV        g515(.A(new_new_n191_), .Y(new_new_n538_));
  OR2        g516(.A(new_new_n535_), .B(new_new_n242_), .Y(new_new_n539_));
  AOI210     g517(.A0(new_new_n539_), .A1(new_new_n533_), .B0(new_new_n62_), .Y(new_new_n540_));
  NOi21      g518(.An(i_11_), .B(i_7_), .Y(new_new_n541_));
  AO210      g519(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n542_));
  NO2        g520(.A(new_new_n542_), .B(new_new_n541_), .Y(new_new_n543_));
  NA2        g521(.A(new_new_n543_), .B(new_new_n197_), .Y(new_new_n544_));
  NA3        g522(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n545_));
  NAi31      g523(.An(new_new_n545_), .B(new_new_n204_), .C(i_11_), .Y(new_new_n546_));
  AOI210     g524(.A0(new_new_n546_), .A1(new_new_n544_), .B0(new_new_n62_), .Y(new_new_n547_));
  NA2        g525(.A(new_new_n85_), .B(new_new_n62_), .Y(new_new_n548_));
  AO210      g526(.A0(new_new_n548_), .A1(new_new_n336_), .B0(new_new_n41_), .Y(new_new_n549_));
  NO3        g527(.A(new_new_n235_), .B(new_new_n198_), .C(new_new_n521_), .Y(new_new_n550_));
  OAI210     g528(.A0(new_new_n550_), .A1(new_new_n213_), .B0(new_new_n62_), .Y(new_new_n551_));
  NA2        g529(.A(new_new_n369_), .B(new_new_n31_), .Y(new_new_n552_));
  OR2        g530(.A(new_new_n198_), .B(new_new_n108_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n553_), .B(new_new_n552_), .Y(new_new_n554_));
  NO2        g532(.A(i_1_), .B(i_4_), .Y(new_new_n555_));
  NA2        g533(.A(new_new_n555_), .B(new_new_n554_), .Y(new_new_n556_));
  NO2        g534(.A(i_1_), .B(i_12_), .Y(new_new_n557_));
  NA3        g535(.A(new_new_n557_), .B(new_new_n109_), .C(new_new_n24_), .Y(new_new_n558_));
  BUFFER     g536(.A(new_new_n558_), .Y(new_new_n559_));
  NA4        g537(.A(new_new_n559_), .B(new_new_n556_), .C(new_new_n551_), .D(new_new_n549_), .Y(new_new_n560_));
  OAI210     g538(.A0(new_new_n560_), .A1(new_new_n547_), .B0(i_6_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n545_), .B(new_new_n108_), .Y(new_new_n562_));
  NA2        g540(.A(new_new_n562_), .B(new_new_n505_), .Y(new_new_n563_));
  NO2        g541(.A(new_new_n220_), .B(new_new_n83_), .Y(new_new_n564_));
  NO2        g542(.A(new_new_n564_), .B(i_11_), .Y(new_new_n565_));
  NA2        g543(.A(new_new_n563_), .B(new_new_n408_), .Y(new_new_n566_));
  NO3        g544(.A(new_new_n536_), .B(new_new_n218_), .C(new_new_n23_), .Y(new_new_n567_));
  NA3        g545(.A(new_new_n465_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n568_));
  INV        g546(.A(i_2_), .Y(new_new_n569_));
  NA2        g547(.A(new_new_n138_), .B(i_9_), .Y(new_new_n570_));
  NO2        g548(.A(new_new_n46_), .B(i_1_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n570_), .B(new_new_n569_), .Y(new_new_n572_));
  AOI210     g550(.A0(new_new_n427_), .A1(new_new_n376_), .B0(new_new_n224_), .Y(new_new_n573_));
  NO2        g551(.A(new_new_n573_), .B(new_new_n527_), .Y(new_new_n574_));
  NAi21      g552(.An(new_new_n568_), .B(new_new_n91_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n571_), .B(new_new_n241_), .Y(new_new_n576_));
  NO2        g554(.A(i_11_), .B(new_new_n37_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n577_), .B(new_new_n24_), .Y(new_new_n578_));
  OAI210     g556(.A0(new_new_n578_), .A1(new_new_n576_), .B0(new_new_n575_), .Y(new_new_n579_));
  OR3        g557(.A(new_new_n579_), .B(new_new_n574_), .C(new_new_n572_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n580_), .B(new_new_n566_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n220_), .B(new_new_n101_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n582_), .B(new_new_n541_), .Y(new_new_n583_));
  NA2        g561(.A(new_new_n583_), .B(i_1_), .Y(new_new_n584_));
  NO2        g562(.A(new_new_n584_), .B(new_new_n537_), .Y(new_new_n585_));
  NO2        g563(.A(new_new_n372_), .B(new_new_n83_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n585_), .B(new_new_n46_), .Y(new_new_n587_));
  NA2        g565(.A(i_3_), .B(new_new_n186_), .Y(new_new_n588_));
  NO2        g566(.A(new_new_n588_), .B(new_new_n114_), .Y(new_new_n589_));
  AN2        g567(.A(new_new_n589_), .B(new_new_n470_), .Y(new_new_n590_));
  NO2        g568(.A(new_new_n218_), .B(new_new_n44_), .Y(new_new_n591_));
  NO3        g569(.A(new_new_n591_), .B(new_new_n280_), .C(new_new_n221_), .Y(new_new_n592_));
  NO2        g570(.A(new_new_n117_), .B(new_new_n37_), .Y(new_new_n593_));
  NO2        g571(.A(new_new_n593_), .B(i_6_), .Y(new_new_n594_));
  NO2        g572(.A(new_new_n83_), .B(i_9_), .Y(new_new_n595_));
  NO2        g573(.A(new_new_n595_), .B(new_new_n62_), .Y(new_new_n596_));
  NO2        g574(.A(new_new_n596_), .B(new_new_n557_), .Y(new_new_n597_));
  NO4        g575(.A(new_new_n597_), .B(new_new_n594_), .C(new_new_n592_), .D(i_4_), .Y(new_new_n598_));
  NA2        g576(.A(i_1_), .B(i_3_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n409_), .B(new_new_n92_), .Y(new_new_n600_));
  AOI210     g578(.A0(new_new_n591_), .A1(new_new_n493_), .B0(new_new_n600_), .Y(new_new_n601_));
  NO2        g579(.A(new_new_n601_), .B(new_new_n599_), .Y(new_new_n602_));
  NO3        g580(.A(new_new_n602_), .B(new_new_n598_), .C(new_new_n590_), .Y(new_new_n603_));
  NA4        g581(.A(new_new_n603_), .B(new_new_n587_), .C(new_new_n581_), .D(new_new_n561_), .Y(new_new_n604_));
  NO3        g582(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n605_));
  NOi21      g583(.An(new_new_n605_), .B(i_10_), .Y(new_new_n606_));
  OA210      g584(.A0(new_new_n606_), .A1(new_new_n228_), .B0(new_new_n83_), .Y(new_new_n607_));
  NO3        g585(.A(new_new_n428_), .B(new_new_n530_), .C(new_new_n83_), .Y(new_new_n608_));
  NA2        g586(.A(new_new_n608_), .B(new_new_n25_), .Y(new_new_n609_));
  INV        g587(.A(new_new_n609_), .Y(new_new_n610_));
  OAI210     g588(.A0(new_new_n610_), .A1(new_new_n607_), .B0(i_1_), .Y(new_new_n611_));
  AOI210     g589(.A0(new_new_n241_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n326_), .B(i_2_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n613_), .B(new_new_n612_), .Y(new_new_n614_));
  AOI210     g592(.A0(new_new_n614_), .A1(new_new_n611_), .B0(i_13_), .Y(new_new_n615_));
  OR2        g593(.A(i_11_), .B(i_7_), .Y(new_new_n616_));
  NA3        g594(.A(new_new_n616_), .B(new_new_n106_), .C(new_new_n138_), .Y(new_new_n617_));
  AOI220     g595(.A0(new_new_n423_), .A1(new_new_n159_), .B0(new_new_n402_), .B1(new_new_n138_), .Y(new_new_n618_));
  OAI210     g596(.A0(new_new_n618_), .A1(new_new_n44_), .B0(new_new_n617_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n54_), .B(i_12_), .Y(new_new_n620_));
  NO2        g598(.A(new_new_n428_), .B(new_new_n24_), .Y(new_new_n621_));
  NA2        g599(.A(new_new_n621_), .B(new_new_n586_), .Y(new_new_n622_));
  OAI220     g600(.A0(new_new_n622_), .A1(new_new_n41_), .B0(new_new_n924_), .B1(new_new_n92_), .Y(new_new_n623_));
  AOI210     g601(.A0(new_new_n619_), .A1(new_new_n301_), .B0(new_new_n623_), .Y(new_new_n624_));
  NA2        g602(.A(new_new_n344_), .B(new_new_n571_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(new_new_n225_), .Y(new_new_n626_));
  AOI210     g604(.A0(new_new_n400_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n627_));
  NOi31      g605(.An(new_new_n627_), .B(new_new_n520_), .C(new_new_n44_), .Y(new_new_n628_));
  NA2        g606(.A(new_new_n127_), .B(i_13_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n629_), .B(new_new_n612_), .Y(new_new_n630_));
  NO3        g608(.A(new_new_n70_), .B(new_new_n32_), .C(new_new_n101_), .Y(new_new_n631_));
  NA2        g609(.A(new_new_n26_), .B(new_new_n186_), .Y(new_new_n632_));
  NA2        g610(.A(new_new_n632_), .B(i_7_), .Y(new_new_n633_));
  AOI220     g611(.A0(new_new_n344_), .A1(new_new_n571_), .B0(new_new_n91_), .B1(new_new_n102_), .Y(new_new_n634_));
  OAI220     g612(.A0(new_new_n634_), .A1(new_new_n525_), .B0(new_new_n925_), .B1(new_new_n538_), .Y(new_new_n635_));
  NO4        g613(.A(new_new_n635_), .B(new_new_n630_), .C(new_new_n628_), .D(new_new_n626_), .Y(new_new_n636_));
  OR2        g614(.A(i_11_), .B(i_6_), .Y(new_new_n637_));
  NA3        g615(.A(new_new_n524_), .B(new_new_n632_), .C(i_7_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n638_), .B(new_new_n637_), .Y(new_new_n639_));
  NA3        g617(.A(new_new_n369_), .B(new_new_n529_), .C(new_new_n97_), .Y(new_new_n640_));
  NA2        g618(.A(new_new_n565_), .B(i_13_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n102_), .B(new_new_n632_), .Y(new_new_n642_));
  NAi21      g620(.An(i_11_), .B(i_12_), .Y(new_new_n643_));
  NOi41      g621(.An(new_new_n110_), .B(new_new_n643_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n644_));
  NO3        g622(.A(new_new_n428_), .B(new_new_n505_), .C(new_new_n530_), .Y(new_new_n645_));
  AOI220     g623(.A0(new_new_n645_), .A1(new_new_n283_), .B0(new_new_n644_), .B1(new_new_n642_), .Y(new_new_n646_));
  NA3        g624(.A(new_new_n646_), .B(new_new_n641_), .C(new_new_n640_), .Y(new_new_n647_));
  OAI210     g625(.A0(new_new_n647_), .A1(new_new_n639_), .B0(new_new_n62_), .Y(new_new_n648_));
  NO2        g626(.A(i_2_), .B(i_12_), .Y(new_new_n649_));
  NA2        g627(.A(new_new_n325_), .B(new_new_n649_), .Y(new_new_n650_));
  NO2        g628(.A(new_new_n128_), .B(i_2_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n651_), .B(new_new_n557_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n652_), .B(new_new_n650_), .Y(new_new_n653_));
  NA3        g631(.A(new_new_n653_), .B(new_new_n45_), .C(new_new_n212_), .Y(new_new_n654_));
  NA4        g632(.A(new_new_n654_), .B(new_new_n648_), .C(new_new_n636_), .D(new_new_n624_), .Y(new_new_n655_));
  OR4        g633(.A(new_new_n655_), .B(new_new_n615_), .C(new_new_n604_), .D(new_new_n540_), .Y(ori5));
  NA2        g634(.A(new_new_n583_), .B(new_new_n244_), .Y(new_new_n657_));
  AN2        g635(.A(new_new_n24_), .B(i_10_), .Y(new_new_n658_));
  NA3        g636(.A(new_new_n658_), .B(new_new_n649_), .C(new_new_n108_), .Y(new_new_n659_));
  NO2        g637(.A(new_new_n525_), .B(i_11_), .Y(new_new_n660_));
  NA2        g638(.A(new_new_n86_), .B(new_new_n660_), .Y(new_new_n661_));
  NA3        g639(.A(new_new_n661_), .B(new_new_n659_), .C(new_new_n657_), .Y(new_new_n662_));
  NO3        g640(.A(i_11_), .B(new_new_n220_), .C(i_13_), .Y(new_new_n663_));
  NO2        g641(.A(new_new_n124_), .B(new_new_n23_), .Y(new_new_n664_));
  NA2        g642(.A(i_12_), .B(i_8_), .Y(new_new_n665_));
  OAI210     g643(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n665_), .Y(new_new_n666_));
  INV        g644(.A(new_new_n399_), .Y(new_new_n667_));
  AOI220     g645(.A0(new_new_n289_), .A1(new_new_n497_), .B0(new_new_n666_), .B1(new_new_n664_), .Y(new_new_n668_));
  INV        g646(.A(new_new_n668_), .Y(new_new_n669_));
  NO2        g647(.A(new_new_n669_), .B(new_new_n662_), .Y(new_new_n670_));
  INV        g648(.A(new_new_n168_), .Y(new_new_n671_));
  INV        g649(.A(new_new_n228_), .Y(new_new_n672_));
  OAI210     g650(.A0(new_new_n613_), .A1(new_new_n401_), .B0(new_new_n110_), .Y(new_new_n673_));
  AOI210     g651(.A0(new_new_n673_), .A1(new_new_n672_), .B0(new_new_n671_), .Y(new_new_n674_));
  NO2        g652(.A(new_new_n409_), .B(new_new_n26_), .Y(new_new_n675_));
  NO2        g653(.A(new_new_n675_), .B(new_new_n376_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n676_), .B(i_2_), .Y(new_new_n677_));
  INV        g655(.A(new_new_n677_), .Y(new_new_n678_));
  AOI210     g656(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n373_), .Y(new_new_n679_));
  AOI210     g657(.A0(new_new_n679_), .A1(new_new_n678_), .B0(new_new_n674_), .Y(new_new_n680_));
  NO2        g658(.A(new_new_n184_), .B(new_new_n125_), .Y(new_new_n681_));
  OAI210     g659(.A0(new_new_n681_), .A1(new_new_n664_), .B0(i_2_), .Y(new_new_n682_));
  INV        g660(.A(new_new_n169_), .Y(new_new_n683_));
  NO3        g661(.A(new_new_n542_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n684_));
  AOI210     g662(.A0(new_new_n683_), .A1(new_new_n86_), .B0(new_new_n684_), .Y(new_new_n685_));
  AOI210     g663(.A0(new_new_n685_), .A1(new_new_n682_), .B0(new_new_n186_), .Y(new_new_n686_));
  OA210      g664(.A0(new_new_n543_), .A1(new_new_n126_), .B0(i_13_), .Y(new_new_n687_));
  NA2        g665(.A(new_new_n191_), .B(new_new_n192_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n151_), .B(new_new_n521_), .Y(new_new_n689_));
  AOI210     g667(.A0(new_new_n689_), .A1(new_new_n688_), .B0(new_new_n330_), .Y(new_new_n690_));
  AOI210     g668(.A0(new_new_n198_), .A1(new_new_n148_), .B0(new_new_n456_), .Y(new_new_n691_));
  NA2        g669(.A(new_new_n691_), .B(new_new_n376_), .Y(new_new_n692_));
  NO2        g670(.A(new_new_n102_), .B(new_new_n44_), .Y(new_new_n693_));
  INV        g671(.A(new_new_n276_), .Y(new_new_n694_));
  NA4        g672(.A(new_new_n694_), .B(new_new_n278_), .C(new_new_n124_), .D(new_new_n42_), .Y(new_new_n695_));
  OAI210     g673(.A0(new_new_n695_), .A1(new_new_n693_), .B0(new_new_n692_), .Y(new_new_n696_));
  NO4        g674(.A(new_new_n696_), .B(new_new_n690_), .C(new_new_n687_), .D(new_new_n686_), .Y(new_new_n697_));
  NA2        g675(.A(new_new_n497_), .B(new_new_n28_), .Y(new_new_n698_));
  NA2        g676(.A(new_new_n663_), .B(new_new_n251_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n699_), .B(new_new_n698_), .Y(new_new_n700_));
  NO2        g678(.A(new_new_n61_), .B(i_12_), .Y(new_new_n701_));
  NO2        g679(.A(new_new_n701_), .B(new_new_n126_), .Y(new_new_n702_));
  NO2        g680(.A(new_new_n702_), .B(new_new_n521_), .Y(new_new_n703_));
  AOI220     g681(.A0(new_new_n703_), .A1(new_new_n36_), .B0(new_new_n700_), .B1(new_new_n46_), .Y(new_new_n704_));
  NA4        g682(.A(new_new_n704_), .B(new_new_n697_), .C(new_new_n680_), .D(new_new_n670_), .Y(ori6));
  NO3        g683(.A(i_9_), .B(new_new_n279_), .C(i_1_), .Y(new_new_n706_));
  NA2        g684(.A(new_new_n706_), .B(new_new_n651_), .Y(new_new_n707_));
  NA4        g685(.A(new_new_n348_), .B(new_new_n429_), .C(new_new_n70_), .D(new_new_n101_), .Y(new_new_n708_));
  INV        g686(.A(new_new_n708_), .Y(new_new_n709_));
  NO2        g687(.A(new_new_n207_), .B(new_new_n432_), .Y(new_new_n710_));
  NO2        g688(.A(new_new_n709_), .B(new_new_n296_), .Y(new_new_n711_));
  AO210      g689(.A0(new_new_n711_), .A1(new_new_n707_), .B0(i_12_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n505_), .B(new_new_n62_), .Y(new_new_n713_));
  NA2        g691(.A(new_new_n606_), .B(new_new_n70_), .Y(new_new_n714_));
  BUFFER     g692(.A(new_new_n548_), .Y(new_new_n715_));
  NA3        g693(.A(new_new_n715_), .B(new_new_n714_), .C(new_new_n713_), .Y(new_new_n716_));
  NA2        g694(.A(new_new_n716_), .B(new_new_n72_), .Y(new_new_n717_));
  INV        g695(.A(new_new_n295_), .Y(new_new_n718_));
  NA2        g696(.A(new_new_n74_), .B(new_new_n131_), .Y(new_new_n719_));
  INV        g697(.A(new_new_n124_), .Y(new_new_n720_));
  NA2        g698(.A(new_new_n720_), .B(new_new_n46_), .Y(new_new_n721_));
  AOI210     g699(.A0(new_new_n721_), .A1(new_new_n719_), .B0(new_new_n718_), .Y(new_new_n722_));
  NO2        g700(.A(new_new_n231_), .B(i_9_), .Y(new_new_n723_));
  NA2        g701(.A(new_new_n723_), .B(new_new_n701_), .Y(new_new_n724_));
  AOI210     g702(.A0(new_new_n724_), .A1(new_new_n454_), .B0(new_new_n180_), .Y(new_new_n725_));
  NO2        g703(.A(new_new_n32_), .B(i_11_), .Y(new_new_n726_));
  NA3        g704(.A(new_new_n726_), .B(new_new_n426_), .C(new_new_n348_), .Y(new_new_n727_));
  NAi32      g705(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n728_));
  NO2        g706(.A(new_new_n637_), .B(new_new_n728_), .Y(new_new_n729_));
  OAI210     g707(.A0(new_new_n605_), .A1(new_new_n488_), .B0(new_new_n487_), .Y(new_new_n730_));
  NAi31      g708(.An(new_new_n729_), .B(new_new_n730_), .C(new_new_n727_), .Y(new_new_n731_));
  OR3        g709(.A(new_new_n731_), .B(new_new_n725_), .C(new_new_n722_), .Y(new_new_n732_));
  NO2        g710(.A(new_new_n616_), .B(i_2_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n734_));
  NO2        g712(.A(new_new_n734_), .B(new_new_n368_), .Y(new_new_n735_));
  NA2        g713(.A(new_new_n735_), .B(new_new_n733_), .Y(new_new_n736_));
  OR2        g714(.A(new_new_n543_), .B(new_new_n401_), .Y(new_new_n737_));
  NA3        g715(.A(new_new_n737_), .B(new_new_n147_), .C(new_new_n68_), .Y(new_new_n738_));
  AO210      g716(.A0(new_new_n439_), .A1(new_new_n667_), .B0(new_new_n36_), .Y(new_new_n739_));
  NA3        g717(.A(new_new_n739_), .B(new_new_n738_), .C(new_new_n736_), .Y(new_new_n740_));
  OAI210     g718(.A0(new_new_n564_), .A1(i_11_), .B0(new_new_n84_), .Y(new_new_n741_));
  AOI220     g719(.A0(new_new_n741_), .A1(new_new_n487_), .B0(new_new_n710_), .B1(new_new_n633_), .Y(new_new_n742_));
  NA3        g720(.A(new_new_n330_), .B(new_new_n222_), .C(new_new_n147_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n356_), .B(new_new_n69_), .Y(new_new_n744_));
  NA4        g722(.A(new_new_n744_), .B(new_new_n743_), .C(new_new_n742_), .D(new_new_n528_), .Y(new_new_n745_));
  AO210      g723(.A0(new_new_n456_), .A1(new_new_n46_), .B0(new_new_n85_), .Y(new_new_n746_));
  NA3        g724(.A(new_new_n746_), .B(new_new_n430_), .C(new_new_n206_), .Y(new_new_n747_));
  NA2        g725(.A(new_new_n401_), .B(new_new_n399_), .Y(new_new_n748_));
  NO2        g726(.A(new_new_n536_), .B(new_new_n102_), .Y(new_new_n749_));
  OAI210     g727(.A0(new_new_n749_), .A1(new_new_n111_), .B0(new_new_n367_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n227_), .B(new_new_n46_), .Y(new_new_n751_));
  INV        g729(.A(new_new_n510_), .Y(new_new_n752_));
  NA3        g730(.A(new_new_n752_), .B(new_new_n295_), .C(i_7_), .Y(new_new_n753_));
  NA4        g731(.A(new_new_n753_), .B(new_new_n750_), .C(new_new_n748_), .D(new_new_n747_), .Y(new_new_n754_));
  NO4        g732(.A(new_new_n754_), .B(new_new_n745_), .C(new_new_n740_), .D(new_new_n732_), .Y(new_new_n755_));
  NA4        g733(.A(new_new_n755_), .B(new_new_n717_), .C(new_new_n712_), .D(new_new_n338_), .Y(ori3));
  NA3        g734(.A(new_new_n743_), .B(new_new_n528_), .C(new_new_n329_), .Y(new_new_n757_));
  NA2        g735(.A(new_new_n757_), .B(new_new_n40_), .Y(new_new_n758_));
  NOi21      g736(.An(new_new_n96_), .B(new_new_n676_), .Y(new_new_n759_));
  NO3        g737(.A(new_new_n553_), .B(new_new_n409_), .C(new_new_n131_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n369_), .B(new_new_n45_), .Y(new_new_n761_));
  AN2        g739(.A(new_new_n407_), .B(new_new_n55_), .Y(new_new_n762_));
  NO3        g740(.A(new_new_n762_), .B(new_new_n760_), .C(new_new_n759_), .Y(new_new_n763_));
  AOI210     g741(.A0(new_new_n763_), .A1(new_new_n758_), .B0(new_new_n48_), .Y(new_new_n764_));
  NO4        g742(.A(new_new_n334_), .B(new_new_n341_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n765_));
  NA2        g743(.A(new_new_n180_), .B(new_new_n493_), .Y(new_new_n766_));
  NOi21      g744(.An(new_new_n766_), .B(new_new_n765_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n627_), .B(new_new_n595_), .Y(new_new_n768_));
  NA2        g746(.A(new_new_n302_), .B(new_new_n392_), .Y(new_new_n769_));
  OAI220     g747(.A0(new_new_n769_), .A1(new_new_n768_), .B0(new_new_n767_), .B1(new_new_n62_), .Y(new_new_n770_));
  NOi21      g748(.An(i_5_), .B(i_9_), .Y(new_new_n771_));
  NA2        g749(.A(new_new_n771_), .B(new_new_n398_), .Y(new_new_n772_));
  BUFFER     g750(.A(new_new_n241_), .Y(new_new_n773_));
  AOI210     g751(.A0(new_new_n773_), .A1(new_new_n427_), .B0(new_new_n608_), .Y(new_new_n774_));
  NO3        g752(.A(new_new_n370_), .B(new_new_n241_), .C(new_new_n72_), .Y(new_new_n775_));
  NO2        g753(.A(new_new_n171_), .B(new_new_n148_), .Y(new_new_n776_));
  AOI210     g754(.A0(new_new_n776_), .A1(new_new_n227_), .B0(new_new_n775_), .Y(new_new_n777_));
  OAI220     g755(.A0(new_new_n777_), .A1(new_new_n175_), .B0(new_new_n774_), .B1(new_new_n772_), .Y(new_new_n778_));
  NO3        g756(.A(new_new_n778_), .B(new_new_n770_), .C(new_new_n764_), .Y(new_new_n779_));
  NA2        g757(.A(new_new_n180_), .B(new_new_n24_), .Y(new_new_n780_));
  NO2        g758(.A(new_new_n593_), .B(new_new_n518_), .Y(new_new_n781_));
  NO2        g759(.A(new_new_n781_), .B(new_new_n780_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n283_), .B(new_new_n129_), .Y(new_new_n783_));
  NAi21      g761(.An(new_new_n160_), .B(new_new_n392_), .Y(new_new_n784_));
  OAI220     g762(.A0(new_new_n784_), .A1(new_new_n751_), .B0(new_new_n783_), .B1(new_new_n361_), .Y(new_new_n785_));
  NO2        g763(.A(new_new_n785_), .B(new_new_n782_), .Y(new_new_n786_));
  NA2        g764(.A(new_new_n494_), .B(i_0_), .Y(new_new_n787_));
  NO3        g765(.A(new_new_n787_), .B(new_new_n343_), .C(new_new_n86_), .Y(new_new_n788_));
  NO4        g766(.A(new_new_n509_), .B(new_new_n204_), .C(new_new_n373_), .D(new_new_n368_), .Y(new_new_n789_));
  AOI210     g767(.A0(new_new_n789_), .A1(i_11_), .B0(new_new_n788_), .Y(new_new_n790_));
  INV        g768(.A(new_new_n426_), .Y(new_new_n791_));
  AN2        g769(.A(new_new_n96_), .B(new_new_n226_), .Y(new_new_n792_));
  NA2        g770(.A(new_new_n663_), .B(new_new_n296_), .Y(new_new_n793_));
  AOI210     g771(.A0(new_new_n430_), .A1(new_new_n86_), .B0(new_new_n57_), .Y(new_new_n794_));
  OAI220     g772(.A0(new_new_n794_), .A1(new_new_n793_), .B0(new_new_n578_), .B1(new_new_n467_), .Y(new_new_n795_));
  NO2        g773(.A(new_new_n233_), .B(new_new_n152_), .Y(new_new_n796_));
  NA2        g774(.A(i_0_), .B(i_10_), .Y(new_new_n797_));
  INV        g775(.A(new_new_n469_), .Y(new_new_n798_));
  NO4        g776(.A(new_new_n114_), .B(new_new_n57_), .C(new_new_n588_), .D(i_5_), .Y(new_new_n799_));
  AO220      g777(.A0(new_new_n799_), .A1(new_new_n798_), .B0(new_new_n796_), .B1(i_6_), .Y(new_new_n800_));
  NA2        g778(.A(new_new_n183_), .B(new_new_n192_), .Y(new_new_n801_));
  NO2        g779(.A(new_new_n801_), .B(new_new_n793_), .Y(new_new_n802_));
  NO4        g780(.A(new_new_n802_), .B(new_new_n800_), .C(new_new_n795_), .D(new_new_n792_), .Y(new_new_n803_));
  NA3        g781(.A(new_new_n803_), .B(new_new_n790_), .C(new_new_n786_), .Y(new_new_n804_));
  NO2        g782(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n805_));
  NA2        g783(.A(i_11_), .B(i_9_), .Y(new_new_n806_));
  NO3        g784(.A(i_12_), .B(new_new_n806_), .C(new_new_n527_), .Y(new_new_n807_));
  AN2        g785(.A(new_new_n807_), .B(new_new_n805_), .Y(new_new_n808_));
  NO2        g786(.A(new_new_n48_), .B(i_7_), .Y(new_new_n809_));
  NA2        g787(.A(new_new_n353_), .B(new_new_n173_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n810_), .B(new_new_n158_), .Y(new_new_n811_));
  NO2        g789(.A(new_new_n171_), .B(i_0_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n811_), .B(new_new_n808_), .Y(new_new_n813_));
  NA2        g791(.A(new_new_n577_), .B(new_new_n121_), .Y(new_new_n814_));
  NO2        g792(.A(i_6_), .B(new_new_n814_), .Y(new_new_n815_));
  AOI210     g793(.A0(new_new_n400_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n816_));
  NA2        g794(.A(new_new_n168_), .B(new_new_n103_), .Y(new_new_n817_));
  NOi32      g795(.An(new_new_n816_), .Bn(new_new_n183_), .C(new_new_n817_), .Y(new_new_n818_));
  NA2        g796(.A(new_new_n529_), .B(new_new_n296_), .Y(new_new_n819_));
  NO2        g797(.A(new_new_n819_), .B(new_new_n761_), .Y(new_new_n820_));
  NO3        g798(.A(new_new_n820_), .B(new_new_n818_), .C(new_new_n815_), .Y(new_new_n821_));
  NOi21      g799(.An(i_7_), .B(i_5_), .Y(new_new_n822_));
  NOi31      g800(.An(new_new_n822_), .B(i_0_), .C(new_new_n643_), .Y(new_new_n823_));
  NA3        g801(.A(new_new_n823_), .B(new_new_n342_), .C(i_6_), .Y(new_new_n824_));
  OA210      g802(.A0(new_new_n817_), .A1(new_new_n454_), .B0(new_new_n824_), .Y(new_new_n825_));
  INV        g803(.A(new_new_n290_), .Y(new_new_n826_));
  NA3        g804(.A(new_new_n825_), .B(new_new_n821_), .C(new_new_n813_), .Y(new_new_n827_));
  OA210      g805(.A0(new_new_n426_), .A1(new_new_n210_), .B0(new_new_n425_), .Y(new_new_n828_));
  NA3        g806(.A(new_new_n425_), .B(new_new_n369_), .C(new_new_n45_), .Y(new_new_n829_));
  OAI210     g807(.A0(new_new_n784_), .A1(new_new_n791_), .B0(new_new_n829_), .Y(new_new_n830_));
  NO2        g808(.A(i_3_), .B(new_new_n182_), .Y(new_new_n831_));
  AOI220     g809(.A0(new_new_n831_), .A1(new_new_n426_), .B0(new_new_n830_), .B1(new_new_n72_), .Y(new_new_n832_));
  NA3        g810(.A(new_new_n734_), .B(new_new_n340_), .C(new_new_n564_), .Y(new_new_n833_));
  NA2        g811(.A(new_new_n92_), .B(new_new_n44_), .Y(new_new_n834_));
  NO2        g812(.A(new_new_n74_), .B(new_new_n665_), .Y(new_new_n835_));
  AOI220     g813(.A0(new_new_n835_), .A1(new_new_n834_), .B0(new_new_n170_), .B1(new_new_n518_), .Y(new_new_n836_));
  AOI210     g814(.A0(new_new_n836_), .A1(new_new_n833_), .B0(new_new_n47_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n837_), .B(new_new_n458_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n838_), .B(new_new_n832_), .Y(new_new_n839_));
  NO3        g817(.A(new_new_n839_), .B(new_new_n827_), .C(new_new_n804_), .Y(new_new_n840_));
  NO2        g818(.A(i_0_), .B(new_new_n643_), .Y(new_new_n841_));
  NA2        g819(.A(new_new_n72_), .B(new_new_n44_), .Y(new_new_n842_));
  AN2        g820(.A(new_new_n841_), .B(new_new_n170_), .Y(new_new_n843_));
  NO2        g821(.A(new_new_n713_), .B(new_new_n817_), .Y(new_new_n844_));
  AOI210     g822(.A0(new_new_n843_), .A1(new_new_n309_), .B0(new_new_n844_), .Y(new_new_n845_));
  NO2        g823(.A(new_new_n730_), .B(new_new_n362_), .Y(new_new_n846_));
  NA2        g824(.A(new_new_n227_), .B(new_new_n217_), .Y(new_new_n847_));
  AOI210     g825(.A0(new_new_n847_), .A1(new_new_n787_), .B0(new_new_n152_), .Y(new_new_n848_));
  NO2        g826(.A(new_new_n848_), .B(new_new_n846_), .Y(new_new_n849_));
  NA2        g827(.A(new_new_n849_), .B(new_new_n845_), .Y(new_new_n850_));
  NO3        g828(.A(new_new_n797_), .B(new_new_n771_), .C(new_new_n184_), .Y(new_new_n851_));
  AOI220     g829(.A0(new_new_n851_), .A1(i_11_), .B0(new_new_n490_), .B1(new_new_n74_), .Y(new_new_n852_));
  NO3        g830(.A(new_new_n199_), .B(new_new_n341_), .C(i_0_), .Y(new_new_n853_));
  OAI210     g831(.A0(new_new_n853_), .A1(new_new_n75_), .B0(i_13_), .Y(new_new_n854_));
  NA2        g832(.A(new_new_n854_), .B(new_new_n852_), .Y(new_new_n855_));
  AOI210     g833(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n171_), .Y(new_new_n856_));
  NA2        g834(.A(new_new_n856_), .B(new_new_n828_), .Y(new_new_n857_));
  INV        g835(.A(new_new_n475_), .Y(new_new_n858_));
  NO3        g836(.A(new_new_n761_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n859_));
  NA2        g837(.A(new_new_n438_), .B(new_new_n431_), .Y(new_new_n860_));
  NO3        g838(.A(new_new_n860_), .B(new_new_n859_), .C(new_new_n858_), .Y(new_new_n861_));
  NA3        g839(.A(new_new_n348_), .B(new_new_n168_), .C(new_new_n167_), .Y(new_new_n862_));
  NA3        g840(.A(new_new_n809_), .B(new_new_n266_), .C(new_new_n217_), .Y(new_new_n863_));
  NA2        g841(.A(new_new_n863_), .B(new_new_n862_), .Y(new_new_n864_));
  NA3        g842(.A(new_new_n348_), .B(new_new_n303_), .C(new_new_n208_), .Y(new_new_n865_));
  INV        g843(.A(new_new_n865_), .Y(new_new_n866_));
  NOi31      g844(.An(new_new_n347_), .B(new_new_n842_), .C(new_new_n223_), .Y(new_new_n867_));
  NO3        g845(.A(new_new_n806_), .B(new_new_n206_), .C(new_new_n184_), .Y(new_new_n868_));
  NO4        g846(.A(new_new_n868_), .B(new_new_n867_), .C(new_new_n866_), .D(new_new_n864_), .Y(new_new_n869_));
  NA3        g847(.A(new_new_n869_), .B(new_new_n861_), .C(new_new_n857_), .Y(new_new_n870_));
  NA3        g848(.A(new_new_n278_), .B(i_5_), .C(new_new_n186_), .Y(new_new_n871_));
  NAi31      g849(.An(new_new_n224_), .B(new_new_n871_), .C(new_new_n225_), .Y(new_new_n872_));
  NO4        g850(.A(new_new_n223_), .B(new_new_n199_), .C(i_0_), .D(i_12_), .Y(new_new_n873_));
  AOI220     g851(.A0(new_new_n873_), .A1(new_new_n872_), .B0(new_new_n709_), .B1(new_new_n172_), .Y(new_new_n874_));
  AN2        g852(.A(new_new_n797_), .B(new_new_n152_), .Y(new_new_n875_));
  NO4        g853(.A(new_new_n875_), .B(i_12_), .C(new_new_n568_), .D(new_new_n131_), .Y(new_new_n876_));
  NA2        g854(.A(new_new_n876_), .B(new_new_n206_), .Y(new_new_n877_));
  NA3        g855(.A(new_new_n98_), .B(new_new_n493_), .C(i_11_), .Y(new_new_n878_));
  NO2        g856(.A(new_new_n878_), .B(new_new_n154_), .Y(new_new_n879_));
  NA2        g857(.A(new_new_n822_), .B(new_new_n423_), .Y(new_new_n880_));
  NA2        g858(.A(new_new_n63_), .B(new_new_n101_), .Y(new_new_n881_));
  OAI220     g859(.A0(new_new_n881_), .A1(new_new_n871_), .B0(new_new_n880_), .B1(new_new_n596_), .Y(new_new_n882_));
  AOI210     g860(.A0(new_new_n882_), .A1(new_new_n812_), .B0(new_new_n879_), .Y(new_new_n883_));
  NA3        g861(.A(new_new_n883_), .B(new_new_n877_), .C(new_new_n874_), .Y(new_new_n884_));
  NO4        g862(.A(new_new_n884_), .B(new_new_n870_), .C(new_new_n855_), .D(new_new_n850_), .Y(new_new_n885_));
  OAI210     g863(.A0(new_new_n733_), .A1(new_new_n726_), .B0(new_new_n37_), .Y(new_new_n886_));
  NA3        g864(.A(new_new_n816_), .B(new_new_n325_), .C(i_5_), .Y(new_new_n887_));
  NA3        g865(.A(new_new_n887_), .B(new_new_n886_), .C(new_new_n535_), .Y(new_new_n888_));
  NA2        g866(.A(new_new_n888_), .B(new_new_n197_), .Y(new_new_n889_));
  AN2        g867(.A(new_new_n616_), .B(new_new_n326_), .Y(new_new_n890_));
  NA2        g868(.A(new_new_n181_), .B(new_new_n183_), .Y(new_new_n891_));
  AO210      g869(.A0(new_new_n890_), .A1(new_new_n33_), .B0(new_new_n891_), .Y(new_new_n892_));
  NAi31      g870(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n893_));
  AOI210     g871(.A0(new_new_n117_), .A1(new_new_n69_), .B0(new_new_n893_), .Y(new_new_n894_));
  NO2        g872(.A(new_new_n894_), .B(new_new_n567_), .Y(new_new_n895_));
  NA2        g873(.A(new_new_n895_), .B(new_new_n892_), .Y(new_new_n896_));
  NO2        g874(.A(new_new_n417_), .B(new_new_n241_), .Y(new_new_n897_));
  NO2        g875(.A(new_new_n897_), .B(new_new_n789_), .Y(new_new_n898_));
  OAI210     g876(.A0(new_new_n878_), .A1(new_new_n148_), .B0(new_new_n898_), .Y(new_new_n899_));
  AOI210     g877(.A0(new_new_n896_), .A1(new_new_n48_), .B0(new_new_n899_), .Y(new_new_n900_));
  AOI210     g878(.A0(new_new_n900_), .A1(new_new_n889_), .B0(new_new_n72_), .Y(new_new_n901_));
  INV        g879(.A(new_new_n337_), .Y(new_new_n902_));
  NO2        g880(.A(new_new_n902_), .B(new_new_n671_), .Y(new_new_n903_));
  OAI210     g881(.A0(new_new_n79_), .A1(new_new_n54_), .B0(new_new_n108_), .Y(new_new_n904_));
  NA2        g882(.A(new_new_n904_), .B(new_new_n75_), .Y(new_new_n905_));
  AOI210     g883(.A0(new_new_n856_), .A1(new_new_n809_), .B0(new_new_n823_), .Y(new_new_n906_));
  AOI210     g884(.A0(new_new_n906_), .A1(new_new_n905_), .B0(new_new_n599_), .Y(new_new_n907_));
  INV        g885(.A(new_new_n907_), .Y(new_new_n908_));
  OAI210     g886(.A0(new_new_n243_), .A1(new_new_n156_), .B0(new_new_n86_), .Y(new_new_n909_));
  NO2        g887(.A(new_new_n909_), .B(i_11_), .Y(new_new_n910_));
  NA2        g888(.A(new_new_n530_), .B(new_new_n204_), .Y(new_new_n911_));
  OAI210     g889(.A0(new_new_n911_), .A1(new_new_n816_), .B0(new_new_n197_), .Y(new_new_n912_));
  NA2        g890(.A(new_new_n162_), .B(i_5_), .Y(new_new_n913_));
  NO2        g891(.A(new_new_n912_), .B(new_new_n913_), .Y(new_new_n914_));
  NO3        g892(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n915_));
  OAI210     g893(.A0(new_new_n826_), .A1(new_new_n279_), .B0(new_new_n915_), .Y(new_new_n916_));
  NO2        g894(.A(new_new_n916_), .B(new_new_n643_), .Y(new_new_n917_));
  NO3        g895(.A(new_new_n917_), .B(new_new_n914_), .C(new_new_n910_), .Y(new_new_n918_));
  OAI210     g896(.A0(new_new_n908_), .A1(i_4_), .B0(new_new_n918_), .Y(new_new_n919_));
  NO3        g897(.A(new_new_n919_), .B(new_new_n903_), .C(new_new_n901_), .Y(new_new_n920_));
  NA4        g898(.A(new_new_n920_), .B(new_new_n885_), .C(new_new_n840_), .D(new_new_n779_), .Y(ori4));
  INV        g899(.A(new_new_n620_), .Y(new_new_n924_));
  INV        g900(.A(new_new_n631_), .Y(new_new_n925_));
endmodule


