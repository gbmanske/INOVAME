//Benchmark atmr_misex3_1774_0.0313

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1227_, ori_ori_n1228_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1522_, mai_mai_n1523_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1597_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  NO2        o0001(.A(d), .B(c), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NOi32      o0003(.An(m), .Bn(l), .C(n), .Y(ori_ori_n32_));
  NOi32      o0004(.An(i), .Bn(g), .C(h), .Y(ori_ori_n33_));
  NA2        o0005(.A(ori_ori_n33_), .B(ori_ori_n32_), .Y(ori_ori_n34_));
  AN2        o0006(.A(m), .B(l), .Y(ori_ori_n35_));
  NOi32      o0007(.An(j), .Bn(g), .C(k), .Y(ori_ori_n36_));
  NA2        o0008(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n37_));
  NO2        o0009(.A(ori_ori_n37_), .B(n), .Y(ori_ori_n38_));
  INV        o0010(.A(h), .Y(ori_ori_n39_));
  NAi21      o0011(.An(j), .B(l), .Y(ori_ori_n40_));
  NAi32      o0012(.An(n), .Bn(g), .C(m), .Y(ori_ori_n41_));
  NO3        o0013(.A(ori_ori_n41_), .B(ori_ori_n40_), .C(ori_ori_n39_), .Y(ori_ori_n42_));
  NAi31      o0014(.An(n), .B(m), .C(l), .Y(ori_ori_n43_));
  INV        o0015(.A(i), .Y(ori_ori_n44_));
  AN2        o0016(.A(h), .B(g), .Y(ori_ori_n45_));
  NA2        o0017(.A(ori_ori_n45_), .B(ori_ori_n44_), .Y(ori_ori_n46_));
  NO2        o0018(.A(ori_ori_n46_), .B(ori_ori_n43_), .Y(ori_ori_n47_));
  NAi21      o0019(.An(n), .B(m), .Y(ori_ori_n48_));
  NOi32      o0020(.An(k), .Bn(h), .C(l), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(g), .Y(ori_ori_n50_));
  INV        o0022(.A(ori_ori_n50_), .Y(ori_ori_n51_));
  NO2        o0023(.A(ori_ori_n51_), .B(ori_ori_n48_), .Y(ori_ori_n52_));
  INV        o0024(.A(c), .Y(ori_ori_n53_));
  NA2        o0025(.A(e), .B(b), .Y(ori_ori_n54_));
  NO2        o0026(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  INV        o0027(.A(d), .Y(ori_ori_n56_));
  NAi21      o0028(.An(i), .B(h), .Y(ori_ori_n57_));
  NAi41      o0029(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n58_));
  NA2        o0030(.A(g), .B(f), .Y(ori_ori_n59_));
  NAi21      o0031(.An(i), .B(j), .Y(ori_ori_n60_));
  NAi32      o0032(.An(n), .Bn(k), .C(m), .Y(ori_ori_n61_));
  NAi31      o0033(.An(l), .B(m), .C(k), .Y(ori_ori_n62_));
  NAi21      o0034(.An(e), .B(h), .Y(ori_ori_n63_));
  NAi41      o0035(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n64_));
  INV        o0036(.A(m), .Y(ori_ori_n65_));
  NOi21      o0037(.An(k), .B(l), .Y(ori_ori_n66_));
  NA2        o0038(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n67_));
  AN4        o0039(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n68_));
  NOi31      o0040(.An(h), .B(g), .C(f), .Y(ori_ori_n69_));
  NA2        o0041(.A(ori_ori_n69_), .B(ori_ori_n68_), .Y(ori_ori_n70_));
  NAi32      o0042(.An(m), .Bn(k), .C(j), .Y(ori_ori_n71_));
  NOi32      o0043(.An(h), .Bn(g), .C(f), .Y(ori_ori_n72_));
  NA2        o0044(.A(ori_ori_n72_), .B(ori_ori_n68_), .Y(ori_ori_n73_));
  OA220      o0045(.A0(ori_ori_n73_), .A1(ori_ori_n71_), .B0(ori_ori_n70_), .B1(ori_ori_n67_), .Y(ori_ori_n74_));
  INV        o0046(.A(ori_ori_n74_), .Y(ori_ori_n75_));
  INV        o0047(.A(n), .Y(ori_ori_n76_));
  NOi32      o0048(.An(e), .Bn(b), .C(d), .Y(ori_ori_n77_));
  NA2        o0049(.A(ori_ori_n77_), .B(ori_ori_n76_), .Y(ori_ori_n78_));
  INV        o0050(.A(j), .Y(ori_ori_n79_));
  AN3        o0051(.A(m), .B(k), .C(i), .Y(ori_ori_n80_));
  NA3        o0052(.A(ori_ori_n80_), .B(ori_ori_n79_), .C(g), .Y(ori_ori_n81_));
  NO2        o0053(.A(ori_ori_n81_), .B(f), .Y(ori_ori_n82_));
  NAi32      o0054(.An(g), .Bn(f), .C(h), .Y(ori_ori_n83_));
  NAi31      o0055(.An(j), .B(m), .C(l), .Y(ori_ori_n84_));
  NO2        o0056(.A(ori_ori_n84_), .B(ori_ori_n83_), .Y(ori_ori_n85_));
  NA2        o0057(.A(m), .B(l), .Y(ori_ori_n86_));
  NAi31      o0058(.An(k), .B(j), .C(g), .Y(ori_ori_n87_));
  NO3        o0059(.A(ori_ori_n87_), .B(ori_ori_n86_), .C(f), .Y(ori_ori_n88_));
  AN2        o0060(.A(j), .B(g), .Y(ori_ori_n89_));
  NOi32      o0061(.An(m), .Bn(l), .C(i), .Y(ori_ori_n90_));
  NOi21      o0062(.An(g), .B(i), .Y(ori_ori_n91_));
  NOi32      o0063(.An(m), .Bn(j), .C(k), .Y(ori_ori_n92_));
  AOI220     o0064(.A0(ori_ori_n92_), .A1(ori_ori_n91_), .B0(ori_ori_n90_), .B1(ori_ori_n89_), .Y(ori_ori_n93_));
  NO2        o0065(.A(ori_ori_n93_), .B(f), .Y(ori_ori_n94_));
  NO4        o0066(.A(ori_ori_n94_), .B(ori_ori_n88_), .C(ori_ori_n85_), .D(ori_ori_n82_), .Y(ori_ori_n95_));
  NAi41      o0067(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n96_));
  AN2        o0068(.A(e), .B(b), .Y(ori_ori_n97_));
  NOi31      o0069(.An(c), .B(h), .C(f), .Y(ori_ori_n98_));
  NA2        o0070(.A(ori_ori_n98_), .B(ori_ori_n97_), .Y(ori_ori_n99_));
  NO2        o0071(.A(ori_ori_n99_), .B(ori_ori_n96_), .Y(ori_ori_n100_));
  NOi21      o0072(.An(g), .B(f), .Y(ori_ori_n101_));
  NOi21      o0073(.An(i), .B(h), .Y(ori_ori_n102_));
  INV        o0074(.A(a), .Y(ori_ori_n103_));
  NA2        o0075(.A(ori_ori_n97_), .B(ori_ori_n103_), .Y(ori_ori_n104_));
  INV        o0076(.A(l), .Y(ori_ori_n105_));
  NOi21      o0077(.An(m), .B(n), .Y(ori_ori_n106_));
  AN2        o0078(.A(k), .B(h), .Y(ori_ori_n107_));
  INV        o0079(.A(b), .Y(ori_ori_n108_));
  NA2        o0080(.A(l), .B(j), .Y(ori_ori_n109_));
  AN2        o0081(.A(k), .B(i), .Y(ori_ori_n110_));
  NA2        o0082(.A(g), .B(e), .Y(ori_ori_n111_));
  NOi32      o0083(.An(c), .Bn(a), .C(d), .Y(ori_ori_n112_));
  NA2        o0084(.A(ori_ori_n112_), .B(ori_ori_n106_), .Y(ori_ori_n113_));
  INV        o0085(.A(ori_ori_n100_), .Y(ori_ori_n114_));
  OAI210     o0086(.A0(ori_ori_n95_), .A1(ori_ori_n78_), .B0(ori_ori_n114_), .Y(ori_ori_n115_));
  NOi31      o0087(.An(k), .B(m), .C(j), .Y(ori_ori_n116_));
  NA3        o0088(.A(ori_ori_n116_), .B(ori_ori_n69_), .C(ori_ori_n68_), .Y(ori_ori_n117_));
  NOi31      o0089(.An(k), .B(m), .C(i), .Y(ori_ori_n118_));
  INV        o0090(.A(ori_ori_n117_), .Y(ori_ori_n119_));
  NOi32      o0091(.An(f), .Bn(b), .C(e), .Y(ori_ori_n120_));
  NAi21      o0092(.An(g), .B(h), .Y(ori_ori_n121_));
  NAi21      o0093(.An(m), .B(n), .Y(ori_ori_n122_));
  NAi21      o0094(.An(j), .B(k), .Y(ori_ori_n123_));
  NO3        o0095(.A(ori_ori_n123_), .B(ori_ori_n122_), .C(ori_ori_n121_), .Y(ori_ori_n124_));
  NAi41      o0096(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n125_));
  NAi31      o0097(.An(j), .B(k), .C(h), .Y(ori_ori_n126_));
  NA2        o0098(.A(ori_ori_n124_), .B(ori_ori_n120_), .Y(ori_ori_n127_));
  NO2        o0099(.A(k), .B(j), .Y(ori_ori_n128_));
  NO2        o0100(.A(ori_ori_n128_), .B(ori_ori_n122_), .Y(ori_ori_n129_));
  AN2        o0101(.A(k), .B(j), .Y(ori_ori_n130_));
  NAi21      o0102(.An(c), .B(b), .Y(ori_ori_n131_));
  NA2        o0103(.A(f), .B(d), .Y(ori_ori_n132_));
  NO4        o0104(.A(ori_ori_n132_), .B(ori_ori_n131_), .C(ori_ori_n130_), .D(ori_ori_n121_), .Y(ori_ori_n133_));
  NA2        o0105(.A(h), .B(c), .Y(ori_ori_n134_));
  NAi31      o0106(.An(f), .B(e), .C(b), .Y(ori_ori_n135_));
  NA2        o0107(.A(ori_ori_n133_), .B(ori_ori_n129_), .Y(ori_ori_n136_));
  NA2        o0108(.A(d), .B(b), .Y(ori_ori_n137_));
  NAi21      o0109(.An(e), .B(f), .Y(ori_ori_n138_));
  NO2        o0110(.A(ori_ori_n138_), .B(ori_ori_n137_), .Y(ori_ori_n139_));
  NAi21      o0111(.An(e), .B(g), .Y(ori_ori_n140_));
  NAi21      o0112(.An(c), .B(d), .Y(ori_ori_n141_));
  NAi31      o0113(.An(l), .B(k), .C(h), .Y(ori_ori_n142_));
  NO2        o0114(.A(ori_ori_n122_), .B(ori_ori_n142_), .Y(ori_ori_n143_));
  NA2        o0115(.A(ori_ori_n143_), .B(ori_ori_n139_), .Y(ori_ori_n144_));
  NAi41      o0116(.An(ori_ori_n119_), .B(ori_ori_n144_), .C(ori_ori_n136_), .D(ori_ori_n127_), .Y(ori_ori_n145_));
  NAi31      o0117(.An(e), .B(f), .C(b), .Y(ori_ori_n146_));
  NOi21      o0118(.An(g), .B(d), .Y(ori_ori_n147_));
  NO2        o0119(.A(ori_ori_n147_), .B(ori_ori_n146_), .Y(ori_ori_n148_));
  NOi21      o0120(.An(h), .B(i), .Y(ori_ori_n149_));
  NOi21      o0121(.An(k), .B(m), .Y(ori_ori_n150_));
  NA3        o0122(.A(ori_ori_n150_), .B(ori_ori_n149_), .C(n), .Y(ori_ori_n151_));
  NOi21      o0123(.An(ori_ori_n148_), .B(ori_ori_n151_), .Y(ori_ori_n152_));
  NOi21      o0124(.An(h), .B(g), .Y(ori_ori_n153_));
  NAi31      o0125(.An(l), .B(j), .C(h), .Y(ori_ori_n154_));
  NOi32      o0126(.An(n), .Bn(k), .C(m), .Y(ori_ori_n155_));
  NAi31      o0127(.An(d), .B(f), .C(c), .Y(ori_ori_n156_));
  NAi31      o0128(.An(e), .B(f), .C(c), .Y(ori_ori_n157_));
  NA2        o0129(.A(ori_ori_n157_), .B(ori_ori_n156_), .Y(ori_ori_n158_));
  NA2        o0130(.A(j), .B(h), .Y(ori_ori_n159_));
  OR3        o0131(.A(n), .B(m), .C(k), .Y(ori_ori_n160_));
  NO2        o0132(.A(ori_ori_n160_), .B(ori_ori_n159_), .Y(ori_ori_n161_));
  NAi32      o0133(.An(m), .Bn(k), .C(n), .Y(ori_ori_n162_));
  NO2        o0134(.A(ori_ori_n162_), .B(ori_ori_n159_), .Y(ori_ori_n163_));
  AOI220     o0135(.A0(ori_ori_n163_), .A1(ori_ori_n148_), .B0(ori_ori_n161_), .B1(ori_ori_n158_), .Y(ori_ori_n164_));
  NO2        o0136(.A(n), .B(m), .Y(ori_ori_n165_));
  NA2        o0137(.A(ori_ori_n165_), .B(ori_ori_n49_), .Y(ori_ori_n166_));
  NAi21      o0138(.An(f), .B(e), .Y(ori_ori_n167_));
  NA2        o0139(.A(d), .B(c), .Y(ori_ori_n168_));
  NO2        o0140(.A(ori_ori_n168_), .B(ori_ori_n167_), .Y(ori_ori_n169_));
  NOi21      o0141(.An(ori_ori_n169_), .B(ori_ori_n166_), .Y(ori_ori_n170_));
  NAi31      o0142(.An(m), .B(n), .C(b), .Y(ori_ori_n171_));
  NA2        o0143(.A(k), .B(i), .Y(ori_ori_n172_));
  NAi21      o0144(.An(h), .B(f), .Y(ori_ori_n173_));
  NO2        o0145(.A(ori_ori_n173_), .B(ori_ori_n172_), .Y(ori_ori_n174_));
  NO2        o0146(.A(ori_ori_n171_), .B(ori_ori_n141_), .Y(ori_ori_n175_));
  NA2        o0147(.A(ori_ori_n175_), .B(ori_ori_n174_), .Y(ori_ori_n176_));
  NOi32      o0148(.An(f), .Bn(c), .C(d), .Y(ori_ori_n177_));
  NOi32      o0149(.An(f), .Bn(c), .C(e), .Y(ori_ori_n178_));
  NO2        o0150(.A(ori_ori_n178_), .B(ori_ori_n177_), .Y(ori_ori_n179_));
  NO3        o0151(.A(n), .B(m), .C(j), .Y(ori_ori_n180_));
  NA2        o0152(.A(ori_ori_n180_), .B(ori_ori_n107_), .Y(ori_ori_n181_));
  AO210      o0153(.A0(ori_ori_n181_), .A1(ori_ori_n166_), .B0(ori_ori_n179_), .Y(ori_ori_n182_));
  NAi41      o0154(.An(ori_ori_n170_), .B(ori_ori_n182_), .C(ori_ori_n176_), .D(ori_ori_n164_), .Y(ori_ori_n183_));
  OR3        o0155(.A(ori_ori_n183_), .B(ori_ori_n152_), .C(ori_ori_n145_), .Y(ori_ori_n184_));
  NO3        o0156(.A(ori_ori_n184_), .B(ori_ori_n115_), .C(ori_ori_n75_), .Y(ori_ori_n185_));
  NA3        o0157(.A(m), .B(ori_ori_n105_), .C(j), .Y(ori_ori_n186_));
  NAi31      o0158(.An(n), .B(h), .C(g), .Y(ori_ori_n187_));
  NO2        o0159(.A(ori_ori_n187_), .B(ori_ori_n186_), .Y(ori_ori_n188_));
  NOi32      o0160(.An(m), .Bn(k), .C(l), .Y(ori_ori_n189_));
  NA3        o0161(.A(ori_ori_n189_), .B(ori_ori_n79_), .C(g), .Y(ori_ori_n190_));
  NO2        o0162(.A(ori_ori_n190_), .B(n), .Y(ori_ori_n191_));
  NOi21      o0163(.An(k), .B(j), .Y(ori_ori_n192_));
  NA4        o0164(.A(ori_ori_n192_), .B(ori_ori_n106_), .C(i), .D(g), .Y(ori_ori_n193_));
  NAi41      o0165(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n194_));
  INV        o0166(.A(ori_ori_n194_), .Y(ori_ori_n195_));
  INV        o0167(.A(f), .Y(ori_ori_n196_));
  INV        o0168(.A(g), .Y(ori_ori_n197_));
  NOi31      o0169(.An(i), .B(j), .C(h), .Y(ori_ori_n198_));
  NOi21      o0170(.An(l), .B(m), .Y(ori_ori_n199_));
  NA2        o0171(.A(ori_ori_n199_), .B(ori_ori_n198_), .Y(ori_ori_n200_));
  NO3        o0172(.A(ori_ori_n200_), .B(ori_ori_n197_), .C(ori_ori_n196_), .Y(ori_ori_n201_));
  NA2        o0173(.A(ori_ori_n201_), .B(ori_ori_n195_), .Y(ori_ori_n202_));
  INV        o0174(.A(ori_ori_n202_), .Y(ori_ori_n203_));
  NOi21      o0175(.An(n), .B(m), .Y(ori_ori_n204_));
  OR2        o0176(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n205_));
  NAi21      o0177(.An(j), .B(h), .Y(ori_ori_n206_));
  XN2        o0178(.A(i), .B(h), .Y(ori_ori_n207_));
  NA2        o0179(.A(ori_ori_n207_), .B(ori_ori_n206_), .Y(ori_ori_n208_));
  NOi31      o0180(.An(k), .B(n), .C(m), .Y(ori_ori_n209_));
  NOi31      o0181(.An(ori_ori_n209_), .B(ori_ori_n168_), .C(ori_ori_n167_), .Y(ori_ori_n210_));
  NA2        o0182(.A(ori_ori_n210_), .B(ori_ori_n208_), .Y(ori_ori_n211_));
  NAi31      o0183(.An(f), .B(e), .C(c), .Y(ori_ori_n212_));
  NO4        o0184(.A(ori_ori_n212_), .B(ori_ori_n160_), .C(ori_ori_n159_), .D(ori_ori_n56_), .Y(ori_ori_n213_));
  NA3        o0185(.A(e), .B(c), .C(b), .Y(ori_ori_n214_));
  NAi32      o0186(.An(m), .Bn(i), .C(k), .Y(ori_ori_n215_));
  INV        o0187(.A(k), .Y(ori_ori_n216_));
  INV        o0188(.A(ori_ori_n213_), .Y(ori_ori_n217_));
  NAi21      o0189(.An(n), .B(a), .Y(ori_ori_n218_));
  NO2        o0190(.A(ori_ori_n218_), .B(ori_ori_n137_), .Y(ori_ori_n219_));
  NAi41      o0191(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n220_));
  NO2        o0192(.A(ori_ori_n220_), .B(e), .Y(ori_ori_n221_));
  NA2        o0193(.A(ori_ori_n221_), .B(ori_ori_n219_), .Y(ori_ori_n222_));
  AN4        o0194(.A(ori_ori_n222_), .B(ori_ori_n217_), .C(ori_ori_n211_), .D(ori_ori_n205_), .Y(ori_ori_n223_));
  OR2        o0195(.A(h), .B(g), .Y(ori_ori_n224_));
  NO2        o0196(.A(ori_ori_n224_), .B(ori_ori_n96_), .Y(ori_ori_n225_));
  NA2        o0197(.A(ori_ori_n225_), .B(ori_ori_n120_), .Y(ori_ori_n226_));
  NAi41      o0198(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n227_));
  NO2        o0199(.A(ori_ori_n227_), .B(ori_ori_n196_), .Y(ori_ori_n228_));
  NA2        o0200(.A(ori_ori_n150_), .B(ori_ori_n102_), .Y(ori_ori_n229_));
  NAi21      o0201(.An(ori_ori_n229_), .B(ori_ori_n228_), .Y(ori_ori_n230_));
  NO2        o0202(.A(n), .B(a), .Y(ori_ori_n231_));
  NAi31      o0203(.An(ori_ori_n220_), .B(ori_ori_n231_), .C(ori_ori_n97_), .Y(ori_ori_n232_));
  AN2        o0204(.A(ori_ori_n232_), .B(ori_ori_n230_), .Y(ori_ori_n233_));
  NAi21      o0205(.An(h), .B(i), .Y(ori_ori_n234_));
  NA2        o0206(.A(ori_ori_n165_), .B(k), .Y(ori_ori_n235_));
  NO2        o0207(.A(ori_ori_n235_), .B(ori_ori_n234_), .Y(ori_ori_n236_));
  NA2        o0208(.A(ori_ori_n236_), .B(ori_ori_n177_), .Y(ori_ori_n237_));
  NA3        o0209(.A(ori_ori_n237_), .B(ori_ori_n233_), .C(ori_ori_n226_), .Y(ori_ori_n238_));
  NOi21      o0210(.An(g), .B(e), .Y(ori_ori_n239_));
  NO2        o0211(.A(ori_ori_n64_), .B(ori_ori_n65_), .Y(ori_ori_n240_));
  NA2        o0212(.A(ori_ori_n240_), .B(ori_ori_n239_), .Y(ori_ori_n241_));
  NOi32      o0213(.An(l), .Bn(j), .C(i), .Y(ori_ori_n242_));
  AOI210     o0214(.A0(ori_ori_n66_), .A1(ori_ori_n79_), .B0(ori_ori_n242_), .Y(ori_ori_n243_));
  NAi21      o0215(.An(f), .B(g), .Y(ori_ori_n244_));
  NO2        o0216(.A(ori_ori_n244_), .B(ori_ori_n58_), .Y(ori_ori_n245_));
  NO2        o0217(.A(ori_ori_n243_), .B(ori_ori_n241_), .Y(ori_ori_n246_));
  NOi41      o0218(.An(ori_ori_n223_), .B(ori_ori_n246_), .C(ori_ori_n238_), .D(ori_ori_n203_), .Y(ori_ori_n247_));
  NO4        o0219(.A(ori_ori_n188_), .B(ori_ori_n47_), .C(ori_ori_n42_), .D(ori_ori_n38_), .Y(ori_ori_n248_));
  NO2        o0220(.A(ori_ori_n248_), .B(ori_ori_n104_), .Y(ori_ori_n249_));
  NA3        o0221(.A(ori_ori_n56_), .B(c), .C(b), .Y(ori_ori_n250_));
  NAi21      o0222(.An(h), .B(g), .Y(ori_ori_n251_));
  NO2        o0223(.A(ori_ori_n229_), .B(ori_ori_n244_), .Y(ori_ori_n252_));
  NAi31      o0224(.An(g), .B(k), .C(h), .Y(ori_ori_n253_));
  NA4        o0225(.A(ori_ori_n150_), .B(ori_ori_n72_), .C(ori_ori_n68_), .D(ori_ori_n109_), .Y(ori_ori_n254_));
  NA3        o0226(.A(ori_ori_n150_), .B(ori_ori_n149_), .C(ori_ori_n76_), .Y(ori_ori_n255_));
  NO2        o0227(.A(ori_ori_n255_), .B(ori_ori_n179_), .Y(ori_ori_n256_));
  NOi21      o0228(.An(ori_ori_n254_), .B(ori_ori_n256_), .Y(ori_ori_n257_));
  NA3        o0229(.A(e), .B(c), .C(b), .Y(ori_ori_n258_));
  NAi31      o0230(.An(h), .B(l), .C(i), .Y(ori_ori_n259_));
  NA2        o0231(.A(ori_ori_n259_), .B(ori_ori_n154_), .Y(ori_ori_n260_));
  NOi21      o0232(.An(ori_ori_n260_), .B(ori_ori_n48_), .Y(ori_ori_n261_));
  NA2        o0233(.A(ori_ori_n245_), .B(ori_ori_n261_), .Y(ori_ori_n262_));
  NAi21      o0234(.An(l), .B(k), .Y(ori_ori_n263_));
  NO2        o0235(.A(ori_ori_n263_), .B(ori_ori_n48_), .Y(ori_ori_n264_));
  NOi21      o0236(.An(l), .B(j), .Y(ori_ori_n265_));
  NA2        o0237(.A(ori_ori_n153_), .B(ori_ori_n265_), .Y(ori_ori_n266_));
  NAi32      o0238(.An(j), .Bn(h), .C(i), .Y(ori_ori_n267_));
  NAi21      o0239(.An(m), .B(l), .Y(ori_ori_n268_));
  NO3        o0240(.A(ori_ori_n268_), .B(ori_ori_n267_), .C(ori_ori_n76_), .Y(ori_ori_n269_));
  NA2        o0241(.A(h), .B(g), .Y(ori_ori_n270_));
  NA2        o0242(.A(ori_ori_n262_), .B(ori_ori_n257_), .Y(ori_ori_n271_));
  NO2        o0243(.A(ori_ori_n135_), .B(d), .Y(ori_ori_n272_));
  NA2        o0244(.A(ori_ori_n272_), .B(ori_ori_n52_), .Y(ori_ori_n273_));
  NO2        o0245(.A(ori_ori_n99_), .B(ori_ori_n96_), .Y(ori_ori_n274_));
  NAi32      o0246(.An(n), .Bn(m), .C(l), .Y(ori_ori_n275_));
  NO2        o0247(.A(ori_ori_n275_), .B(ori_ori_n267_), .Y(ori_ori_n276_));
  NA2        o0248(.A(ori_ori_n276_), .B(ori_ori_n169_), .Y(ori_ori_n277_));
  NAi31      o0249(.An(k), .B(l), .C(j), .Y(ori_ori_n278_));
  OAI210     o0250(.A0(ori_ori_n263_), .A1(j), .B0(ori_ori_n278_), .Y(ori_ori_n279_));
  NOi21      o0251(.An(ori_ori_n279_), .B(ori_ori_n111_), .Y(ori_ori_n280_));
  NA2        o0252(.A(ori_ori_n277_), .B(ori_ori_n273_), .Y(ori_ori_n281_));
  NO3        o0253(.A(ori_ori_n281_), .B(ori_ori_n271_), .C(ori_ori_n249_), .Y(ori_ori_n282_));
  NA2        o0254(.A(ori_ori_n236_), .B(ori_ori_n178_), .Y(ori_ori_n283_));
  NAi21      o0255(.An(m), .B(k), .Y(ori_ori_n284_));
  NO2        o0256(.A(ori_ori_n207_), .B(ori_ori_n284_), .Y(ori_ori_n285_));
  NAi41      o0257(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n286_));
  NO2        o0258(.A(ori_ori_n286_), .B(ori_ori_n140_), .Y(ori_ori_n287_));
  NA2        o0259(.A(ori_ori_n287_), .B(ori_ori_n285_), .Y(ori_ori_n288_));
  NA2        o0260(.A(e), .B(c), .Y(ori_ori_n289_));
  NO3        o0261(.A(ori_ori_n289_), .B(n), .C(d), .Y(ori_ori_n290_));
  NOi21      o0262(.An(f), .B(h), .Y(ori_ori_n291_));
  NA2        o0263(.A(ori_ori_n291_), .B(ori_ori_n110_), .Y(ori_ori_n292_));
  NO2        o0264(.A(ori_ori_n292_), .B(ori_ori_n197_), .Y(ori_ori_n293_));
  NAi31      o0265(.An(d), .B(e), .C(b), .Y(ori_ori_n294_));
  NO2        o0266(.A(ori_ori_n122_), .B(ori_ori_n294_), .Y(ori_ori_n295_));
  NA2        o0267(.A(ori_ori_n295_), .B(ori_ori_n293_), .Y(ori_ori_n296_));
  NA3        o0268(.A(ori_ori_n296_), .B(ori_ori_n288_), .C(ori_ori_n283_), .Y(ori_ori_n297_));
  NO4        o0269(.A(ori_ori_n286_), .B(ori_ori_n71_), .C(ori_ori_n63_), .D(ori_ori_n197_), .Y(ori_ori_n298_));
  NA2        o0270(.A(ori_ori_n231_), .B(ori_ori_n97_), .Y(ori_ori_n299_));
  OR2        o0271(.A(ori_ori_n299_), .B(ori_ori_n190_), .Y(ori_ori_n300_));
  NOi31      o0272(.An(l), .B(n), .C(m), .Y(ori_ori_n301_));
  NA2        o0273(.A(ori_ori_n301_), .B(ori_ori_n198_), .Y(ori_ori_n302_));
  NO2        o0274(.A(ori_ori_n302_), .B(ori_ori_n179_), .Y(ori_ori_n303_));
  NAi32      o0275(.An(ori_ori_n303_), .Bn(ori_ori_n298_), .C(ori_ori_n300_), .Y(ori_ori_n304_));
  NAi32      o0276(.An(m), .Bn(j), .C(k), .Y(ori_ori_n305_));
  NAi41      o0277(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n306_));
  OAI210     o0278(.A0(ori_ori_n194_), .A1(ori_ori_n305_), .B0(ori_ori_n306_), .Y(ori_ori_n307_));
  NOi31      o0279(.An(j), .B(m), .C(k), .Y(ori_ori_n308_));
  NO2        o0280(.A(ori_ori_n116_), .B(ori_ori_n308_), .Y(ori_ori_n309_));
  AN3        o0281(.A(h), .B(g), .C(f), .Y(ori_ori_n310_));
  NAi31      o0282(.An(ori_ori_n309_), .B(ori_ori_n310_), .C(ori_ori_n307_), .Y(ori_ori_n311_));
  NOi32      o0283(.An(m), .Bn(j), .C(l), .Y(ori_ori_n312_));
  NO2        o0284(.A(ori_ori_n312_), .B(ori_ori_n90_), .Y(ori_ori_n313_));
  NAi32      o0285(.An(ori_ori_n313_), .Bn(ori_ori_n187_), .C(ori_ori_n272_), .Y(ori_ori_n314_));
  NO2        o0286(.A(ori_ori_n268_), .B(ori_ori_n267_), .Y(ori_ori_n315_));
  NO2        o0287(.A(ori_ori_n200_), .B(g), .Y(ori_ori_n316_));
  NO2        o0288(.A(ori_ori_n146_), .B(ori_ori_n76_), .Y(ori_ori_n317_));
  AOI220     o0289(.A0(ori_ori_n317_), .A1(ori_ori_n316_), .B0(ori_ori_n228_), .B1(ori_ori_n315_), .Y(ori_ori_n318_));
  NA2        o0290(.A(ori_ori_n215_), .B(ori_ori_n71_), .Y(ori_ori_n319_));
  NA3        o0291(.A(ori_ori_n319_), .B(ori_ori_n310_), .C(ori_ori_n195_), .Y(ori_ori_n320_));
  NA4        o0292(.A(ori_ori_n320_), .B(ori_ori_n318_), .C(ori_ori_n314_), .D(ori_ori_n311_), .Y(ori_ori_n321_));
  NA3        o0293(.A(h), .B(g), .C(f), .Y(ori_ori_n322_));
  NO2        o0294(.A(ori_ori_n322_), .B(ori_ori_n67_), .Y(ori_ori_n323_));
  NA2        o0295(.A(ori_ori_n153_), .B(e), .Y(ori_ori_n324_));
  NO2        o0296(.A(ori_ori_n324_), .B(ori_ori_n40_), .Y(ori_ori_n325_));
  NOi32      o0297(.An(j), .Bn(g), .C(i), .Y(ori_ori_n326_));
  NA3        o0298(.A(ori_ori_n326_), .B(ori_ori_n263_), .C(ori_ori_n106_), .Y(ori_ori_n327_));
  OR2        o0299(.A(ori_ori_n104_), .B(ori_ori_n327_), .Y(ori_ori_n328_));
  NOi32      o0300(.An(e), .Bn(b), .C(a), .Y(ori_ori_n329_));
  AN2        o0301(.A(l), .B(j), .Y(ori_ori_n330_));
  NO2        o0302(.A(ori_ori_n284_), .B(ori_ori_n330_), .Y(ori_ori_n331_));
  NO3        o0303(.A(ori_ori_n286_), .B(ori_ori_n63_), .C(ori_ori_n197_), .Y(ori_ori_n332_));
  NA2        o0304(.A(ori_ori_n193_), .B(ori_ori_n34_), .Y(ori_ori_n333_));
  AOI220     o0305(.A0(ori_ori_n333_), .A1(ori_ori_n329_), .B0(ori_ori_n332_), .B1(ori_ori_n331_), .Y(ori_ori_n334_));
  NA4        o0306(.A(ori_ori_n189_), .B(ori_ori_n79_), .C(g), .D(ori_ori_n196_), .Y(ori_ori_n335_));
  NA2        o0307(.A(ori_ori_n50_), .B(ori_ori_n106_), .Y(ori_ori_n336_));
  NA2        o0308(.A(ori_ori_n334_), .B(ori_ori_n328_), .Y(ori_ori_n337_));
  NO4        o0309(.A(ori_ori_n337_), .B(ori_ori_n321_), .C(ori_ori_n304_), .D(ori_ori_n297_), .Y(ori_ori_n338_));
  NA4        o0310(.A(ori_ori_n338_), .B(ori_ori_n282_), .C(ori_ori_n247_), .D(ori_ori_n185_), .Y(ori10));
  NA3        o0311(.A(m), .B(k), .C(i), .Y(ori_ori_n340_));
  NOi21      o0312(.An(e), .B(f), .Y(ori_ori_n341_));
  NO4        o0313(.A(ori_ori_n141_), .B(ori_ori_n341_), .C(n), .D(ori_ori_n103_), .Y(ori_ori_n342_));
  NAi31      o0314(.An(b), .B(f), .C(c), .Y(ori_ori_n343_));
  INV        o0315(.A(ori_ori_n343_), .Y(ori_ori_n344_));
  NOi32      o0316(.An(k), .Bn(h), .C(j), .Y(ori_ori_n345_));
  NA2        o0317(.A(ori_ori_n345_), .B(ori_ori_n204_), .Y(ori_ori_n346_));
  NA2        o0318(.A(ori_ori_n151_), .B(ori_ori_n346_), .Y(ori_ori_n347_));
  NA2        o0319(.A(ori_ori_n347_), .B(ori_ori_n344_), .Y(ori_ori_n348_));
  AN2        o0320(.A(j), .B(h), .Y(ori_ori_n349_));
  NO3        o0321(.A(n), .B(m), .C(k), .Y(ori_ori_n350_));
  NA2        o0322(.A(ori_ori_n350_), .B(ori_ori_n349_), .Y(ori_ori_n351_));
  NO3        o0323(.A(ori_ori_n351_), .B(ori_ori_n141_), .C(ori_ori_n196_), .Y(ori_ori_n352_));
  OR2        o0324(.A(m), .B(k), .Y(ori_ori_n353_));
  NO2        o0325(.A(ori_ori_n159_), .B(ori_ori_n353_), .Y(ori_ori_n354_));
  NA4        o0326(.A(n), .B(f), .C(c), .D(ori_ori_n108_), .Y(ori_ori_n355_));
  NOi21      o0327(.An(ori_ori_n354_), .B(ori_ori_n355_), .Y(ori_ori_n356_));
  NOi32      o0328(.An(d), .Bn(a), .C(c), .Y(ori_ori_n357_));
  NA2        o0329(.A(ori_ori_n357_), .B(ori_ori_n167_), .Y(ori_ori_n358_));
  NO2        o0330(.A(ori_ori_n356_), .B(ori_ori_n352_), .Y(ori_ori_n359_));
  NO2        o0331(.A(ori_ori_n355_), .B(ori_ori_n268_), .Y(ori_ori_n360_));
  NOi32      o0332(.An(f), .Bn(d), .C(c), .Y(ori_ori_n361_));
  AOI220     o0333(.A0(ori_ori_n361_), .A1(ori_ori_n276_), .B0(ori_ori_n360_), .B1(ori_ori_n198_), .Y(ori_ori_n362_));
  NA3        o0334(.A(ori_ori_n362_), .B(ori_ori_n359_), .C(ori_ori_n348_), .Y(ori_ori_n363_));
  NO2        o0335(.A(ori_ori_n56_), .B(ori_ori_n108_), .Y(ori_ori_n364_));
  NA2        o0336(.A(ori_ori_n231_), .B(ori_ori_n364_), .Y(ori_ori_n365_));
  INV        o0337(.A(e), .Y(ori_ori_n366_));
  NA2        o0338(.A(ori_ori_n45_), .B(e), .Y(ori_ori_n367_));
  OAI220     o0339(.A0(ori_ori_n367_), .A1(ori_ori_n186_), .B0(ori_ori_n190_), .B1(ori_ori_n366_), .Y(ori_ori_n368_));
  NO2        o0340(.A(ori_ori_n81_), .B(ori_ori_n366_), .Y(ori_ori_n369_));
  NO2        o0341(.A(ori_ori_n93_), .B(ori_ori_n366_), .Y(ori_ori_n370_));
  NO3        o0342(.A(ori_ori_n370_), .B(ori_ori_n369_), .C(ori_ori_n368_), .Y(ori_ori_n371_));
  NOi32      o0343(.An(h), .Bn(e), .C(g), .Y(ori_ori_n372_));
  NA3        o0344(.A(ori_ori_n372_), .B(ori_ori_n265_), .C(m), .Y(ori_ori_n373_));
  NOi21      o0345(.An(g), .B(h), .Y(ori_ori_n374_));
  AN3        o0346(.A(m), .B(l), .C(i), .Y(ori_ori_n375_));
  NA3        o0347(.A(ori_ori_n375_), .B(ori_ori_n374_), .C(e), .Y(ori_ori_n376_));
  AN3        o0348(.A(h), .B(g), .C(e), .Y(ori_ori_n377_));
  NA2        o0349(.A(ori_ori_n377_), .B(ori_ori_n90_), .Y(ori_ori_n378_));
  AN3        o0350(.A(ori_ori_n378_), .B(ori_ori_n376_), .C(ori_ori_n373_), .Y(ori_ori_n379_));
  AOI210     o0351(.A0(ori_ori_n379_), .A1(ori_ori_n371_), .B0(ori_ori_n365_), .Y(ori_ori_n380_));
  NA3        o0352(.A(ori_ori_n357_), .B(ori_ori_n167_), .C(ori_ori_n76_), .Y(ori_ori_n381_));
  NAi31      o0353(.An(b), .B(c), .C(a), .Y(ori_ori_n382_));
  NO2        o0354(.A(ori_ori_n382_), .B(n), .Y(ori_ori_n383_));
  NA2        o0355(.A(ori_ori_n50_), .B(m), .Y(ori_ori_n384_));
  NO2        o0356(.A(ori_ori_n384_), .B(ori_ori_n138_), .Y(ori_ori_n385_));
  NA2        o0357(.A(ori_ori_n385_), .B(ori_ori_n383_), .Y(ori_ori_n386_));
  INV        o0358(.A(ori_ori_n386_), .Y(ori_ori_n387_));
  NO3        o0359(.A(ori_ori_n387_), .B(ori_ori_n380_), .C(ori_ori_n363_), .Y(ori_ori_n388_));
  NA2        o0360(.A(i), .B(g), .Y(ori_ori_n389_));
  NOi21      o0361(.An(a), .B(n), .Y(ori_ori_n390_));
  NOi21      o0362(.An(d), .B(c), .Y(ori_ori_n391_));
  NA2        o0363(.A(ori_ori_n391_), .B(ori_ori_n390_), .Y(ori_ori_n392_));
  NA3        o0364(.A(i), .B(g), .C(f), .Y(ori_ori_n393_));
  OR2        o0365(.A(ori_ori_n393_), .B(ori_ori_n62_), .Y(ori_ori_n394_));
  NA3        o0366(.A(ori_ori_n375_), .B(ori_ori_n374_), .C(ori_ori_n167_), .Y(ori_ori_n395_));
  AOI210     o0367(.A0(ori_ori_n395_), .A1(ori_ori_n394_), .B0(ori_ori_n392_), .Y(ori_ori_n396_));
  INV        o0368(.A(ori_ori_n396_), .Y(ori_ori_n397_));
  OR2        o0369(.A(n), .B(m), .Y(ori_ori_n398_));
  NO2        o0370(.A(ori_ori_n398_), .B(ori_ori_n142_), .Y(ori_ori_n399_));
  NO2        o0371(.A(ori_ori_n168_), .B(ori_ori_n138_), .Y(ori_ori_n400_));
  OAI210     o0372(.A0(ori_ori_n399_), .A1(ori_ori_n161_), .B0(ori_ori_n400_), .Y(ori_ori_n401_));
  INV        o0373(.A(ori_ori_n336_), .Y(ori_ori_n402_));
  NA3        o0374(.A(ori_ori_n402_), .B(ori_ori_n329_), .C(d), .Y(ori_ori_n403_));
  NO2        o0375(.A(ori_ori_n382_), .B(ori_ori_n48_), .Y(ori_ori_n404_));
  NO3        o0376(.A(ori_ori_n59_), .B(ori_ori_n105_), .C(e), .Y(ori_ori_n405_));
  NAi21      o0377(.An(k), .B(j), .Y(ori_ori_n406_));
  NA2        o0378(.A(ori_ori_n234_), .B(ori_ori_n406_), .Y(ori_ori_n407_));
  NA3        o0379(.A(ori_ori_n407_), .B(ori_ori_n405_), .C(ori_ori_n404_), .Y(ori_ori_n408_));
  NAi21      o0380(.An(e), .B(d), .Y(ori_ori_n409_));
  INV        o0381(.A(ori_ori_n409_), .Y(ori_ori_n410_));
  NO2        o0382(.A(ori_ori_n235_), .B(ori_ori_n196_), .Y(ori_ori_n411_));
  NA3        o0383(.A(ori_ori_n411_), .B(ori_ori_n410_), .C(ori_ori_n208_), .Y(ori_ori_n412_));
  NA4        o0384(.A(ori_ori_n412_), .B(ori_ori_n408_), .C(ori_ori_n403_), .D(ori_ori_n401_), .Y(ori_ori_n413_));
  NO2        o0385(.A(ori_ori_n302_), .B(ori_ori_n196_), .Y(ori_ori_n414_));
  NA2        o0386(.A(ori_ori_n414_), .B(ori_ori_n410_), .Y(ori_ori_n415_));
  NOi31      o0387(.An(n), .B(m), .C(k), .Y(ori_ori_n416_));
  AOI220     o0388(.A0(ori_ori_n416_), .A1(ori_ori_n349_), .B0(ori_ori_n204_), .B1(ori_ori_n49_), .Y(ori_ori_n417_));
  NAi31      o0389(.An(g), .B(f), .C(c), .Y(ori_ori_n418_));
  OR3        o0390(.A(ori_ori_n418_), .B(ori_ori_n417_), .C(e), .Y(ori_ori_n419_));
  NA3        o0391(.A(ori_ori_n419_), .B(ori_ori_n415_), .C(ori_ori_n277_), .Y(ori_ori_n420_));
  NOi41      o0392(.An(ori_ori_n397_), .B(ori_ori_n420_), .C(ori_ori_n413_), .D(ori_ori_n246_), .Y(ori_ori_n421_));
  NOi32      o0393(.An(c), .Bn(a), .C(b), .Y(ori_ori_n422_));
  NA2        o0394(.A(ori_ori_n422_), .B(ori_ori_n106_), .Y(ori_ori_n423_));
  NA2        o0395(.A(ori_ori_n253_), .B(ori_ori_n142_), .Y(ori_ori_n424_));
  AN2        o0396(.A(e), .B(d), .Y(ori_ori_n425_));
  NA2        o0397(.A(ori_ori_n425_), .B(ori_ori_n424_), .Y(ori_ori_n426_));
  INV        o0398(.A(ori_ori_n138_), .Y(ori_ori_n427_));
  NO2        o0399(.A(ori_ori_n121_), .B(ori_ori_n40_), .Y(ori_ori_n428_));
  NO2        o0400(.A(ori_ori_n59_), .B(e), .Y(ori_ori_n429_));
  NA2        o0401(.A(ori_ori_n154_), .B(ori_ori_n243_), .Y(ori_ori_n430_));
  AOI220     o0402(.A0(ori_ori_n430_), .A1(ori_ori_n429_), .B0(ori_ori_n428_), .B1(ori_ori_n427_), .Y(ori_ori_n431_));
  AOI210     o0403(.A0(ori_ori_n431_), .A1(ori_ori_n426_), .B0(ori_ori_n423_), .Y(ori_ori_n432_));
  INV        o0404(.A(ori_ori_n191_), .Y(ori_ori_n433_));
  NOi21      o0405(.An(a), .B(b), .Y(ori_ori_n434_));
  NA3        o0406(.A(e), .B(d), .C(c), .Y(ori_ori_n435_));
  NAi21      o0407(.An(ori_ori_n435_), .B(ori_ori_n434_), .Y(ori_ori_n436_));
  NO2        o0408(.A(ori_ori_n381_), .B(ori_ori_n190_), .Y(ori_ori_n437_));
  NOi21      o0409(.An(ori_ori_n436_), .B(ori_ori_n437_), .Y(ori_ori_n438_));
  AOI210     o0410(.A0(ori_ori_n248_), .A1(ori_ori_n433_), .B0(ori_ori_n438_), .Y(ori_ori_n439_));
  NO4        o0411(.A(ori_ori_n173_), .B(ori_ori_n96_), .C(ori_ori_n53_), .D(b), .Y(ori_ori_n440_));
  NA2        o0412(.A(ori_ori_n344_), .B(ori_ori_n143_), .Y(ori_ori_n441_));
  OR2        o0413(.A(k), .B(j), .Y(ori_ori_n442_));
  NA2        o0414(.A(l), .B(k), .Y(ori_ori_n443_));
  NA3        o0415(.A(ori_ori_n443_), .B(ori_ori_n442_), .C(ori_ori_n204_), .Y(ori_ori_n444_));
  AOI210     o0416(.A0(ori_ori_n215_), .A1(ori_ori_n305_), .B0(ori_ori_n76_), .Y(ori_ori_n445_));
  NOi21      o0417(.An(ori_ori_n444_), .B(ori_ori_n445_), .Y(ori_ori_n446_));
  OR3        o0418(.A(ori_ori_n446_), .B(ori_ori_n134_), .C(ori_ori_n125_), .Y(ori_ori_n447_));
  NA2        o0419(.A(ori_ori_n254_), .B(ori_ori_n117_), .Y(ori_ori_n448_));
  NO3        o0420(.A(ori_ori_n381_), .B(ori_ori_n84_), .C(ori_ori_n121_), .Y(ori_ori_n449_));
  NO2        o0421(.A(ori_ori_n449_), .B(ori_ori_n448_), .Y(ori_ori_n450_));
  NA3        o0422(.A(ori_ori_n450_), .B(ori_ori_n447_), .C(ori_ori_n441_), .Y(ori_ori_n451_));
  NO4        o0423(.A(ori_ori_n451_), .B(ori_ori_n440_), .C(ori_ori_n439_), .D(ori_ori_n432_), .Y(ori_ori_n452_));
  INV        o0424(.A(e), .Y(ori_ori_n453_));
  NO2        o0425(.A(ori_ori_n173_), .B(ori_ori_n53_), .Y(ori_ori_n454_));
  NAi31      o0426(.An(j), .B(l), .C(i), .Y(ori_ori_n455_));
  OAI210     o0427(.A0(ori_ori_n455_), .A1(ori_ori_n122_), .B0(ori_ori_n96_), .Y(ori_ori_n456_));
  NA3        o0428(.A(ori_ori_n456_), .B(ori_ori_n454_), .C(ori_ori_n453_), .Y(ori_ori_n457_));
  NO3        o0429(.A(ori_ori_n358_), .B(ori_ori_n313_), .C(ori_ori_n187_), .Y(ori_ori_n458_));
  NO2        o0430(.A(ori_ori_n358_), .B(ori_ori_n336_), .Y(ori_ori_n459_));
  NO4        o0431(.A(ori_ori_n459_), .B(ori_ori_n458_), .C(ori_ori_n170_), .D(ori_ori_n274_), .Y(ori_ori_n460_));
  NA3        o0432(.A(ori_ori_n460_), .B(ori_ori_n457_), .C(ori_ori_n223_), .Y(ori_ori_n461_));
  OAI210     o0433(.A0(ori_ori_n118_), .A1(ori_ori_n116_), .B0(n), .Y(ori_ori_n462_));
  NO2        o0434(.A(ori_ori_n462_), .B(ori_ori_n121_), .Y(ori_ori_n463_));
  AN2        o0435(.A(ori_ori_n463_), .B(ori_ori_n178_), .Y(ori_ori_n464_));
  XO2        o0436(.A(i), .B(h), .Y(ori_ori_n465_));
  NA3        o0437(.A(ori_ori_n465_), .B(ori_ori_n150_), .C(n), .Y(ori_ori_n466_));
  NAi41      o0438(.An(ori_ori_n269_), .B(ori_ori_n466_), .C(ori_ori_n417_), .D(ori_ori_n346_), .Y(ori_ori_n467_));
  NOi32      o0439(.An(ori_ori_n467_), .Bn(ori_ori_n429_), .C(ori_ori_n250_), .Y(ori_ori_n468_));
  NAi31      o0440(.An(c), .B(f), .C(d), .Y(ori_ori_n469_));
  AOI210     o0441(.A0(ori_ori_n255_), .A1(ori_ori_n181_), .B0(ori_ori_n469_), .Y(ori_ori_n470_));
  NOi21      o0442(.An(ori_ori_n74_), .B(ori_ori_n470_), .Y(ori_ori_n471_));
  NA2        o0443(.A(ori_ori_n209_), .B(ori_ori_n102_), .Y(ori_ori_n472_));
  AOI210     o0444(.A0(ori_ori_n472_), .A1(ori_ori_n166_), .B0(ori_ori_n469_), .Y(ori_ori_n473_));
  AOI210     o0445(.A0(ori_ori_n327_), .A1(ori_ori_n34_), .B0(ori_ori_n436_), .Y(ori_ori_n474_));
  NO2        o0446(.A(ori_ori_n474_), .B(ori_ori_n473_), .Y(ori_ori_n475_));
  AN2        o0447(.A(ori_ori_n261_), .B(ori_ori_n245_), .Y(ori_ori_n476_));
  NA3        o0448(.A(ori_ori_n36_), .B(ori_ori_n35_), .C(f), .Y(ori_ori_n477_));
  NAi31      o0449(.An(ori_ori_n476_), .B(ori_ori_n475_), .C(ori_ori_n471_), .Y(ori_ori_n478_));
  NO4        o0450(.A(ori_ori_n478_), .B(ori_ori_n468_), .C(ori_ori_n464_), .D(ori_ori_n461_), .Y(ori_ori_n479_));
  NA4        o0451(.A(ori_ori_n479_), .B(ori_ori_n452_), .C(ori_ori_n421_), .D(ori_ori_n388_), .Y(ori11));
  NO2        o0452(.A(ori_ori_n64_), .B(f), .Y(ori_ori_n481_));
  NA2        o0453(.A(j), .B(g), .Y(ori_ori_n482_));
  NAi31      o0454(.An(i), .B(m), .C(l), .Y(ori_ori_n483_));
  NA3        o0455(.A(m), .B(k), .C(j), .Y(ori_ori_n484_));
  OAI220     o0456(.A0(ori_ori_n484_), .A1(ori_ori_n121_), .B0(ori_ori_n483_), .B1(ori_ori_n482_), .Y(ori_ori_n485_));
  NA2        o0457(.A(ori_ori_n485_), .B(ori_ori_n481_), .Y(ori_ori_n486_));
  NOi32      o0458(.An(e), .Bn(b), .C(f), .Y(ori_ori_n487_));
  NA2        o0459(.A(ori_ori_n45_), .B(j), .Y(ori_ori_n488_));
  NAi31      o0460(.An(d), .B(e), .C(a), .Y(ori_ori_n489_));
  NO2        o0461(.A(ori_ori_n489_), .B(n), .Y(ori_ori_n490_));
  NA2        o0462(.A(ori_ori_n490_), .B(ori_ori_n94_), .Y(ori_ori_n491_));
  NO2        o0463(.A(ori_ori_n358_), .B(ori_ori_n251_), .Y(ori_ori_n492_));
  NA2        o0464(.A(j), .B(i), .Y(ori_ori_n493_));
  NAi31      o0465(.An(n), .B(m), .C(k), .Y(ori_ori_n494_));
  NO3        o0466(.A(ori_ori_n494_), .B(ori_ori_n493_), .C(ori_ori_n105_), .Y(ori_ori_n495_));
  NO4        o0467(.A(n), .B(d), .C(ori_ori_n108_), .D(a), .Y(ori_ori_n496_));
  INV        o0468(.A(ori_ori_n496_), .Y(ori_ori_n497_));
  NA2        o0469(.A(ori_ori_n485_), .B(f), .Y(ori_ori_n498_));
  NO2        o0470(.A(ori_ori_n253_), .B(ori_ori_n48_), .Y(ori_ori_n499_));
  NO2        o0471(.A(ori_ori_n498_), .B(ori_ori_n497_), .Y(ori_ori_n500_));
  AOI210     o0472(.A0(ori_ori_n495_), .A1(ori_ori_n492_), .B0(ori_ori_n500_), .Y(ori_ori_n501_));
  NA2        o0473(.A(ori_ori_n130_), .B(ori_ori_n33_), .Y(ori_ori_n502_));
  OAI220     o0474(.A0(ori_ori_n502_), .A1(m), .B0(ori_ori_n488_), .B1(ori_ori_n215_), .Y(ori_ori_n503_));
  NOi41      o0475(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n504_));
  NAi32      o0476(.An(e), .Bn(b), .C(c), .Y(ori_ori_n505_));
  OR2        o0477(.A(ori_ori_n505_), .B(ori_ori_n76_), .Y(ori_ori_n506_));
  AN2        o0478(.A(ori_ori_n306_), .B(ori_ori_n286_), .Y(ori_ori_n507_));
  NA2        o0479(.A(ori_ori_n507_), .B(ori_ori_n506_), .Y(ori_ori_n508_));
  OA210      o0480(.A0(ori_ori_n508_), .A1(ori_ori_n504_), .B0(ori_ori_n503_), .Y(ori_ori_n509_));
  NO2        o0481(.A(ori_ori_n483_), .B(ori_ori_n482_), .Y(ori_ori_n510_));
  INV        o0482(.A(ori_ori_n383_), .Y(ori_ori_n511_));
  NA2        o0483(.A(ori_ori_n510_), .B(f), .Y(ori_ori_n512_));
  NAi32      o0484(.An(d), .Bn(a), .C(b), .Y(ori_ori_n513_));
  NO2        o0485(.A(ori_ori_n513_), .B(ori_ori_n48_), .Y(ori_ori_n514_));
  NA2        o0486(.A(h), .B(f), .Y(ori_ori_n515_));
  NO2        o0487(.A(ori_ori_n515_), .B(ori_ori_n87_), .Y(ori_ori_n516_));
  NO3        o0488(.A(ori_ori_n162_), .B(ori_ori_n159_), .C(g), .Y(ori_ori_n517_));
  AOI220     o0489(.A0(ori_ori_n517_), .A1(ori_ori_n55_), .B0(ori_ori_n516_), .B1(ori_ori_n514_), .Y(ori_ori_n518_));
  OAI210     o0490(.A0(ori_ori_n512_), .A1(ori_ori_n511_), .B0(ori_ori_n518_), .Y(ori_ori_n519_));
  AN3        o0491(.A(j), .B(h), .C(g), .Y(ori_ori_n520_));
  NO2        o0492(.A(ori_ori_n137_), .B(c), .Y(ori_ori_n521_));
  NA3        o0493(.A(ori_ori_n521_), .B(ori_ori_n520_), .C(ori_ori_n416_), .Y(ori_ori_n522_));
  NA3        o0494(.A(f), .B(d), .C(b), .Y(ori_ori_n523_));
  NO4        o0495(.A(ori_ori_n523_), .B(ori_ori_n162_), .C(ori_ori_n159_), .D(g), .Y(ori_ori_n524_));
  NAi21      o0496(.An(ori_ori_n524_), .B(ori_ori_n522_), .Y(ori_ori_n525_));
  NO3        o0497(.A(ori_ori_n525_), .B(ori_ori_n519_), .C(ori_ori_n509_), .Y(ori_ori_n526_));
  AN4        o0498(.A(ori_ori_n526_), .B(ori_ori_n501_), .C(ori_ori_n491_), .D(ori_ori_n486_), .Y(ori_ori_n527_));
  INV        o0499(.A(k), .Y(ori_ori_n528_));
  NA3        o0500(.A(l), .B(ori_ori_n528_), .C(i), .Y(ori_ori_n529_));
  INV        o0501(.A(ori_ori_n529_), .Y(ori_ori_n530_));
  NA4        o0502(.A(ori_ori_n357_), .B(ori_ori_n374_), .C(ori_ori_n167_), .D(ori_ori_n106_), .Y(ori_ori_n531_));
  NAi32      o0503(.An(h), .Bn(f), .C(g), .Y(ori_ori_n532_));
  NAi41      o0504(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n533_));
  OAI210     o0505(.A0(ori_ori_n489_), .A1(n), .B0(ori_ori_n533_), .Y(ori_ori_n534_));
  NA2        o0506(.A(ori_ori_n534_), .B(m), .Y(ori_ori_n535_));
  NAi31      o0507(.An(h), .B(g), .C(f), .Y(ori_ori_n536_));
  OR2        o0508(.A(ori_ori_n535_), .B(ori_ori_n532_), .Y(ori_ori_n537_));
  NO3        o0509(.A(ori_ori_n532_), .B(ori_ori_n64_), .C(ori_ori_n65_), .Y(ori_ori_n538_));
  NAi31      o0510(.An(ori_ori_n538_), .B(ori_ori_n537_), .C(ori_ori_n531_), .Y(ori_ori_n539_));
  NAi31      o0511(.An(f), .B(h), .C(g), .Y(ori_ori_n540_));
  NOi32      o0512(.An(d), .Bn(a), .C(e), .Y(ori_ori_n541_));
  NOi32      o0513(.An(e), .Bn(a), .C(d), .Y(ori_ori_n542_));
  AOI210     o0514(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n542_), .Y(ori_ori_n543_));
  NO2        o0515(.A(ori_ori_n230_), .B(ori_ori_n79_), .Y(ori_ori_n544_));
  AOI210     o0516(.A0(ori_ori_n539_), .A1(ori_ori_n530_), .B0(ori_ori_n544_), .Y(ori_ori_n545_));
  NO3        o0517(.A(ori_ori_n284_), .B(ori_ori_n57_), .C(n), .Y(ori_ori_n546_));
  NA3        o0518(.A(ori_ori_n469_), .B(ori_ori_n157_), .C(ori_ori_n156_), .Y(ori_ori_n547_));
  NA2        o0519(.A(ori_ori_n418_), .B(ori_ori_n212_), .Y(ori_ori_n548_));
  OR2        o0520(.A(ori_ori_n548_), .B(ori_ori_n547_), .Y(ori_ori_n549_));
  NA2        o0521(.A(ori_ori_n66_), .B(ori_ori_n106_), .Y(ori_ori_n550_));
  NA2        o0522(.A(ori_ori_n549_), .B(ori_ori_n546_), .Y(ori_ori_n551_));
  NO2        o0523(.A(ori_ori_n551_), .B(ori_ori_n79_), .Y(ori_ori_n552_));
  NA3        o0524(.A(ori_ori_n504_), .B(ori_ori_n308_), .C(ori_ori_n45_), .Y(ori_ori_n553_));
  NOi32      o0525(.An(e), .Bn(c), .C(f), .Y(ori_ori_n554_));
  NOi21      o0526(.An(f), .B(g), .Y(ori_ori_n555_));
  NO2        o0527(.A(ori_ori_n555_), .B(ori_ori_n194_), .Y(ori_ori_n556_));
  AOI220     o0528(.A0(ori_ori_n556_), .A1(ori_ori_n354_), .B0(ori_ori_n554_), .B1(ori_ori_n161_), .Y(ori_ori_n557_));
  NA3        o0529(.A(ori_ori_n557_), .B(ori_ori_n553_), .C(ori_ori_n164_), .Y(ori_ori_n558_));
  NOi21      o0530(.An(j), .B(l), .Y(ori_ori_n559_));
  NAi21      o0531(.An(k), .B(h), .Y(ori_ori_n560_));
  NO2        o0532(.A(ori_ori_n560_), .B(ori_ori_n244_), .Y(ori_ori_n561_));
  NA2        o0533(.A(ori_ori_n561_), .B(ori_ori_n559_), .Y(ori_ori_n562_));
  OR2        o0534(.A(ori_ori_n562_), .B(ori_ori_n535_), .Y(ori_ori_n563_));
  NO2        o0535(.A(ori_ori_n278_), .B(ori_ori_n540_), .Y(ori_ori_n564_));
  NO2        o0536(.A(ori_ori_n489_), .B(ori_ori_n48_), .Y(ori_ori_n565_));
  NA2        o0537(.A(ori_ori_n565_), .B(ori_ori_n564_), .Y(ori_ori_n566_));
  NA2        o0538(.A(ori_ori_n566_), .B(ori_ori_n563_), .Y(ori_ori_n567_));
  NA2        o0539(.A(ori_ori_n102_), .B(ori_ori_n35_), .Y(ori_ori_n568_));
  NO2        o0540(.A(k), .B(ori_ori_n197_), .Y(ori_ori_n569_));
  INV        o0541(.A(ori_ori_n329_), .Y(ori_ori_n570_));
  NO2        o0542(.A(ori_ori_n570_), .B(n), .Y(ori_ori_n571_));
  NAi31      o0543(.An(ori_ori_n568_), .B(ori_ori_n571_), .C(ori_ori_n569_), .Y(ori_ori_n572_));
  NO2        o0544(.A(ori_ori_n488_), .B(ori_ori_n162_), .Y(ori_ori_n573_));
  NA3        o0545(.A(ori_ori_n505_), .B(ori_ori_n250_), .C(ori_ori_n135_), .Y(ori_ori_n574_));
  NA2        o0546(.A(ori_ori_n465_), .B(ori_ori_n150_), .Y(ori_ori_n575_));
  NO3        o0547(.A(ori_ori_n355_), .B(ori_ori_n575_), .C(ori_ori_n79_), .Y(ori_ori_n576_));
  AOI210     o0548(.A0(ori_ori_n574_), .A1(ori_ori_n573_), .B0(ori_ori_n576_), .Y(ori_ori_n577_));
  AN3        o0549(.A(f), .B(d), .C(b), .Y(ori_ori_n578_));
  OAI210     o0550(.A0(ori_ori_n578_), .A1(ori_ori_n120_), .B0(n), .Y(ori_ori_n579_));
  NA3        o0551(.A(ori_ori_n465_), .B(ori_ori_n150_), .C(ori_ori_n197_), .Y(ori_ori_n580_));
  AOI210     o0552(.A0(ori_ori_n579_), .A1(ori_ori_n214_), .B0(ori_ori_n580_), .Y(ori_ori_n581_));
  NAi31      o0553(.An(m), .B(n), .C(k), .Y(ori_ori_n582_));
  OR2        o0554(.A(ori_ori_n125_), .B(ori_ori_n57_), .Y(ori_ori_n583_));
  OAI210     o0555(.A0(ori_ori_n583_), .A1(ori_ori_n582_), .B0(ori_ori_n232_), .Y(ori_ori_n584_));
  OAI210     o0556(.A0(ori_ori_n584_), .A1(ori_ori_n581_), .B0(j), .Y(ori_ori_n585_));
  NA3        o0557(.A(ori_ori_n585_), .B(ori_ori_n577_), .C(ori_ori_n572_), .Y(ori_ori_n586_));
  NO4        o0558(.A(ori_ori_n586_), .B(ori_ori_n567_), .C(ori_ori_n558_), .D(ori_ori_n552_), .Y(ori_ori_n587_));
  NA2        o0559(.A(ori_ori_n342_), .B(ori_ori_n153_), .Y(ori_ori_n588_));
  NAi31      o0560(.An(g), .B(h), .C(f), .Y(ori_ori_n589_));
  OA210      o0561(.A0(ori_ori_n489_), .A1(n), .B0(ori_ori_n533_), .Y(ori_ori_n590_));
  NO2        o0562(.A(ori_ori_n590_), .B(ori_ori_n83_), .Y(ori_ori_n591_));
  INV        o0563(.A(ori_ori_n591_), .Y(ori_ori_n592_));
  AOI210     o0564(.A0(ori_ori_n592_), .A1(ori_ori_n588_), .B0(ori_ori_n484_), .Y(ori_ori_n593_));
  NO3        o0565(.A(g), .B(ori_ori_n196_), .C(ori_ori_n53_), .Y(ori_ori_n594_));
  NAi21      o0566(.An(h), .B(j), .Y(ori_ori_n595_));
  NO2        o0567(.A(ori_ori_n472_), .B(ori_ori_n79_), .Y(ori_ori_n596_));
  OAI210     o0568(.A0(ori_ori_n596_), .A1(ori_ori_n354_), .B0(ori_ori_n594_), .Y(ori_ori_n597_));
  OR2        o0569(.A(ori_ori_n64_), .B(ori_ori_n65_), .Y(ori_ori_n598_));
  OR2        o0570(.A(ori_ori_n562_), .B(ori_ori_n598_), .Y(ori_ori_n599_));
  AN2        o0571(.A(h), .B(f), .Y(ori_ori_n600_));
  NA2        o0572(.A(ori_ori_n600_), .B(ori_ori_n36_), .Y(ori_ori_n601_));
  NA2        o0573(.A(ori_ori_n92_), .B(ori_ori_n45_), .Y(ori_ori_n602_));
  OAI220     o0574(.A0(ori_ori_n602_), .A1(ori_ori_n299_), .B0(ori_ori_n601_), .B1(ori_ori_n423_), .Y(ori_ori_n603_));
  AOI210     o0575(.A0(ori_ori_n513_), .A1(ori_ori_n382_), .B0(ori_ori_n48_), .Y(ori_ori_n604_));
  OAI220     o0576(.A0(ori_ori_n536_), .A1(ori_ori_n529_), .B0(ori_ori_n292_), .B1(ori_ori_n482_), .Y(ori_ori_n605_));
  AOI210     o0577(.A0(ori_ori_n605_), .A1(ori_ori_n604_), .B0(ori_ori_n603_), .Y(ori_ori_n606_));
  NA3        o0578(.A(ori_ori_n606_), .B(ori_ori_n599_), .C(ori_ori_n597_), .Y(ori_ori_n607_));
  NO2        o0579(.A(ori_ori_n555_), .B(ori_ori_n57_), .Y(ori_ori_n608_));
  NO2        o0580(.A(ori_ori_n608_), .B(ori_ori_n33_), .Y(ori_ori_n609_));
  NA2        o0581(.A(ori_ori_n295_), .B(ori_ori_n130_), .Y(ori_ori_n610_));
  NA2        o0582(.A(ori_ori_n122_), .B(ori_ori_n48_), .Y(ori_ori_n611_));
  AOI220     o0583(.A0(ori_ori_n611_), .A1(ori_ori_n487_), .B0(ori_ori_n329_), .B1(ori_ori_n106_), .Y(ori_ori_n612_));
  OA220      o0584(.A0(ori_ori_n612_), .A1(ori_ori_n502_), .B0(ori_ori_n327_), .B1(ori_ori_n104_), .Y(ori_ori_n613_));
  OAI210     o0585(.A0(ori_ori_n610_), .A1(ori_ori_n609_), .B0(ori_ori_n613_), .Y(ori_ori_n614_));
  NO3        o0586(.A(ori_ori_n361_), .B(ori_ori_n178_), .C(ori_ori_n177_), .Y(ori_ori_n615_));
  NA2        o0587(.A(ori_ori_n615_), .B(ori_ori_n212_), .Y(ori_ori_n616_));
  NA3        o0588(.A(ori_ori_n616_), .B(ori_ori_n236_), .C(j), .Y(ori_ori_n617_));
  NO3        o0589(.A(ori_ori_n418_), .B(ori_ori_n159_), .C(i), .Y(ori_ori_n618_));
  NA2        o0590(.A(ori_ori_n422_), .B(ori_ori_n76_), .Y(ori_ori_n619_));
  NO4        o0591(.A(ori_ori_n484_), .B(ori_ori_n619_), .C(ori_ori_n121_), .D(ori_ori_n196_), .Y(ori_ori_n620_));
  INV        o0592(.A(ori_ori_n620_), .Y(ori_ori_n621_));
  NA3        o0593(.A(ori_ori_n621_), .B(ori_ori_n617_), .C(ori_ori_n359_), .Y(ori_ori_n622_));
  NO4        o0594(.A(ori_ori_n622_), .B(ori_ori_n614_), .C(ori_ori_n607_), .D(ori_ori_n593_), .Y(ori_ori_n623_));
  NA4        o0595(.A(ori_ori_n623_), .B(ori_ori_n587_), .C(ori_ori_n545_), .D(ori_ori_n527_), .Y(ori08));
  NO2        o0596(.A(k), .B(h), .Y(ori_ori_n625_));
  AO210      o0597(.A0(ori_ori_n234_), .A1(ori_ori_n406_), .B0(ori_ori_n625_), .Y(ori_ori_n626_));
  NO2        o0598(.A(ori_ori_n626_), .B(ori_ori_n268_), .Y(ori_ori_n627_));
  NA2        o0599(.A(ori_ori_n554_), .B(ori_ori_n76_), .Y(ori_ori_n628_));
  NA2        o0600(.A(ori_ori_n628_), .B(ori_ori_n418_), .Y(ori_ori_n629_));
  AOI210     o0601(.A0(ori_ori_n629_), .A1(ori_ori_n627_), .B0(ori_ori_n449_), .Y(ori_ori_n630_));
  NA2        o0602(.A(ori_ori_n76_), .B(ori_ori_n103_), .Y(ori_ori_n631_));
  NO2        o0603(.A(ori_ori_n631_), .B(ori_ori_n54_), .Y(ori_ori_n632_));
  NO4        o0604(.A(ori_ori_n340_), .B(ori_ori_n105_), .C(j), .D(ori_ori_n197_), .Y(ori_ori_n633_));
  NA2        o0605(.A(ori_ori_n523_), .B(ori_ori_n214_), .Y(ori_ori_n634_));
  AOI220     o0606(.A0(ori_ori_n634_), .A1(ori_ori_n316_), .B0(ori_ori_n633_), .B1(ori_ori_n632_), .Y(ori_ori_n635_));
  AOI210     o0607(.A0(ori_ori_n523_), .A1(ori_ori_n146_), .B0(ori_ori_n76_), .Y(ori_ori_n636_));
  NA4        o0608(.A(ori_ori_n199_), .B(ori_ori_n130_), .C(ori_ori_n44_), .D(h), .Y(ori_ori_n637_));
  AN2        o0609(.A(l), .B(k), .Y(ori_ori_n638_));
  NA4        o0610(.A(ori_ori_n638_), .B(ori_ori_n102_), .C(ori_ori_n65_), .D(ori_ori_n197_), .Y(ori_ori_n639_));
  OAI210     o0611(.A0(ori_ori_n637_), .A1(g), .B0(ori_ori_n639_), .Y(ori_ori_n640_));
  NA2        o0612(.A(ori_ori_n640_), .B(ori_ori_n636_), .Y(ori_ori_n641_));
  NA4        o0613(.A(ori_ori_n641_), .B(ori_ori_n635_), .C(ori_ori_n630_), .D(ori_ori_n318_), .Y(ori_ori_n642_));
  AN2        o0614(.A(ori_ori_n490_), .B(ori_ori_n88_), .Y(ori_ori_n643_));
  NO4        o0615(.A(ori_ori_n159_), .B(ori_ori_n353_), .C(ori_ori_n105_), .D(g), .Y(ori_ori_n644_));
  NA2        o0616(.A(ori_ori_n644_), .B(ori_ori_n634_), .Y(ori_ori_n645_));
  NO2        o0617(.A(ori_ori_n37_), .B(ori_ori_n196_), .Y(ori_ori_n646_));
  NA2        o0618(.A(ori_ori_n556_), .B(ori_ori_n315_), .Y(ori_ori_n647_));
  NAi31      o0619(.An(ori_ori_n643_), .B(ori_ori_n647_), .C(ori_ori_n645_), .Y(ori_ori_n648_));
  OAI210     o0620(.A0(ori_ori_n505_), .A1(ori_ori_n46_), .B0(ori_ori_n583_), .Y(ori_ori_n649_));
  NO2        o0621(.A(ori_ori_n443_), .B(ori_ori_n122_), .Y(ori_ori_n650_));
  NA2        o0622(.A(ori_ori_n650_), .B(ori_ori_n649_), .Y(ori_ori_n651_));
  NO3        o0623(.A(ori_ori_n284_), .B(ori_ori_n121_), .C(ori_ori_n40_), .Y(ori_ori_n652_));
  NAi21      o0624(.An(ori_ori_n652_), .B(ori_ori_n639_), .Y(ori_ori_n653_));
  NA2        o0625(.A(ori_ori_n626_), .B(ori_ori_n126_), .Y(ori_ori_n654_));
  AOI220     o0626(.A0(ori_ori_n654_), .A1(ori_ori_n360_), .B0(ori_ori_n653_), .B1(ori_ori_n68_), .Y(ori_ori_n655_));
  NA2        o0627(.A(ori_ori_n651_), .B(ori_ori_n655_), .Y(ori_ori_n656_));
  NA2        o0628(.A(ori_ori_n329_), .B(ori_ori_n42_), .Y(ori_ori_n657_));
  NA3        o0629(.A(ori_ori_n616_), .B(ori_ori_n301_), .C(ori_ori_n345_), .Y(ori_ori_n658_));
  NA3        o0630(.A(m), .B(l), .C(k), .Y(ori_ori_n659_));
  NA4        o0631(.A(ori_ori_n106_), .B(l), .C(k), .D(ori_ori_n79_), .Y(ori_ori_n660_));
  NA2        o0632(.A(ori_ori_n658_), .B(ori_ori_n657_), .Y(ori_ori_n661_));
  NO4        o0633(.A(ori_ori_n661_), .B(ori_ori_n656_), .C(ori_ori_n648_), .D(ori_ori_n642_), .Y(ori_ori_n662_));
  NA2        o0634(.A(ori_ori_n556_), .B(ori_ori_n354_), .Y(ori_ori_n663_));
  NO3        o0635(.A(ori_ori_n358_), .B(ori_ori_n482_), .C(h), .Y(ori_ori_n664_));
  AOI210     o0636(.A0(ori_ori_n664_), .A1(ori_ori_n106_), .B0(ori_ori_n459_), .Y(ori_ori_n665_));
  NA3        o0637(.A(ori_ori_n665_), .B(ori_ori_n663_), .C(ori_ori_n233_), .Y(ori_ori_n666_));
  NA2        o0638(.A(ori_ori_n638_), .B(ori_ori_n65_), .Y(ori_ori_n667_));
  NO4        o0639(.A(ori_ori_n615_), .B(ori_ori_n159_), .C(n), .D(i), .Y(ori_ori_n668_));
  NOi21      o0640(.An(h), .B(j), .Y(ori_ori_n669_));
  NA2        o0641(.A(ori_ori_n669_), .B(f), .Y(ori_ori_n670_));
  NO2        o0642(.A(ori_ori_n668_), .B(ori_ori_n618_), .Y(ori_ori_n671_));
  NO2        o0643(.A(ori_ori_n671_), .B(ori_ori_n667_), .Y(ori_ori_n672_));
  AOI210     o0644(.A0(ori_ori_n666_), .A1(l), .B0(ori_ori_n672_), .Y(ori_ori_n673_));
  NO2        o0645(.A(j), .B(i), .Y(ori_ori_n674_));
  NA3        o0646(.A(ori_ori_n674_), .B(ori_ori_n72_), .C(l), .Y(ori_ori_n675_));
  NA2        o0647(.A(ori_ori_n674_), .B(ori_ori_n32_), .Y(ori_ori_n676_));
  OR2        o0648(.A(ori_ori_n675_), .B(ori_ori_n535_), .Y(ori_ori_n677_));
  NO3        o0649(.A(ori_ori_n141_), .B(ori_ori_n48_), .C(ori_ori_n103_), .Y(ori_ori_n678_));
  NO3        o0650(.A(ori_ori_n443_), .B(ori_ori_n393_), .C(j), .Y(ori_ori_n679_));
  NA2        o0651(.A(k), .B(j), .Y(ori_ori_n680_));
  NO3        o0652(.A(ori_ori_n268_), .B(ori_ori_n680_), .C(ori_ori_n39_), .Y(ori_ori_n681_));
  AOI210     o0653(.A0(ori_ori_n487_), .A1(n), .B0(ori_ori_n504_), .Y(ori_ori_n682_));
  NA2        o0654(.A(ori_ori_n682_), .B(ori_ori_n507_), .Y(ori_ori_n683_));
  AN3        o0655(.A(ori_ori_n683_), .B(ori_ori_n681_), .C(ori_ori_n91_), .Y(ori_ori_n684_));
  NA2        o0656(.A(ori_ori_n548_), .B(ori_ori_n276_), .Y(ori_ori_n685_));
  NAi31      o0657(.An(ori_ori_n543_), .B(ori_ori_n85_), .C(ori_ori_n76_), .Y(ori_ori_n686_));
  NA2        o0658(.A(ori_ori_n686_), .B(ori_ori_n685_), .Y(ori_ori_n687_));
  NO2        o0659(.A(ori_ori_n268_), .B(ori_ori_n126_), .Y(ori_ori_n688_));
  AOI220     o0660(.A0(ori_ori_n688_), .A1(ori_ori_n556_), .B0(ori_ori_n652_), .B1(ori_ori_n636_), .Y(ori_ori_n689_));
  NO2        o0661(.A(ori_ori_n659_), .B(ori_ori_n83_), .Y(ori_ori_n690_));
  NA2        o0662(.A(ori_ori_n690_), .B(ori_ori_n534_), .Y(ori_ori_n691_));
  NO2        o0663(.A(ori_ori_n536_), .B(ori_ori_n109_), .Y(ori_ori_n692_));
  OAI210     o0664(.A0(ori_ori_n692_), .A1(ori_ori_n679_), .B0(ori_ori_n604_), .Y(ori_ori_n693_));
  NA3        o0665(.A(ori_ori_n693_), .B(ori_ori_n691_), .C(ori_ori_n689_), .Y(ori_ori_n694_));
  OR3        o0666(.A(ori_ori_n694_), .B(ori_ori_n687_), .C(ori_ori_n684_), .Y(ori_ori_n695_));
  NA3        o0667(.A(ori_ori_n682_), .B(ori_ori_n507_), .C(ori_ori_n506_), .Y(ori_ori_n696_));
  NA4        o0668(.A(ori_ori_n696_), .B(ori_ori_n199_), .C(ori_ori_n406_), .D(ori_ori_n33_), .Y(ori_ori_n697_));
  NO4        o0669(.A(ori_ori_n443_), .B(ori_ori_n389_), .C(j), .D(f), .Y(ori_ori_n698_));
  OAI220     o0670(.A0(ori_ori_n637_), .A1(ori_ori_n628_), .B0(ori_ori_n299_), .B1(ori_ori_n37_), .Y(ori_ori_n699_));
  AOI210     o0671(.A0(ori_ori_n698_), .A1(ori_ori_n240_), .B0(ori_ori_n699_), .Y(ori_ori_n700_));
  NO2        o0672(.A(ori_ori_n84_), .B(ori_ori_n46_), .Y(ori_ori_n701_));
  NA2        o0673(.A(ori_ori_n701_), .B(ori_ori_n571_), .Y(ori_ori_n702_));
  NA3        o0674(.A(ori_ori_n702_), .B(ori_ori_n700_), .C(ori_ori_n697_), .Y(ori_ori_n703_));
  BUFFER     o0675(.A(ori_ori_n690_), .Y(ori_ori_n704_));
  NA2        o0676(.A(ori_ori_n704_), .B(ori_ori_n219_), .Y(ori_ori_n705_));
  NO2        o0677(.A(ori_ori_n590_), .B(ori_ori_n65_), .Y(ori_ori_n706_));
  AOI210     o0678(.A0(ori_ori_n698_), .A1(ori_ori_n706_), .B0(ori_ori_n303_), .Y(ori_ori_n707_));
  OAI210     o0679(.A0(ori_ori_n659_), .A1(ori_ori_n589_), .B0(ori_ori_n477_), .Y(ori_ori_n708_));
  NA3        o0680(.A(ori_ori_n231_), .B(ori_ori_n56_), .C(b), .Y(ori_ori_n709_));
  NA2        o0681(.A(ori_ori_n422_), .B(ori_ori_n76_), .Y(ori_ori_n710_));
  NA2        o0682(.A(ori_ori_n710_), .B(ori_ori_n709_), .Y(ori_ori_n711_));
  NA2        o0683(.A(ori_ori_n711_), .B(ori_ori_n708_), .Y(ori_ori_n712_));
  NA3        o0684(.A(ori_ori_n712_), .B(ori_ori_n707_), .C(ori_ori_n705_), .Y(ori_ori_n713_));
  NOi41      o0685(.An(ori_ori_n677_), .B(ori_ori_n713_), .C(ori_ori_n703_), .D(ori_ori_n695_), .Y(ori_ori_n714_));
  NO3        o0686(.A(ori_ori_n309_), .B(ori_ori_n270_), .C(ori_ori_n105_), .Y(ori_ori_n715_));
  NA2        o0687(.A(ori_ori_n715_), .B(ori_ori_n683_), .Y(ori_ori_n716_));
  NO3        o0688(.A(ori_ori_n482_), .B(ori_ori_n86_), .C(h), .Y(ori_ori_n717_));
  NA2        o0689(.A(ori_ori_n717_), .B(ori_ori_n632_), .Y(ori_ori_n718_));
  NA3        o0690(.A(ori_ori_n718_), .B(ori_ori_n716_), .C(ori_ori_n362_), .Y(ori_ori_n719_));
  OR2        o0691(.A(ori_ori_n589_), .B(ori_ori_n84_), .Y(ori_ori_n720_));
  NOi31      o0692(.An(b), .B(d), .C(a), .Y(ori_ori_n721_));
  NO2        o0693(.A(ori_ori_n721_), .B(ori_ori_n541_), .Y(ori_ori_n722_));
  NO2        o0694(.A(ori_ori_n722_), .B(n), .Y(ori_ori_n723_));
  NOi21      o0695(.An(ori_ori_n710_), .B(ori_ori_n723_), .Y(ori_ori_n724_));
  NO2        o0696(.A(ori_ori_n724_), .B(ori_ori_n720_), .Y(ori_ori_n725_));
  NO2        o0697(.A(ori_ori_n505_), .B(ori_ori_n76_), .Y(ori_ori_n726_));
  NA2        o0698(.A(ori_ori_n715_), .B(ori_ori_n726_), .Y(ori_ori_n727_));
  OAI210     o0699(.A0(ori_ori_n637_), .A1(ori_ori_n355_), .B0(ori_ori_n727_), .Y(ori_ori_n728_));
  NO2        o0700(.A(ori_ori_n615_), .B(n), .Y(ori_ori_n729_));
  AOI220     o0701(.A0(ori_ori_n688_), .A1(ori_ori_n594_), .B0(ori_ori_n729_), .B1(ori_ori_n627_), .Y(ori_ori_n730_));
  NO2        o0702(.A(ori_ori_n289_), .B(ori_ori_n218_), .Y(ori_ori_n731_));
  OAI210     o0703(.A0(ori_ori_n88_), .A1(ori_ori_n85_), .B0(ori_ori_n731_), .Y(ori_ori_n732_));
  INV        o0704(.A(ori_ori_n732_), .Y(ori_ori_n733_));
  NA2        o0705(.A(ori_ori_n644_), .B(ori_ori_n317_), .Y(ori_ori_n734_));
  NA2        o0706(.A(ori_ori_n538_), .B(ori_ori_n330_), .Y(ori_ori_n735_));
  AN2        o0707(.A(ori_ori_n735_), .B(ori_ori_n734_), .Y(ori_ori_n736_));
  NAi31      o0708(.An(ori_ori_n733_), .B(ori_ori_n736_), .C(ori_ori_n730_), .Y(ori_ori_n737_));
  NO4        o0709(.A(ori_ori_n737_), .B(ori_ori_n728_), .C(ori_ori_n725_), .D(ori_ori_n719_), .Y(ori_ori_n738_));
  NA4        o0710(.A(ori_ori_n738_), .B(ori_ori_n714_), .C(ori_ori_n673_), .D(ori_ori_n662_), .Y(ori09));
  INV        o0711(.A(ori_ori_n113_), .Y(ori_ori_n740_));
  NA2        o0712(.A(f), .B(e), .Y(ori_ori_n741_));
  NO2        o0713(.A(ori_ori_n207_), .B(ori_ori_n105_), .Y(ori_ori_n742_));
  NA2        o0714(.A(ori_ori_n742_), .B(g), .Y(ori_ori_n743_));
  NA3        o0715(.A(ori_ori_n278_), .B(ori_ori_n154_), .C(ori_ori_n243_), .Y(ori_ori_n744_));
  AOI210     o0716(.A0(ori_ori_n744_), .A1(g), .B0(ori_ori_n428_), .Y(ori_ori_n745_));
  AOI210     o0717(.A0(ori_ori_n745_), .A1(ori_ori_n743_), .B0(ori_ori_n741_), .Y(ori_ori_n746_));
  NA2        o0718(.A(ori_ori_n399_), .B(e), .Y(ori_ori_n747_));
  NO2        o0719(.A(ori_ori_n747_), .B(ori_ori_n469_), .Y(ori_ori_n748_));
  AOI210     o0720(.A0(ori_ori_n746_), .A1(ori_ori_n740_), .B0(ori_ori_n748_), .Y(ori_ori_n749_));
  NA3        o0721(.A(m), .B(l), .C(i), .Y(ori_ori_n750_));
  OAI220     o0722(.A0(ori_ori_n536_), .A1(ori_ori_n750_), .B0(ori_ori_n322_), .B1(ori_ori_n483_), .Y(ori_ori_n751_));
  NAi21      o0723(.An(ori_ori_n751_), .B(ori_ori_n394_), .Y(ori_ori_n752_));
  NA3        o0724(.A(ori_ori_n720_), .B(ori_ori_n512_), .C(ori_ori_n477_), .Y(ori_ori_n753_));
  OA210      o0725(.A0(ori_ori_n753_), .A1(ori_ori_n752_), .B0(ori_ori_n723_), .Y(ori_ori_n754_));
  INV        o0726(.A(ori_ori_n306_), .Y(ori_ori_n755_));
  NO2        o0727(.A(ori_ori_n118_), .B(ori_ori_n116_), .Y(ori_ori_n756_));
  NOi31      o0728(.An(k), .B(m), .C(l), .Y(ori_ori_n757_));
  NO2        o0729(.A(ori_ori_n308_), .B(ori_ori_n757_), .Y(ori_ori_n758_));
  AOI210     o0730(.A0(ori_ori_n758_), .A1(ori_ori_n756_), .B0(ori_ori_n540_), .Y(ori_ori_n759_));
  NA2        o0731(.A(ori_ori_n709_), .B(ori_ori_n299_), .Y(ori_ori_n760_));
  NA2        o0732(.A(ori_ori_n310_), .B(ori_ori_n312_), .Y(ori_ori_n761_));
  OAI210     o0733(.A0(ori_ori_n190_), .A1(ori_ori_n196_), .B0(ori_ori_n761_), .Y(ori_ori_n762_));
  AOI220     o0734(.A0(ori_ori_n762_), .A1(ori_ori_n760_), .B0(ori_ori_n759_), .B1(ori_ori_n755_), .Y(ori_ori_n763_));
  NA2        o0735(.A(ori_ori_n626_), .B(ori_ori_n126_), .Y(ori_ori_n764_));
  NA3        o0736(.A(ori_ori_n764_), .B(ori_ori_n175_), .C(ori_ori_n31_), .Y(ori_ori_n765_));
  NA4        o0737(.A(ori_ori_n765_), .B(ori_ori_n763_), .C(ori_ori_n557_), .D(ori_ori_n74_), .Y(ori_ori_n766_));
  NO2        o0738(.A(ori_ori_n532_), .B(ori_ori_n455_), .Y(ori_ori_n767_));
  NA2        o0739(.A(ori_ori_n767_), .B(ori_ori_n175_), .Y(ori_ori_n768_));
  NOi21      o0740(.An(f), .B(d), .Y(ori_ori_n769_));
  NA2        o0741(.A(ori_ori_n769_), .B(m), .Y(ori_ori_n770_));
  NO2        o0742(.A(ori_ori_n770_), .B(ori_ori_n51_), .Y(ori_ori_n771_));
  NA2        o0743(.A(ori_ori_n278_), .B(ori_ori_n243_), .Y(ori_ori_n772_));
  AN2        o0744(.A(f), .B(d), .Y(ori_ori_n773_));
  NA3        o0745(.A(ori_ori_n434_), .B(ori_ori_n773_), .C(ori_ori_n76_), .Y(ori_ori_n774_));
  NO3        o0746(.A(ori_ori_n774_), .B(ori_ori_n65_), .C(ori_ori_n197_), .Y(ori_ori_n775_));
  NA2        o0747(.A(ori_ori_n772_), .B(ori_ori_n775_), .Y(ori_ori_n776_));
  NAi31      o0748(.An(ori_ori_n448_), .B(ori_ori_n776_), .C(ori_ori_n768_), .Y(ori_ori_n777_));
  NO2        o0749(.A(ori_ori_n582_), .B(ori_ori_n294_), .Y(ori_ori_n778_));
  NA3        o0750(.A(ori_ori_n150_), .B(ori_ori_n102_), .C(ori_ori_n101_), .Y(ori_ori_n779_));
  OAI220     o0751(.A0(ori_ori_n774_), .A1(ori_ori_n384_), .B0(ori_ori_n306_), .B1(ori_ori_n779_), .Y(ori_ori_n780_));
  NOi31      o0752(.An(ori_ori_n205_), .B(ori_ori_n780_), .C(ori_ori_n274_), .Y(ori_ori_n781_));
  NA2        o0753(.A(c), .B(ori_ori_n108_), .Y(ori_ori_n782_));
  NO2        o0754(.A(ori_ori_n782_), .B(ori_ori_n366_), .Y(ori_ori_n783_));
  NA3        o0755(.A(ori_ori_n783_), .B(ori_ori_n467_), .C(f), .Y(ori_ori_n784_));
  OR2        o0756(.A(ori_ori_n589_), .B(ori_ori_n494_), .Y(ori_ori_n785_));
  INV        o0757(.A(ori_ori_n785_), .Y(ori_ori_n786_));
  NA2        o0758(.A(ori_ori_n722_), .B(ori_ori_n104_), .Y(ori_ori_n787_));
  NA2        o0759(.A(ori_ori_n787_), .B(ori_ori_n786_), .Y(ori_ori_n788_));
  NA3        o0760(.A(ori_ori_n788_), .B(ori_ori_n784_), .C(ori_ori_n781_), .Y(ori_ori_n789_));
  NO4        o0761(.A(ori_ori_n789_), .B(ori_ori_n777_), .C(ori_ori_n766_), .D(ori_ori_n754_), .Y(ori_ori_n790_));
  OR2        o0762(.A(ori_ori_n774_), .B(ori_ori_n65_), .Y(ori_ori_n791_));
  NA2        o0763(.A(ori_ori_n742_), .B(g), .Y(ori_ori_n792_));
  AOI210     o0764(.A0(ori_ori_n792_), .A1(ori_ori_n266_), .B0(ori_ori_n791_), .Y(ori_ori_n793_));
  NO2        o0765(.A(ori_ori_n126_), .B(ori_ori_n122_), .Y(ori_ori_n794_));
  NO2        o0766(.A(ori_ori_n212_), .B(ori_ori_n206_), .Y(ori_ori_n795_));
  AOI220     o0767(.A0(ori_ori_n795_), .A1(ori_ori_n209_), .B0(ori_ori_n272_), .B1(ori_ori_n794_), .Y(ori_ori_n796_));
  NO2        o0768(.A(ori_ori_n384_), .B(ori_ori_n741_), .Y(ori_ori_n797_));
  INV        o0769(.A(ori_ori_n796_), .Y(ori_ori_n798_));
  NA2        o0770(.A(e), .B(d), .Y(ori_ori_n799_));
  OAI220     o0771(.A0(ori_ori_n799_), .A1(c), .B0(ori_ori_n289_), .B1(d), .Y(ori_ori_n800_));
  NA3        o0772(.A(ori_ori_n800_), .B(ori_ori_n411_), .C(ori_ori_n465_), .Y(ori_ori_n801_));
  AOI210     o0773(.A0(ori_ori_n472_), .A1(ori_ori_n166_), .B0(ori_ori_n212_), .Y(ori_ori_n802_));
  AOI210     o0774(.A0(ori_ori_n556_), .A1(ori_ori_n315_), .B0(ori_ori_n802_), .Y(ori_ori_n803_));
  INV        o0775(.A(ori_ori_n154_), .Y(ori_ori_n804_));
  NA2        o0776(.A(ori_ori_n775_), .B(ori_ori_n804_), .Y(ori_ori_n805_));
  NA3        o0777(.A(ori_ori_n155_), .B(ori_ori_n77_), .C(ori_ori_n33_), .Y(ori_ori_n806_));
  NA4        o0778(.A(ori_ori_n806_), .B(ori_ori_n805_), .C(ori_ori_n803_), .D(ori_ori_n801_), .Y(ori_ori_n807_));
  NO3        o0779(.A(ori_ori_n807_), .B(ori_ori_n798_), .C(ori_ori_n793_), .Y(ori_ori_n808_));
  OR2        o0780(.A(ori_ori_n628_), .B(ori_ori_n200_), .Y(ori_ori_n809_));
  OAI220     o0781(.A0(ori_ori_n555_), .A1(ori_ori_n57_), .B0(ori_ori_n270_), .B1(j), .Y(ori_ori_n810_));
  AOI220     o0782(.A0(ori_ori_n810_), .A1(ori_ori_n778_), .B0(ori_ori_n546_), .B1(ori_ori_n554_), .Y(ori_ori_n811_));
  OAI210     o0783(.A0(ori_ori_n747_), .A1(ori_ori_n156_), .B0(ori_ori_n811_), .Y(ori_ori_n812_));
  INV        o0784(.A(ori_ori_n242_), .Y(ori_ori_n813_));
  AN2        o0785(.A(ori_ori_n760_), .B(ori_ori_n751_), .Y(ori_ori_n814_));
  NO2        o0786(.A(ori_ori_n814_), .B(ori_ori_n812_), .Y(ori_ori_n815_));
  AO220      o0787(.A0(ori_ori_n411_), .A1(ori_ori_n669_), .B0(ori_ori_n161_), .B1(f), .Y(ori_ori_n816_));
  OAI210     o0788(.A0(ori_ori_n816_), .A1(ori_ori_n414_), .B0(ori_ori_n800_), .Y(ori_ori_n817_));
  NA2        o0789(.A(ori_ori_n753_), .B(ori_ori_n632_), .Y(ori_ori_n818_));
  AN4        o0790(.A(ori_ori_n818_), .B(ori_ori_n817_), .C(ori_ori_n815_), .D(ori_ori_n809_), .Y(ori_ori_n819_));
  NA4        o0791(.A(ori_ori_n819_), .B(ori_ori_n808_), .C(ori_ori_n790_), .D(ori_ori_n749_), .Y(ori12));
  NO2        o0792(.A(ori_ori_n409_), .B(c), .Y(ori_ori_n821_));
  NO4        o0793(.A(ori_ori_n398_), .B(ori_ori_n234_), .C(ori_ori_n528_), .D(ori_ori_n197_), .Y(ori_ori_n822_));
  NA2        o0794(.A(ori_ori_n822_), .B(ori_ori_n821_), .Y(ori_ori_n823_));
  NO2        o0795(.A(ori_ori_n409_), .B(ori_ori_n108_), .Y(ori_ori_n824_));
  NO2        o0796(.A(ori_ori_n756_), .B(ori_ori_n322_), .Y(ori_ori_n825_));
  NO2        o0797(.A(ori_ori_n589_), .B(ori_ori_n340_), .Y(ori_ori_n826_));
  AOI220     o0798(.A0(ori_ori_n826_), .A1(ori_ori_n496_), .B0(ori_ori_n825_), .B1(ori_ori_n824_), .Y(ori_ori_n827_));
  NA3        o0799(.A(ori_ori_n827_), .B(ori_ori_n823_), .C(ori_ori_n397_), .Y(ori_ori_n828_));
  AOI210     o0800(.A0(ori_ori_n215_), .A1(ori_ori_n305_), .B0(ori_ori_n187_), .Y(ori_ori_n829_));
  OR2        o0801(.A(ori_ori_n829_), .B(ori_ori_n822_), .Y(ori_ori_n830_));
  AOI210     o0802(.A0(ori_ori_n302_), .A1(ori_ori_n351_), .B0(ori_ori_n197_), .Y(ori_ori_n831_));
  OAI210     o0803(.A0(ori_ori_n831_), .A1(ori_ori_n830_), .B0(ori_ori_n361_), .Y(ori_ori_n832_));
  NO2        o0804(.A(ori_ori_n568_), .B(ori_ori_n244_), .Y(ori_ori_n833_));
  NO2        o0805(.A(ori_ori_n536_), .B(ori_ori_n750_), .Y(ori_ori_n834_));
  NO2        o0806(.A(ori_ori_n141_), .B(ori_ori_n218_), .Y(ori_ori_n835_));
  INV        o0807(.A(ori_ori_n832_), .Y(ori_ori_n836_));
  OR2        o0808(.A(ori_ori_n290_), .B(ori_ori_n824_), .Y(ori_ori_n837_));
  NA2        o0809(.A(ori_ori_n837_), .B(ori_ori_n323_), .Y(ori_ori_n838_));
  NO3        o0810(.A(ori_ori_n122_), .B(ori_ori_n142_), .C(ori_ori_n197_), .Y(ori_ori_n839_));
  NA2        o0811(.A(ori_ori_n839_), .B(ori_ori_n487_), .Y(ori_ori_n840_));
  NA4        o0812(.A(ori_ori_n399_), .B(ori_ori_n391_), .C(ori_ori_n167_), .D(g), .Y(ori_ori_n841_));
  NA3        o0813(.A(ori_ori_n841_), .B(ori_ori_n840_), .C(ori_ori_n838_), .Y(ori_ori_n842_));
  NO3        o0814(.A(ori_ori_n592_), .B(ori_ori_n84_), .C(ori_ori_n44_), .Y(ori_ori_n843_));
  NO4        o0815(.A(ori_ori_n843_), .B(ori_ori_n842_), .C(ori_ori_n836_), .D(ori_ori_n828_), .Y(ori_ori_n844_));
  NA2        o0816(.A(ori_ori_n505_), .B(ori_ori_n135_), .Y(ori_ori_n845_));
  NOi21      o0817(.An(ori_ori_n33_), .B(ori_ori_n582_), .Y(ori_ori_n846_));
  NA2        o0818(.A(ori_ori_n846_), .B(ori_ori_n845_), .Y(ori_ori_n847_));
  OAI210     o0819(.A0(ori_ori_n232_), .A1(ori_ori_n44_), .B0(ori_ori_n847_), .Y(ori_ori_n848_));
  INV        o0820(.A(ori_ori_n288_), .Y(ori_ori_n849_));
  NO2        o0821(.A(ori_ori_n48_), .B(ori_ori_n44_), .Y(ori_ori_n850_));
  NO2        o0822(.A(ori_ori_n462_), .B(ori_ori_n270_), .Y(ori_ori_n851_));
  INV        o0823(.A(ori_ori_n851_), .Y(ori_ori_n852_));
  NO2        o0824(.A(ori_ori_n852_), .B(ori_ori_n135_), .Y(ori_ori_n853_));
  INV        o0825(.A(ori_ori_n334_), .Y(ori_ori_n854_));
  NO4        o0826(.A(ori_ori_n854_), .B(ori_ori_n853_), .C(ori_ori_n849_), .D(ori_ori_n848_), .Y(ori_ori_n855_));
  NA2        o0827(.A(ori_ori_n315_), .B(g), .Y(ori_ori_n856_));
  NA2        o0828(.A(ori_ori_n153_), .B(i), .Y(ori_ori_n857_));
  NA2        o0829(.A(ori_ori_n45_), .B(i), .Y(ori_ori_n858_));
  OAI220     o0830(.A0(ori_ori_n858_), .A1(ori_ori_n186_), .B0(ori_ori_n857_), .B1(ori_ori_n84_), .Y(ori_ori_n859_));
  AOI210     o0831(.A0(ori_ori_n375_), .A1(ori_ori_n36_), .B0(ori_ori_n859_), .Y(ori_ori_n860_));
  NO2        o0832(.A(ori_ori_n135_), .B(ori_ori_n76_), .Y(ori_ori_n861_));
  OR2        o0833(.A(ori_ori_n861_), .B(ori_ori_n504_), .Y(ori_ori_n862_));
  NA2        o0834(.A(ori_ori_n505_), .B(ori_ori_n343_), .Y(ori_ori_n863_));
  AOI210     o0835(.A0(ori_ori_n863_), .A1(n), .B0(ori_ori_n862_), .Y(ori_ori_n864_));
  OAI220     o0836(.A0(ori_ori_n864_), .A1(ori_ori_n856_), .B0(ori_ori_n860_), .B1(ori_ori_n299_), .Y(ori_ori_n865_));
  NO2        o0837(.A(ori_ori_n589_), .B(ori_ori_n455_), .Y(ori_ori_n866_));
  NA3        o0838(.A(ori_ori_n310_), .B(ori_ori_n559_), .C(i), .Y(ori_ori_n867_));
  OAI210     o0839(.A0(ori_ori_n393_), .A1(ori_ori_n278_), .B0(ori_ori_n867_), .Y(ori_ori_n868_));
  OAI210     o0840(.A0(ori_ori_n868_), .A1(ori_ori_n866_), .B0(ori_ori_n604_), .Y(ori_ori_n869_));
  NA2        o0841(.A(ori_ori_n542_), .B(ori_ori_n106_), .Y(ori_ori_n870_));
  OR3        o0842(.A(ori_ori_n278_), .B(ori_ori_n389_), .C(f), .Y(ori_ori_n871_));
  NA3        o0843(.A(ori_ori_n559_), .B(ori_ori_n72_), .C(i), .Y(ori_ori_n872_));
  OA220      o0844(.A0(ori_ori_n872_), .A1(ori_ori_n870_), .B0(ori_ori_n871_), .B1(ori_ori_n535_), .Y(ori_ori_n873_));
  NA3        o0845(.A(ori_ori_n291_), .B(ori_ori_n110_), .C(g), .Y(ori_ori_n874_));
  AOI210     o0846(.A0(ori_ori_n601_), .A1(ori_ori_n874_), .B0(m), .Y(ori_ori_n875_));
  OAI210     o0847(.A0(ori_ori_n875_), .A1(ori_ori_n825_), .B0(ori_ori_n290_), .Y(ori_ori_n876_));
  INV        o0848(.A(ori_ori_n619_), .Y(ori_ori_n877_));
  INV        o0849(.A(ori_ori_n394_), .Y(ori_ori_n878_));
  INV        o0850(.A(ori_ori_n872_), .Y(ori_ori_n879_));
  AOI220     o0851(.A0(ori_ori_n879_), .A1(ori_ori_n240_), .B0(ori_ori_n878_), .B1(ori_ori_n877_), .Y(ori_ori_n880_));
  NA4        o0852(.A(ori_ori_n880_), .B(ori_ori_n876_), .C(ori_ori_n873_), .D(ori_ori_n869_), .Y(ori_ori_n881_));
  NO2        o0853(.A(ori_ori_n340_), .B(ori_ori_n83_), .Y(ori_ori_n882_));
  OAI210     o0854(.A0(ori_ori_n882_), .A1(ori_ori_n833_), .B0(ori_ori_n219_), .Y(ori_ori_n883_));
  NA2        o0855(.A(ori_ori_n591_), .B(ori_ori_n80_), .Y(ori_ori_n884_));
  NO2        o0856(.A(ori_ori_n417_), .B(ori_ori_n197_), .Y(ori_ori_n885_));
  AOI220     o0857(.A0(ori_ori_n885_), .A1(ori_ori_n344_), .B0(ori_ori_n837_), .B1(ori_ori_n201_), .Y(ori_ori_n886_));
  AOI220     o0858(.A0(ori_ori_n826_), .A1(ori_ori_n835_), .B0(ori_ori_n534_), .B1(ori_ori_n82_), .Y(ori_ori_n887_));
  NA4        o0859(.A(ori_ori_n887_), .B(ori_ori_n886_), .C(ori_ori_n884_), .D(ori_ori_n883_), .Y(ori_ori_n888_));
  OAI210     o0860(.A0(ori_ori_n878_), .A1(ori_ori_n834_), .B0(ori_ori_n496_), .Y(ori_ori_n889_));
  NA2        o0861(.A(ori_ori_n875_), .B(ori_ori_n824_), .Y(ori_ori_n890_));
  NA2        o0862(.A(ori_ori_n573_), .B(ori_ori_n487_), .Y(ori_ori_n891_));
  NA3        o0863(.A(ori_ori_n891_), .B(ori_ori_n890_), .C(ori_ori_n889_), .Y(ori_ori_n892_));
  NO4        o0864(.A(ori_ori_n892_), .B(ori_ori_n888_), .C(ori_ori_n881_), .D(ori_ori_n865_), .Y(ori_ori_n893_));
  NAi31      o0865(.An(ori_ori_n131_), .B(ori_ori_n377_), .C(n), .Y(ori_ori_n894_));
  NO3        o0866(.A(ori_ori_n116_), .B(ori_ori_n308_), .C(ori_ori_n757_), .Y(ori_ori_n895_));
  NO2        o0867(.A(ori_ori_n895_), .B(ori_ori_n894_), .Y(ori_ori_n896_));
  NO3        o0868(.A(ori_ori_n251_), .B(ori_ori_n131_), .C(ori_ori_n366_), .Y(ori_ori_n897_));
  AOI210     o0869(.A0(ori_ori_n897_), .A1(ori_ori_n456_), .B0(ori_ori_n896_), .Y(ori_ori_n898_));
  NA2        o0870(.A(ori_ori_n449_), .B(i), .Y(ori_ori_n899_));
  NA2        o0871(.A(ori_ori_n899_), .B(ori_ori_n898_), .Y(ori_ori_n900_));
  NA2        o0872(.A(ori_ori_n212_), .B(ori_ori_n157_), .Y(ori_ori_n901_));
  NO3        o0873(.A(ori_ori_n276_), .B(ori_ori_n399_), .C(ori_ori_n161_), .Y(ori_ori_n902_));
  NOi31      o0874(.An(ori_ori_n901_), .B(ori_ori_n902_), .C(ori_ori_n197_), .Y(ori_ori_n903_));
  NAi21      o0875(.An(ori_ori_n505_), .B(ori_ori_n885_), .Y(ori_ori_n904_));
  NA2        o0876(.A(ori_ori_n440_), .B(g), .Y(ori_ori_n905_));
  NA2        o0877(.A(ori_ori_n905_), .B(ori_ori_n904_), .Y(ori_ori_n906_));
  NA2        o0878(.A(ori_ori_n829_), .B(ori_ori_n821_), .Y(ori_ori_n907_));
  OAI210     o0879(.A0(ori_ori_n826_), .A1(ori_ori_n834_), .B0(ori_ori_n383_), .Y(ori_ori_n908_));
  NA3        o0880(.A(ori_ori_n908_), .B(ori_ori_n907_), .C(ori_ori_n553_), .Y(ori_ori_n909_));
  OAI210     o0881(.A0(ori_ori_n829_), .A1(ori_ori_n822_), .B0(ori_ori_n901_), .Y(ori_ori_n910_));
  NA3        o0882(.A(ori_ori_n863_), .B(ori_ori_n445_), .C(ori_ori_n45_), .Y(ori_ori_n911_));
  INV        o0883(.A(ori_ori_n298_), .Y(ori_ori_n912_));
  NA3        o0884(.A(ori_ori_n912_), .B(ori_ori_n911_), .C(ori_ori_n910_), .Y(ori_ori_n913_));
  OR2        o0885(.A(ori_ori_n913_), .B(ori_ori_n909_), .Y(ori_ori_n914_));
  NO4        o0886(.A(ori_ori_n914_), .B(ori_ori_n906_), .C(ori_ori_n903_), .D(ori_ori_n900_), .Y(ori_ori_n915_));
  NA4        o0887(.A(ori_ori_n915_), .B(ori_ori_n893_), .C(ori_ori_n855_), .D(ori_ori_n844_), .Y(ori13));
  AN2        o0888(.A(c), .B(b), .Y(ori_ori_n917_));
  NAi32      o0889(.An(d), .Bn(c), .C(e), .Y(ori_ori_n918_));
  AN2        o0890(.A(d), .B(c), .Y(ori_ori_n919_));
  NA2        o0891(.A(ori_ori_n919_), .B(ori_ori_n108_), .Y(ori_ori_n920_));
  NO3        o0892(.A(m), .B(i), .C(h), .Y(ori_ori_n921_));
  NA3        o0893(.A(k), .B(j), .C(i), .Y(ori_ori_n922_));
  NO2        o0894(.A(f), .B(c), .Y(ori_ori_n923_));
  NOi21      o0895(.An(ori_ori_n923_), .B(ori_ori_n398_), .Y(ori_ori_n924_));
  OR3        o0896(.A(n), .B(m), .C(i), .Y(ori_ori_n925_));
  AN3        o0897(.A(g), .B(f), .C(c), .Y(ori_ori_n926_));
  NA3        o0898(.A(l), .B(k), .C(j), .Y(ori_ori_n927_));
  NA2        o0899(.A(i), .B(h), .Y(ori_ori_n928_));
  NO3        o0900(.A(ori_ori_n928_), .B(ori_ori_n927_), .C(ori_ori_n122_), .Y(ori_ori_n929_));
  NO3        o0901(.A(ori_ori_n132_), .B(ori_ori_n258_), .C(ori_ori_n197_), .Y(ori_ori_n930_));
  NA3        o0902(.A(c), .B(b), .C(a), .Y(ori_ori_n931_));
  NO2        o0903(.A(ori_ori_n483_), .B(ori_ori_n540_), .Y(ori_ori_n932_));
  NA4        o0904(.A(ori_ori_n80_), .B(ori_ori_n79_), .C(g), .D(ori_ori_n196_), .Y(ori_ori_n933_));
  NA4        o0905(.A(ori_ori_n520_), .B(m), .C(ori_ori_n105_), .D(ori_ori_n196_), .Y(ori_ori_n934_));
  NA3        o0906(.A(ori_ori_n934_), .B(ori_ori_n335_), .C(ori_ori_n933_), .Y(ori_ori_n935_));
  NO2        o0907(.A(ori_ori_n935_), .B(ori_ori_n932_), .Y(ori_ori_n936_));
  NOi41      o0908(.An(ori_ori_n720_), .B(ori_ori_n762_), .C(ori_ori_n752_), .D(ori_ori_n646_), .Y(ori_ori_n937_));
  OAI220     o0909(.A0(ori_ori_n937_), .A1(ori_ori_n619_), .B0(ori_ori_n936_), .B1(ori_ori_n533_), .Y(ori_ori_n938_));
  NOi31      o0910(.An(m), .B(n), .C(f), .Y(ori_ori_n939_));
  NA2        o0911(.A(ori_ori_n939_), .B(ori_ori_n50_), .Y(ori_ori_n940_));
  AN2        o0912(.A(e), .B(c), .Y(ori_ori_n941_));
  NA2        o0913(.A(ori_ori_n941_), .B(a), .Y(ori_ori_n942_));
  OAI220     o0914(.A0(ori_ori_n942_), .A1(ori_ori_n940_), .B0(ori_ori_n785_), .B1(ori_ori_n382_), .Y(ori_ori_n943_));
  NA2        o0915(.A(ori_ori_n465_), .B(l), .Y(ori_ori_n944_));
  NO2        o0916(.A(ori_ori_n258_), .B(a), .Y(ori_ori_n945_));
  NO2        o0917(.A(ori_ori_n79_), .B(g), .Y(ori_ori_n946_));
  NO3        o0918(.A(ori_ori_n943_), .B(ori_ori_n938_), .C(ori_ori_n733_), .Y(ori_ori_n947_));
  NA2        o0919(.A(c), .B(b), .Y(ori_ori_n948_));
  NO2        o0920(.A(ori_ori_n631_), .B(ori_ori_n948_), .Y(ori_ori_n949_));
  OAI210     o0921(.A0(ori_ori_n770_), .A1(ori_ori_n745_), .B0(ori_ori_n371_), .Y(ori_ori_n950_));
  OAI210     o0922(.A0(ori_ori_n950_), .A1(ori_ori_n771_), .B0(ori_ori_n949_), .Y(ori_ori_n951_));
  NAi21      o0923(.An(ori_ori_n379_), .B(ori_ori_n949_), .Y(ori_ori_n952_));
  NA3        o0924(.A(ori_ori_n383_), .B(ori_ori_n510_), .C(f), .Y(ori_ori_n953_));
  OAI210     o0925(.A0(ori_ori_n499_), .A1(ori_ori_n38_), .B0(ori_ori_n945_), .Y(ori_ori_n954_));
  NA3        o0926(.A(ori_ori_n954_), .B(ori_ori_n953_), .C(ori_ori_n952_), .Y(ori_ori_n955_));
  OAI210     o0927(.A0(ori_ori_n242_), .A1(ori_ori_n260_), .B0(g), .Y(ori_ori_n956_));
  NAi21      o0928(.An(f), .B(d), .Y(ori_ori_n957_));
  NO2        o0929(.A(ori_ori_n957_), .B(ori_ori_n931_), .Y(ori_ori_n958_));
  INV        o0930(.A(ori_ori_n958_), .Y(ori_ori_n959_));
  NO2        o0931(.A(ori_ori_n956_), .B(ori_ori_n959_), .Y(ori_ori_n960_));
  AOI210     o0932(.A0(ori_ori_n960_), .A1(ori_ori_n106_), .B0(ori_ori_n955_), .Y(ori_ori_n961_));
  NA3        o0933(.A(ori_ori_n813_), .B(ori_ori_n944_), .C(ori_ori_n154_), .Y(ori_ori_n962_));
  NA2        o0934(.A(ori_ori_n402_), .B(ori_ori_n958_), .Y(ori_ori_n963_));
  NA4        o0935(.A(ori_ori_n963_), .B(ori_ori_n961_), .C(ori_ori_n951_), .D(ori_ori_n947_), .Y(ori00));
  NA2        o0936(.A(ori_ori_n797_), .B(ori_ori_n835_), .Y(ori_ori_n965_));
  INV        o0937(.A(ori_ori_n643_), .Y(ori_ori_n966_));
  NA2        o0938(.A(ori_ori_n966_), .B(ori_ori_n965_), .Y(ori_ori_n967_));
  NA2        o0939(.A(ori_ori_n467_), .B(f), .Y(ori_ori_n968_));
  OAI210     o0940(.A0(ori_ori_n895_), .A1(ori_ori_n39_), .B0(ori_ori_n575_), .Y(ori_ori_n969_));
  NA3        o0941(.A(ori_ori_n969_), .B(ori_ori_n239_), .C(n), .Y(ori_ori_n970_));
  AOI210     o0942(.A0(ori_ori_n970_), .A1(ori_ori_n968_), .B0(ori_ori_n920_), .Y(ori_ori_n971_));
  NO2        o0943(.A(ori_ori_n971_), .B(ori_ori_n967_), .Y(ori_ori_n972_));
  NA3        o0944(.A(ori_ori_n155_), .B(ori_ori_n45_), .C(ori_ori_n44_), .Y(ori_ori_n973_));
  NA3        o0945(.A(d), .B(ori_ori_n53_), .C(b), .Y(ori_ori_n974_));
  NO2        o0946(.A(ori_ori_n974_), .B(ori_ori_n973_), .Y(ori_ori_n975_));
  NO4        o0947(.A(ori_ori_n446_), .B(ori_ori_n324_), .C(ori_ori_n948_), .D(ori_ori_n56_), .Y(ori_ori_n976_));
  NA3        o0948(.A(ori_ori_n345_), .B(ori_ori_n204_), .C(g), .Y(ori_ori_n977_));
  OR2        o0949(.A(ori_ori_n977_), .B(ori_ori_n974_), .Y(ori_ori_n978_));
  NO2        o0950(.A(h), .B(g), .Y(ori_ori_n979_));
  NA4        o0951(.A(ori_ori_n456_), .B(ori_ori_n425_), .C(ori_ori_n979_), .D(ori_ori_n917_), .Y(ori_ori_n980_));
  OAI220     o0952(.A0(ori_ori_n483_), .A1(ori_ori_n540_), .B0(ori_ori_n84_), .B1(ori_ori_n83_), .Y(ori_ori_n981_));
  AOI220     o0953(.A0(ori_ori_n981_), .A1(ori_ori_n490_), .B0(ori_ori_n839_), .B1(ori_ori_n521_), .Y(ori_ori_n982_));
  AOI220     o0954(.A0(ori_ori_n285_), .A1(ori_ori_n228_), .B0(ori_ori_n163_), .B1(ori_ori_n139_), .Y(ori_ori_n983_));
  NA4        o0955(.A(ori_ori_n983_), .B(ori_ori_n982_), .C(ori_ori_n980_), .D(ori_ori_n978_), .Y(ori_ori_n984_));
  NO3        o0956(.A(ori_ori_n984_), .B(ori_ori_n976_), .C(ori_ori_n246_), .Y(ori_ori_n985_));
  AOI210     o0957(.A0(ori_ori_n228_), .A1(ori_ori_n315_), .B0(ori_ori_n524_), .Y(ori_ori_n986_));
  NA2        o0958(.A(ori_ori_n986_), .B(ori_ori_n144_), .Y(ori_ori_n987_));
  NO2        o0959(.A(ori_ori_n220_), .B(ori_ori_n167_), .Y(ori_ori_n988_));
  NA2        o0960(.A(ori_ori_n988_), .B(ori_ori_n383_), .Y(ori_ori_n989_));
  INV        o0961(.A(ori_ori_n989_), .Y(ori_ori_n990_));
  NO3        o0962(.A(ori_ori_n990_), .B(ori_ori_n987_), .C(ori_ori_n476_), .Y(ori_ori_n991_));
  AN3        o0963(.A(ori_ori_n991_), .B(ori_ori_n985_), .C(ori_ori_n522_), .Y(ori_ori_n992_));
  NA3        o0964(.A(ori_ori_n939_), .B(ori_ori_n542_), .C(ori_ori_n424_), .Y(ori_ori_n993_));
  NA2        o0965(.A(ori_ori_n993_), .B(ori_ori_n222_), .Y(ori_ori_n994_));
  NA2        o0966(.A(ori_ori_n935_), .B(ori_ori_n490_), .Y(ori_ori_n995_));
  NA4        o0967(.A(ori_ori_n578_), .B(ori_ori_n192_), .C(ori_ori_n204_), .D(ori_ori_n153_), .Y(ori_ori_n996_));
  NA2        o0968(.A(ori_ori_n996_), .B(ori_ori_n995_), .Y(ori_ori_n997_));
  NO2        o0969(.A(ori_ori_n423_), .B(ori_ori_n111_), .Y(ori_ori_n998_));
  NA2        o0970(.A(ori_ori_n998_), .B(ori_ori_n962_), .Y(ori_ori_n999_));
  NO2        o0971(.A(ori_ori_n200_), .B(ori_ori_n197_), .Y(ori_ori_n1000_));
  NA2        o0972(.A(n), .B(e), .Y(ori_ori_n1001_));
  NO2        o0973(.A(ori_ori_n1001_), .B(ori_ori_n137_), .Y(ori_ori_n1002_));
  AOI220     o0974(.A0(ori_ori_n1002_), .A1(ori_ori_n252_), .B0(ori_ori_n755_), .B1(ori_ori_n1000_), .Y(ori_ori_n1003_));
  OAI210     o0975(.A0(ori_ori_n325_), .A1(ori_ori_n280_), .B0(ori_ori_n404_), .Y(ori_ori_n1004_));
  NA3        o0976(.A(ori_ori_n1004_), .B(ori_ori_n1003_), .C(ori_ori_n999_), .Y(ori_ori_n1005_));
  NA2        o0977(.A(ori_ori_n1002_), .B(ori_ori_n759_), .Y(ori_ori_n1006_));
  AOI220     o0978(.A0(ori_ori_n846_), .A1(ori_ori_n521_), .B0(ori_ori_n578_), .B1(ori_ori_n225_), .Y(ori_ori_n1007_));
  NO2        o0979(.A(ori_ori_n60_), .B(h), .Y(ori_ori_n1008_));
  NA2        o0980(.A(ori_ori_n1007_), .B(ori_ori_n1006_), .Y(ori_ori_n1009_));
  NO4        o0981(.A(ori_ori_n1009_), .B(ori_ori_n1005_), .C(ori_ori_n997_), .D(ori_ori_n994_), .Y(ori_ori_n1010_));
  NA2        o0982(.A(ori_ori_n746_), .B(ori_ori_n678_), .Y(ori_ori_n1011_));
  NA4        o0983(.A(ori_ori_n1011_), .B(ori_ori_n1010_), .C(ori_ori_n992_), .D(ori_ori_n972_), .Y(ori01));
  NO2        o0984(.A(ori_ori_n437_), .B(ori_ori_n256_), .Y(ori_ori_n1013_));
  NA2        o0985(.A(ori_ori_n356_), .B(i), .Y(ori_ori_n1014_));
  NA3        o0986(.A(ori_ori_n1014_), .B(ori_ori_n1013_), .C(ori_ori_n907_), .Y(ori_ori_n1015_));
  NA2        o0987(.A(ori_ori_n534_), .B(ori_ori_n82_), .Y(ori_ori_n1016_));
  NA2        o0988(.A(ori_ori_n505_), .B(ori_ori_n250_), .Y(ori_ori_n1017_));
  NA2        o0989(.A(ori_ori_n851_), .B(ori_ori_n1017_), .Y(ori_ori_n1018_));
  NA4        o0990(.A(ori_ori_n1018_), .B(ori_ori_n1016_), .C(ori_ori_n811_), .D(ori_ori_n300_), .Y(ori_ori_n1019_));
  NA2        o0991(.A(ori_ori_n44_), .B(f), .Y(ori_ori_n1020_));
  NA2        o0992(.A(ori_ori_n638_), .B(ori_ori_n89_), .Y(ori_ori_n1021_));
  NO2        o0993(.A(ori_ori_n1021_), .B(ori_ori_n1020_), .Y(ori_ori_n1022_));
  NA2        o0994(.A(ori_ori_n110_), .B(l), .Y(ori_ori_n1023_));
  OA220      o0995(.A0(ori_ori_n1023_), .A1(ori_ori_n531_), .B0(ori_ori_n590_), .B1(ori_ori_n335_), .Y(ori_ori_n1024_));
  NAi41      o0996(.An(ori_ori_n152_), .B(ori_ori_n1024_), .C(ori_ori_n996_), .D(ori_ori_n796_), .Y(ori_ori_n1025_));
  NO2        o0997(.A(ori_ori_n603_), .B(ori_ori_n470_), .Y(ori_ori_n1026_));
  NA4        o0998(.A(ori_ori_n638_), .B(ori_ori_n89_), .C(ori_ori_n44_), .D(ori_ori_n196_), .Y(ori_ori_n1027_));
  OA220      o0999(.A0(ori_ori_n1027_), .A1(ori_ori_n598_), .B0(ori_ori_n181_), .B1(ori_ori_n179_), .Y(ori_ori_n1028_));
  NA3        o1000(.A(ori_ori_n1028_), .B(ori_ori_n1026_), .C(ori_ori_n127_), .Y(ori_ori_n1029_));
  NO4        o1001(.A(ori_ori_n1029_), .B(ori_ori_n1025_), .C(ori_ori_n1019_), .D(ori_ori_n1015_), .Y(ori_ori_n1030_));
  INV        o1002(.A(ori_ori_n977_), .Y(ori_ori_n1031_));
  NA2        o1003(.A(ori_ori_n1031_), .B(ori_ori_n487_), .Y(ori_ori_n1032_));
  AOI210     o1004(.A0(ori_ori_n190_), .A1(ori_ori_n81_), .B0(ori_ori_n196_), .Y(ori_ori_n1033_));
  OAI210     o1005(.A0(ori_ori_n723_), .A1(ori_ori_n383_), .B0(ori_ori_n1033_), .Y(ori_ori_n1034_));
  AN3        o1006(.A(m), .B(l), .C(k), .Y(ori_ori_n1035_));
  OAI210     o1007(.A0(ori_ori_n326_), .A1(ori_ori_n33_), .B0(ori_ori_n1035_), .Y(ori_ori_n1036_));
  OR2        o1008(.A(ori_ori_n1036_), .B(ori_ori_n299_), .Y(ori_ori_n1037_));
  NA3        o1009(.A(ori_ori_n1037_), .B(ori_ori_n1034_), .C(ori_ori_n1032_), .Y(ori_ori_n1038_));
  NA2        o1010(.A(ori_ori_n538_), .B(ori_ori_n110_), .Y(ori_ori_n1039_));
  INV        o1011(.A(ori_ori_n1039_), .Y(ori_ori_n1040_));
  NA2        o1012(.A(ori_ori_n255_), .B(ori_ori_n181_), .Y(ori_ori_n1041_));
  OAI210     o1013(.A0(ori_ori_n1041_), .A1(ori_ori_n347_), .B0(ori_ori_n594_), .Y(ori_ori_n1042_));
  OAI210     o1014(.A0(ori_ori_n1022_), .A1(ori_ori_n293_), .B0(ori_ori_n604_), .Y(ori_ori_n1043_));
  NA3        o1015(.A(ori_ori_n1043_), .B(ori_ori_n1042_), .C(ori_ori_n702_), .Y(ori_ori_n1044_));
  NO3        o1016(.A(ori_ori_n1044_), .B(ori_ori_n1040_), .C(ori_ori_n1038_), .Y(ori_ori_n1045_));
  NA2        o1017(.A(ori_ori_n463_), .B(ori_ori_n55_), .Y(ori_ori_n1046_));
  NO2        o1018(.A(ori_ori_n1027_), .B(ori_ori_n870_), .Y(ori_ori_n1047_));
  NO2        o1019(.A(ori_ori_n193_), .B(ori_ori_n104_), .Y(ori_ori_n1048_));
  NO3        o1020(.A(ori_ori_n1048_), .B(ori_ori_n1047_), .C(ori_ori_n975_), .Y(ori_ori_n1049_));
  NA3        o1021(.A(ori_ori_n1049_), .B(ori_ori_n1046_), .C(ori_ori_n677_), .Y(ori_ori_n1050_));
  NO2        o1022(.A(ori_ori_n857_), .B(ori_ori_n214_), .Y(ori_ori_n1051_));
  NO2        o1023(.A(ori_ori_n858_), .B(ori_ori_n507_), .Y(ori_ori_n1052_));
  OAI210     o1024(.A0(ori_ori_n1052_), .A1(ori_ori_n1051_), .B0(ori_ori_n308_), .Y(ori_ori_n1053_));
  NA2        o1025(.A(ori_ori_n516_), .B(ori_ori_n514_), .Y(ori_ori_n1054_));
  NO3        o1026(.A(ori_ori_n71_), .B(ori_ori_n270_), .C(ori_ori_n44_), .Y(ori_ori_n1055_));
  NA2        o1027(.A(ori_ori_n1055_), .B(ori_ori_n504_), .Y(ori_ori_n1056_));
  NA3        o1028(.A(ori_ori_n1056_), .B(ori_ori_n1054_), .C(ori_ori_n599_), .Y(ori_ori_n1057_));
  OR2        o1029(.A(ori_ori_n977_), .B(ori_ori_n974_), .Y(ori_ori_n1058_));
  NA2        o1030(.A(ori_ori_n1055_), .B(ori_ori_n726_), .Y(ori_ori_n1059_));
  NA3        o1031(.A(ori_ori_n1059_), .B(ori_ori_n1058_), .C(ori_ori_n348_), .Y(ori_ori_n1060_));
  NOi41      o1032(.An(ori_ori_n1053_), .B(ori_ori_n1060_), .C(ori_ori_n1057_), .D(ori_ori_n1050_), .Y(ori_ori_n1061_));
  NO2        o1033(.A(ori_ori_n121_), .B(ori_ori_n44_), .Y(ori_ori_n1062_));
  NO2        o1034(.A(ori_ori_n44_), .B(ori_ori_n39_), .Y(ori_ori_n1063_));
  AO220      o1035(.A0(ori_ori_n1063_), .A1(ori_ori_n556_), .B0(ori_ori_n1062_), .B1(ori_ori_n636_), .Y(ori_ori_n1064_));
  NA2        o1036(.A(ori_ori_n1064_), .B(ori_ori_n308_), .Y(ori_ori_n1065_));
  INV        o1037(.A(ori_ori_n125_), .Y(ori_ori_n1066_));
  NO3        o1038(.A(ori_ori_n928_), .B(ori_ori_n162_), .C(ori_ori_n79_), .Y(ori_ori_n1067_));
  AOI220     o1039(.A0(ori_ori_n1067_), .A1(ori_ori_n1066_), .B0(ori_ori_n1055_), .B1(ori_ori_n861_), .Y(ori_ori_n1068_));
  NA2        o1040(.A(ori_ori_n1068_), .B(ori_ori_n1065_), .Y(ori_ori_n1069_));
  NO2        o1041(.A(ori_ori_n548_), .B(ori_ori_n547_), .Y(ori_ori_n1070_));
  NO4        o1042(.A(ori_ori_n928_), .B(ori_ori_n1070_), .C(ori_ori_n160_), .D(ori_ori_n79_), .Y(ori_ori_n1071_));
  NO3        o1043(.A(ori_ori_n1071_), .B(ori_ori_n1069_), .C(ori_ori_n567_), .Y(ori_ori_n1072_));
  NA4        o1044(.A(ori_ori_n1072_), .B(ori_ori_n1061_), .C(ori_ori_n1045_), .D(ori_ori_n1030_), .Y(ori06));
  NO2        o1045(.A(ori_ori_n206_), .B(ori_ori_n96_), .Y(ori_ori_n1074_));
  OAI210     o1046(.A0(ori_ori_n1074_), .A1(ori_ori_n1067_), .B0(ori_ori_n344_), .Y(ori_ori_n1075_));
  INV        o1047(.A(ori_ori_n721_), .Y(ori_ori_n1076_));
  OR2        o1048(.A(ori_ori_n1076_), .B(ori_ori_n785_), .Y(ori_ori_n1077_));
  NA3        o1049(.A(ori_ori_n1077_), .B(ori_ori_n1075_), .C(ori_ori_n1053_), .Y(ori_ori_n1078_));
  NO3        o1050(.A(ori_ori_n1078_), .B(ori_ori_n1057_), .C(ori_ori_n238_), .Y(ori_ori_n1079_));
  NO2        o1051(.A(ori_ori_n270_), .B(ori_ori_n44_), .Y(ori_ori_n1080_));
  AOI210     o1052(.A0(ori_ori_n1080_), .A1(ori_ori_n862_), .B0(ori_ori_n1051_), .Y(ori_ori_n1081_));
  AOI210     o1053(.A0(ori_ori_n1080_), .A1(ori_ori_n508_), .B0(ori_ori_n1064_), .Y(ori_ori_n1082_));
  AOI210     o1054(.A0(ori_ori_n1082_), .A1(ori_ori_n1081_), .B0(ori_ori_n305_), .Y(ori_ori_n1083_));
  OAI210     o1055(.A0(ori_ori_n81_), .A1(ori_ori_n39_), .B0(ori_ori_n602_), .Y(ori_ori_n1084_));
  NA2        o1056(.A(ori_ori_n1084_), .B(ori_ori_n571_), .Y(ori_ori_n1085_));
  NO2        o1057(.A(ori_ori_n472_), .B(ori_ori_n157_), .Y(ori_ori_n1086_));
  NO2        o1058(.A(ori_ori_n543_), .B(ori_ori_n940_), .Y(ori_ori_n1087_));
  OAI210     o1059(.A0(ori_ori_n418_), .A1(ori_ori_n229_), .B0(ori_ori_n806_), .Y(ori_ori_n1088_));
  NO3        o1060(.A(ori_ori_n1088_), .B(ori_ori_n1087_), .C(ori_ori_n1086_), .Y(ori_ori_n1089_));
  NA2        o1061(.A(ori_ori_n1089_), .B(ori_ori_n1085_), .Y(ori_ori_n1090_));
  AN2        o1062(.A(ori_ori_n846_), .B(ori_ori_n574_), .Y(ori_ori_n1091_));
  NO3        o1063(.A(ori_ori_n1091_), .B(ori_ori_n1090_), .C(ori_ori_n1083_), .Y(ori_ori_n1092_));
  OAI220     o1064(.A0(ori_ori_n660_), .A1(ori_ori_n46_), .B0(ori_ori_n206_), .B1(ori_ori_n550_), .Y(ori_ori_n1093_));
  NA2        o1065(.A(ori_ori_n329_), .B(ori_ori_n1093_), .Y(ori_ori_n1094_));
  NO3        o1066(.A(ori_ori_n224_), .B(ori_ori_n96_), .C(ori_ori_n258_), .Y(ori_ori_n1095_));
  OAI220     o1067(.A0(ori_ori_n628_), .A1(ori_ori_n229_), .B0(ori_ori_n469_), .B1(ori_ori_n472_), .Y(ori_ori_n1096_));
  INV        o1068(.A(k), .Y(ori_ori_n1097_));
  NO3        o1069(.A(ori_ori_n1097_), .B(ori_ori_n540_), .C(j), .Y(ori_ori_n1098_));
  NO3        o1070(.A(ori_ori_n1096_), .B(ori_ori_n1095_), .C(ori_ori_n943_), .Y(ori_ori_n1099_));
  NA3        o1071(.A(ori_ori_n710_), .B(ori_ori_n709_), .C(ori_ori_n392_), .Y(ori_ori_n1100_));
  NAi31      o1072(.An(ori_ori_n670_), .B(ori_ori_n1100_), .C(ori_ori_n189_), .Y(ori_ori_n1101_));
  NA4        o1073(.A(ori_ori_n1101_), .B(ori_ori_n1099_), .C(ori_ori_n1094_), .D(ori_ori_n1007_), .Y(ori_ori_n1102_));
  NA2        o1074(.A(ori_ori_n516_), .B(ori_ori_n404_), .Y(ori_ori_n1103_));
  NA2        o1075(.A(ori_ori_n1098_), .B(ori_ori_n706_), .Y(ori_ori_n1104_));
  NA2        o1076(.A(ori_ori_n1104_), .B(ori_ori_n1103_), .Y(ori_ori_n1105_));
  AN2        o1077(.A(ori_ori_n822_), .B(ori_ori_n821_), .Y(ori_ori_n1106_));
  NO3        o1078(.A(ori_ori_n1106_), .B(ori_ori_n459_), .C(ori_ori_n440_), .Y(ori_ori_n1107_));
  NA2        o1079(.A(ori_ori_n1107_), .B(ori_ori_n1059_), .Y(ori_ori_n1108_));
  NAi21      o1080(.An(j), .B(i), .Y(ori_ori_n1109_));
  NO4        o1081(.A(ori_ori_n1070_), .B(ori_ori_n1109_), .C(ori_ori_n398_), .D(ori_ori_n216_), .Y(ori_ori_n1110_));
  NO4        o1082(.A(ori_ori_n1110_), .B(ori_ori_n1108_), .C(ori_ori_n1105_), .D(ori_ori_n1102_), .Y(ori_ori_n1111_));
  NA4        o1083(.A(ori_ori_n1111_), .B(ori_ori_n1092_), .C(ori_ori_n1079_), .D(ori_ori_n1072_), .Y(ori07));
  NAi32      o1084(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1113_));
  NO3        o1085(.A(ori_ori_n1113_), .B(g), .C(f), .Y(ori_ori_n1114_));
  NAi21      o1086(.An(f), .B(c), .Y(ori_ori_n1115_));
  OR2        o1087(.A(e), .B(d), .Y(ori_ori_n1116_));
  NOi31      o1088(.An(n), .B(m), .C(b), .Y(ori_ori_n1117_));
  NOi41      o1089(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1118_));
  NO2        o1090(.A(ori_ori_n922_), .B(ori_ori_n275_), .Y(ori_ori_n1119_));
  NA2        o1091(.A(ori_ori_n495_), .B(ori_ori_n72_), .Y(ori_ori_n1120_));
  NA2        o1092(.A(ori_ori_n1008_), .B(ori_ori_n264_), .Y(ori_ori_n1121_));
  NA2        o1093(.A(ori_ori_n1121_), .B(ori_ori_n1120_), .Y(ori_ori_n1122_));
  NO2        o1094(.A(ori_ori_n1122_), .B(ori_ori_n1114_), .Y(ori_ori_n1123_));
  NO3        o1095(.A(e), .B(d), .C(c), .Y(ori_ori_n1124_));
  NO2        o1096(.A(ori_ori_n122_), .B(ori_ori_n197_), .Y(ori_ori_n1125_));
  NA2        o1097(.A(ori_ori_n1125_), .B(ori_ori_n1124_), .Y(ori_ori_n1126_));
  INV        o1098(.A(ori_ori_n1126_), .Y(ori_ori_n1127_));
  NA3        o1099(.A(ori_ori_n625_), .B(ori_ori_n611_), .C(ori_ori_n105_), .Y(ori_ori_n1128_));
  NO2        o1100(.A(ori_ori_n1128_), .B(ori_ori_n44_), .Y(ori_ori_n1129_));
  NO2        o1101(.A(l), .B(k), .Y(ori_ori_n1130_));
  NO3        o1102(.A(ori_ori_n398_), .B(d), .C(c), .Y(ori_ori_n1131_));
  NO2        o1103(.A(ori_ori_n1129_), .B(ori_ori_n1127_), .Y(ori_ori_n1132_));
  NO2        o1104(.A(g), .B(c), .Y(ori_ori_n1133_));
  NO2        o1105(.A(ori_ori_n409_), .B(a), .Y(ori_ori_n1134_));
  NA2        o1106(.A(ori_ori_n1134_), .B(ori_ori_n106_), .Y(ori_ori_n1135_));
  NA2        o1107(.A(ori_ori_n128_), .B(ori_ori_n204_), .Y(ori_ori_n1136_));
  NO2        o1108(.A(ori_ori_n1136_), .B(ori_ori_n1228_), .Y(ori_ori_n1137_));
  NO2        o1109(.A(ori_ori_n676_), .B(ori_ori_n173_), .Y(ori_ori_n1138_));
  NOi31      o1110(.An(m), .B(n), .C(b), .Y(ori_ori_n1139_));
  NOi31      o1111(.An(f), .B(d), .C(c), .Y(ori_ori_n1140_));
  NA2        o1112(.A(ori_ori_n1140_), .B(ori_ori_n1139_), .Y(ori_ori_n1141_));
  INV        o1113(.A(ori_ori_n1141_), .Y(ori_ori_n1142_));
  NO3        o1114(.A(ori_ori_n1142_), .B(ori_ori_n1138_), .C(ori_ori_n1137_), .Y(ori_ori_n1143_));
  NA2        o1115(.A(ori_ori_n926_), .B(ori_ori_n425_), .Y(ori_ori_n1144_));
  NO2        o1116(.A(ori_ori_n1144_), .B(ori_ori_n398_), .Y(ori_ori_n1145_));
  NO3        o1117(.A(ori_ori_n40_), .B(i), .C(h), .Y(ori_ori_n1146_));
  NO2        o1118(.A(ori_ori_n921_), .B(ori_ori_n1145_), .Y(ori_ori_n1147_));
  AN3        o1119(.A(ori_ori_n1147_), .B(ori_ori_n1143_), .C(ori_ori_n1135_), .Y(ori_ori_n1148_));
  NA2        o1120(.A(ori_ori_n1117_), .B(ori_ori_n341_), .Y(ori_ori_n1149_));
  INV        o1121(.A(ori_ori_n1149_), .Y(ori_ori_n1150_));
  INV        o1122(.A(ori_ori_n929_), .Y(ori_ori_n1151_));
  NAi21      o1123(.An(ori_ori_n1150_), .B(ori_ori_n1151_), .Y(ori_ori_n1152_));
  NO4        o1124(.A(ori_ori_n122_), .B(g), .C(f), .D(e), .Y(ori_ori_n1153_));
  NA2        o1125(.A(ori_ori_n30_), .B(h), .Y(ori_ori_n1154_));
  NO2        o1126(.A(ori_ori_n1154_), .B(ori_ori_n925_), .Y(ori_ori_n1155_));
  NA2        o1127(.A(ori_ori_n1118_), .B(ori_ori_n1130_), .Y(ori_ori_n1156_));
  INV        o1128(.A(ori_ori_n1156_), .Y(ori_ori_n1157_));
  OR3        o1129(.A(ori_ori_n494_), .B(ori_ori_n493_), .C(ori_ori_n105_), .Y(ori_ori_n1158_));
  NA2        o1130(.A(ori_ori_n939_), .B(ori_ori_n366_), .Y(ori_ori_n1159_));
  NO2        o1131(.A(ori_ori_n1159_), .B(ori_ori_n391_), .Y(ori_ori_n1160_));
  AO210      o1132(.A0(ori_ori_n1160_), .A1(ori_ori_n108_), .B0(ori_ori_n1157_), .Y(ori_ori_n1161_));
  NO3        o1133(.A(ori_ori_n1161_), .B(ori_ori_n1155_), .C(ori_ori_n1152_), .Y(ori_ori_n1162_));
  NA4        o1134(.A(ori_ori_n1162_), .B(ori_ori_n1148_), .C(ori_ori_n1132_), .D(ori_ori_n1123_), .Y(ori_ori_n1163_));
  NO2        o1135(.A(ori_ori_n948_), .B(ori_ori_n103_), .Y(ori_ori_n1164_));
  NO2        o1136(.A(ori_ori_n353_), .B(j), .Y(ori_ori_n1165_));
  NA2        o1137(.A(ori_ori_n1146_), .B(ori_ori_n939_), .Y(ori_ori_n1166_));
  NA2        o1138(.A(ori_ori_n924_), .B(ori_ori_n140_), .Y(ori_ori_n1167_));
  NA2        o1139(.A(ori_ori_n1167_), .B(ori_ori_n1166_), .Y(ori_ori_n1168_));
  NA2        o1140(.A(ori_ori_n1165_), .B(ori_ori_n149_), .Y(ori_ori_n1169_));
  INV        o1141(.A(ori_ori_n1169_), .Y(ori_ori_n1170_));
  NO2        o1142(.A(ori_ori_n1170_), .B(ori_ori_n1168_), .Y(ori_ori_n1171_));
  INV        o1143(.A(ori_ori_n48_), .Y(ori_ori_n1172_));
  NA2        o1144(.A(ori_ori_n1172_), .B(ori_ori_n979_), .Y(ori_ori_n1173_));
  INV        o1145(.A(ori_ori_n1173_), .Y(ori_ori_n1174_));
  NO2        o1146(.A(ori_ori_n595_), .B(ori_ori_n162_), .Y(ori_ori_n1175_));
  NO2        o1147(.A(ori_ori_n1175_), .B(ori_ori_n1174_), .Y(ori_ori_n1176_));
  NO3        o1148(.A(ori_ori_n931_), .B(ori_ori_n1116_), .C(ori_ori_n48_), .Y(ori_ori_n1177_));
  NO2        o1149(.A(ori_ori_n925_), .B(h), .Y(ori_ori_n1178_));
  NA3        o1150(.A(ori_ori_n1164_), .B(ori_ori_n425_), .C(f), .Y(ori_ori_n1179_));
  NO2        o1151(.A(ori_ori_n1227_), .B(ori_ori_n1179_), .Y(ori_ori_n1180_));
  NO2        o1152(.A(ori_ori_n1109_), .B(ori_ori_n160_), .Y(ori_ori_n1181_));
  NOi21      o1153(.An(d), .B(f), .Y(ori_ori_n1182_));
  NO2        o1154(.A(ori_ori_n1180_), .B(ori_ori_n1178_), .Y(ori_ori_n1183_));
  NA3        o1155(.A(ori_ori_n1183_), .B(ori_ori_n1176_), .C(ori_ori_n1171_), .Y(ori_ori_n1184_));
  NA2        o1156(.A(h), .B(ori_ori_n1119_), .Y(ori_ori_n1185_));
  OAI210     o1157(.A0(ori_ori_n1153_), .A1(ori_ori_n1117_), .B0(ori_ori_n782_), .Y(ori_ori_n1186_));
  NO2        o1158(.A(ori_ori_n918_), .B(ori_ori_n122_), .Y(ori_ori_n1187_));
  NA2        o1159(.A(ori_ori_n1187_), .B(ori_ori_n555_), .Y(ori_ori_n1188_));
  NA3        o1160(.A(ori_ori_n1188_), .B(ori_ori_n1186_), .C(ori_ori_n1185_), .Y(ori_ori_n1189_));
  NA2        o1161(.A(ori_ori_n1133_), .B(ori_ori_n1182_), .Y(ori_ori_n1190_));
  NO2        o1162(.A(ori_ori_n1190_), .B(m), .Y(ori_ori_n1191_));
  NO2        o1163(.A(ori_ori_n141_), .B(ori_ori_n167_), .Y(ori_ori_n1192_));
  OAI210     o1164(.A0(ori_ori_n1192_), .A1(ori_ori_n103_), .B0(ori_ori_n1139_), .Y(ori_ori_n1193_));
  INV        o1165(.A(ori_ori_n1193_), .Y(ori_ori_n1194_));
  NO3        o1166(.A(ori_ori_n1194_), .B(ori_ori_n1191_), .C(ori_ori_n1189_), .Y(ori_ori_n1195_));
  NO2        o1167(.A(ori_ori_n1115_), .B(e), .Y(ori_ori_n1196_));
  NA2        o1168(.A(ori_ori_n1196_), .B(ori_ori_n364_), .Y(ori_ori_n1197_));
  BUFFER     o1169(.A(ori_ori_n122_), .Y(ori_ori_n1198_));
  NO2        o1170(.A(ori_ori_n1198_), .B(ori_ori_n1197_), .Y(ori_ori_n1199_));
  NO2        o1171(.A(ori_ori_n1158_), .B(ori_ori_n322_), .Y(ori_ori_n1200_));
  NO2        o1172(.A(ori_ori_n1200_), .B(ori_ori_n1199_), .Y(ori_ori_n1201_));
  NA2        o1173(.A(ori_ori_n1196_), .B(ori_ori_n165_), .Y(ori_ori_n1202_));
  INV        o1174(.A(ori_ori_n1202_), .Y(ori_ori_n1203_));
  AOI210     o1175(.A0(i), .A1(ori_ori_n1131_), .B0(ori_ori_n1177_), .Y(ori_ori_n1204_));
  INV        o1176(.A(ori_ori_n946_), .Y(ori_ori_n1205_));
  OAI210     o1177(.A0(ori_ori_n1205_), .A1(ori_ori_n61_), .B0(ori_ori_n1204_), .Y(ori_ori_n1206_));
  OR2        o1178(.A(h), .B(ori_ori_n493_), .Y(ori_ori_n1207_));
  NO2        o1179(.A(ori_ori_n1207_), .B(ori_ori_n160_), .Y(ori_ori_n1208_));
  NA2        o1180(.A(ori_ori_n930_), .B(ori_ori_n204_), .Y(ori_ori_n1209_));
  NO2        o1181(.A(ori_ori_n48_), .B(l), .Y(ori_ori_n1210_));
  INV        o1182(.A(ori_ori_n442_), .Y(ori_ori_n1211_));
  NA2        o1183(.A(ori_ori_n1211_), .B(ori_ori_n1210_), .Y(ori_ori_n1212_));
  NA2        o1184(.A(ori_ori_n1212_), .B(ori_ori_n1209_), .Y(ori_ori_n1213_));
  NO4        o1185(.A(ori_ori_n1213_), .B(ori_ori_n1208_), .C(ori_ori_n1206_), .D(ori_ori_n1203_), .Y(ori_ori_n1214_));
  NA3        o1186(.A(ori_ori_n1214_), .B(ori_ori_n1201_), .C(ori_ori_n1195_), .Y(ori_ori_n1215_));
  NA3        o1187(.A(ori_ori_n850_), .B(ori_ori_n128_), .C(ori_ori_n45_), .Y(ori_ori_n1216_));
  INV        o1188(.A(ori_ori_n1216_), .Y(ori_ori_n1217_));
  NA2        o1189(.A(ori_ori_n1181_), .B(h), .Y(ori_ori_n1218_));
  INV        o1190(.A(ori_ori_n1218_), .Y(ori_ori_n1219_));
  NO2        o1191(.A(ori_ori_n1219_), .B(ori_ori_n1217_), .Y(ori_ori_n1220_));
  NO2        o1192(.A(ori_ori_n1159_), .B(d), .Y(ori_ori_n1221_));
  INV        o1193(.A(ori_ori_n1221_), .Y(ori_ori_n1222_));
  NA2        o1194(.A(ori_ori_n1222_), .B(ori_ori_n1220_), .Y(ori_ori_n1223_));
  OR4        o1195(.A(ori_ori_n1223_), .B(ori_ori_n1215_), .C(ori_ori_n1184_), .D(ori_ori_n1163_), .Y(ori04));
  INV        o1196(.A(ori_ori_n106_), .Y(ori_ori_n1227_));
  INV        o1197(.A(h), .Y(ori_ori_n1228_));
  ZERO       o1198(.Y(ori02));
  ZERO       o1199(.Y(ori03));
  ZERO       o1200(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO4        m0025(.A(mai_mai_n53_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n54_));
  AOI210     m0026(.A0(mai_mai_n54_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NA3        m0031(.A(g), .B(mai_mai_n59_), .C(a), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(h), .Y(mai_mai_n61_));
  NAi31      m0033(.An(i), .B(l), .C(j), .Y(mai_mai_n62_));
  OAI220     m0034(.A0(mai_mai_n62_), .A1(mai_mai_n49_), .B0(mai_mai_n61_), .B1(mai_mai_n44_), .Y(mai_mai_n63_));
  NAi31      m0035(.An(mai_mai_n60_), .B(mai_mai_n63_), .C(mai_mai_n58_), .Y(mai_mai_n64_));
  NAi41      m0036(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n65_));
  NA2        m0037(.A(g), .B(f), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi21      m0039(.An(i), .B(j), .Y(mai_mai_n68_));
  NAi32      m0040(.An(n), .Bn(k), .C(m), .Y(mai_mai_n69_));
  NO2        m0041(.A(mai_mai_n69_), .B(mai_mai_n68_), .Y(mai_mai_n70_));
  NAi31      m0042(.An(l), .B(m), .C(k), .Y(mai_mai_n71_));
  NAi21      m0043(.An(e), .B(h), .Y(mai_mai_n72_));
  NAi41      m0044(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n74_));
  INV        m0046(.A(m), .Y(mai_mai_n75_));
  NOi21      m0047(.An(k), .B(l), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n77_));
  AN4        m0049(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n78_));
  NOi31      m0050(.An(h), .B(g), .C(f), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  NAi32      m0052(.An(m), .Bn(k), .C(j), .Y(mai_mai_n81_));
  NOi32      m0053(.An(h), .Bn(g), .C(f), .Y(mai_mai_n82_));
  NA2        m0054(.A(mai_mai_n82_), .B(mai_mai_n78_), .Y(mai_mai_n83_));
  OA220      m0055(.A0(mai_mai_n83_), .A1(mai_mai_n81_), .B0(mai_mai_n80_), .B1(mai_mai_n77_), .Y(mai_mai_n84_));
  NA3        m0056(.A(mai_mai_n84_), .B(mai_mai_n74_), .C(mai_mai_n64_), .Y(mai_mai_n85_));
  INV        m0057(.A(n), .Y(mai_mai_n86_));
  NOi32      m0058(.An(e), .Bn(b), .C(d), .Y(mai_mai_n87_));
  NA2        m0059(.A(mai_mai_n87_), .B(mai_mai_n86_), .Y(mai_mai_n88_));
  INV        m0060(.A(j), .Y(mai_mai_n89_));
  AN3        m0061(.A(m), .B(k), .C(i), .Y(mai_mai_n90_));
  NA3        m0062(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(g), .Y(mai_mai_n91_));
  NAi32      m0063(.An(g), .Bn(f), .C(h), .Y(mai_mai_n92_));
  NAi31      m0064(.An(j), .B(m), .C(l), .Y(mai_mai_n93_));
  NA2        m0065(.A(m), .B(l), .Y(mai_mai_n94_));
  NAi31      m0066(.An(k), .B(j), .C(g), .Y(mai_mai_n95_));
  NO3        m0067(.A(mai_mai_n95_), .B(mai_mai_n94_), .C(f), .Y(mai_mai_n96_));
  AN2        m0068(.A(j), .B(g), .Y(mai_mai_n97_));
  NOi32      m0069(.An(m), .Bn(l), .C(i), .Y(mai_mai_n98_));
  NOi21      m0070(.An(g), .B(i), .Y(mai_mai_n99_));
  NOi32      m0071(.An(m), .Bn(j), .C(k), .Y(mai_mai_n100_));
  AOI220     m0072(.A0(mai_mai_n100_), .A1(mai_mai_n99_), .B0(mai_mai_n98_), .B1(mai_mai_n97_), .Y(mai_mai_n101_));
  NO2        m0073(.A(mai_mai_n101_), .B(f), .Y(mai_mai_n102_));
  NAi41      m0074(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n103_));
  AN2        m0075(.A(e), .B(b), .Y(mai_mai_n104_));
  NOi31      m0076(.An(c), .B(h), .C(f), .Y(mai_mai_n105_));
  NA2        m0077(.A(mai_mai_n105_), .B(mai_mai_n104_), .Y(mai_mai_n106_));
  NO3        m0078(.A(mai_mai_n106_), .B(mai_mai_n103_), .C(g), .Y(mai_mai_n107_));
  NOi21      m0079(.An(g), .B(f), .Y(mai_mai_n108_));
  NOi21      m0080(.An(i), .B(h), .Y(mai_mai_n109_));
  NA3        m0081(.A(mai_mai_n109_), .B(mai_mai_n108_), .C(mai_mai_n36_), .Y(mai_mai_n110_));
  INV        m0082(.A(a), .Y(mai_mai_n111_));
  NA2        m0083(.A(mai_mai_n104_), .B(mai_mai_n111_), .Y(mai_mai_n112_));
  INV        m0084(.A(l), .Y(mai_mai_n113_));
  NOi21      m0085(.An(m), .B(n), .Y(mai_mai_n114_));
  AN2        m0086(.A(k), .B(h), .Y(mai_mai_n115_));
  NO2        m0087(.A(mai_mai_n110_), .B(mai_mai_n88_), .Y(mai_mai_n116_));
  INV        m0088(.A(b), .Y(mai_mai_n117_));
  NA2        m0089(.A(l), .B(j), .Y(mai_mai_n118_));
  AN2        m0090(.A(k), .B(i), .Y(mai_mai_n119_));
  NA2        m0091(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n120_));
  NA2        m0092(.A(g), .B(e), .Y(mai_mai_n121_));
  NOi32      m0093(.An(c), .Bn(a), .C(d), .Y(mai_mai_n122_));
  NA2        m0094(.A(mai_mai_n122_), .B(mai_mai_n114_), .Y(mai_mai_n123_));
  NO4        m0095(.A(mai_mai_n123_), .B(mai_mai_n121_), .C(mai_mai_n120_), .D(mai_mai_n117_), .Y(mai_mai_n124_));
  NO3        m0096(.A(mai_mai_n124_), .B(mai_mai_n116_), .C(mai_mai_n107_), .Y(mai_mai_n125_));
  OAI210     m0097(.A0(mai_mai_n101_), .A1(mai_mai_n88_), .B0(mai_mai_n125_), .Y(mai_mai_n126_));
  NOi31      m0098(.An(k), .B(m), .C(j), .Y(mai_mai_n127_));
  NOi31      m0099(.An(k), .B(m), .C(i), .Y(mai_mai_n128_));
  NA3        m0100(.A(mai_mai_n128_), .B(mai_mai_n82_), .C(mai_mai_n78_), .Y(mai_mai_n129_));
  INV        m0101(.A(mai_mai_n129_), .Y(mai_mai_n130_));
  NOi32      m0102(.An(f), .Bn(b), .C(e), .Y(mai_mai_n131_));
  NAi21      m0103(.An(g), .B(h), .Y(mai_mai_n132_));
  NAi21      m0104(.An(m), .B(n), .Y(mai_mai_n133_));
  NAi21      m0105(.An(j), .B(k), .Y(mai_mai_n134_));
  NAi41      m0106(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n135_));
  NAi31      m0107(.An(j), .B(k), .C(h), .Y(mai_mai_n136_));
  NO3        m0108(.A(mai_mai_n136_), .B(mai_mai_n135_), .C(mai_mai_n133_), .Y(mai_mai_n137_));
  INV        m0109(.A(mai_mai_n137_), .Y(mai_mai_n138_));
  NO2        m0110(.A(k), .B(j), .Y(mai_mai_n139_));
  AN2        m0111(.A(k), .B(j), .Y(mai_mai_n140_));
  NAi21      m0112(.An(c), .B(b), .Y(mai_mai_n141_));
  NA2        m0113(.A(f), .B(d), .Y(mai_mai_n142_));
  NA2        m0114(.A(h), .B(c), .Y(mai_mai_n143_));
  NAi31      m0115(.An(f), .B(e), .C(b), .Y(mai_mai_n144_));
  NA2        m0116(.A(d), .B(b), .Y(mai_mai_n145_));
  NAi21      m0117(.An(e), .B(f), .Y(mai_mai_n146_));
  NO2        m0118(.A(mai_mai_n146_), .B(mai_mai_n145_), .Y(mai_mai_n147_));
  NA2        m0119(.A(b), .B(a), .Y(mai_mai_n148_));
  NAi21      m0120(.An(e), .B(g), .Y(mai_mai_n149_));
  NAi21      m0121(.An(c), .B(d), .Y(mai_mai_n150_));
  NAi31      m0122(.An(l), .B(k), .C(h), .Y(mai_mai_n151_));
  NO2        m0123(.A(mai_mai_n133_), .B(mai_mai_n151_), .Y(mai_mai_n152_));
  NAi21      m0124(.An(mai_mai_n130_), .B(mai_mai_n138_), .Y(mai_mai_n153_));
  NAi31      m0125(.An(e), .B(f), .C(b), .Y(mai_mai_n154_));
  NOi21      m0126(.An(g), .B(d), .Y(mai_mai_n155_));
  NO2        m0127(.A(mai_mai_n155_), .B(mai_mai_n154_), .Y(mai_mai_n156_));
  NOi21      m0128(.An(h), .B(i), .Y(mai_mai_n157_));
  NOi21      m0129(.An(k), .B(m), .Y(mai_mai_n158_));
  NA3        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .C(n), .Y(mai_mai_n159_));
  NOi21      m0131(.An(mai_mai_n156_), .B(mai_mai_n159_), .Y(mai_mai_n160_));
  NOi21      m0132(.An(h), .B(g), .Y(mai_mai_n161_));
  NO2        m0133(.A(mai_mai_n142_), .B(mai_mai_n141_), .Y(mai_mai_n162_));
  NA2        m0134(.A(mai_mai_n162_), .B(mai_mai_n161_), .Y(mai_mai_n163_));
  NAi31      m0135(.An(l), .B(j), .C(h), .Y(mai_mai_n164_));
  NO2        m0136(.A(mai_mai_n164_), .B(mai_mai_n49_), .Y(mai_mai_n165_));
  NA2        m0137(.A(mai_mai_n165_), .B(mai_mai_n67_), .Y(mai_mai_n166_));
  NOi32      m0138(.An(n), .Bn(k), .C(m), .Y(mai_mai_n167_));
  NA2        m0139(.A(l), .B(i), .Y(mai_mai_n168_));
  NA2        m0140(.A(mai_mai_n168_), .B(mai_mai_n167_), .Y(mai_mai_n169_));
  OAI210     m0141(.A0(mai_mai_n169_), .A1(mai_mai_n163_), .B0(mai_mai_n166_), .Y(mai_mai_n170_));
  NAi31      m0142(.An(d), .B(f), .C(c), .Y(mai_mai_n171_));
  NAi31      m0143(.An(e), .B(f), .C(c), .Y(mai_mai_n172_));
  NA2        m0144(.A(mai_mai_n172_), .B(mai_mai_n171_), .Y(mai_mai_n173_));
  NA2        m0145(.A(j), .B(h), .Y(mai_mai_n174_));
  OR3        m0146(.A(n), .B(m), .C(k), .Y(mai_mai_n175_));
  NO2        m0147(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  NAi32      m0148(.An(m), .Bn(k), .C(n), .Y(mai_mai_n177_));
  NO2        m0149(.A(mai_mai_n177_), .B(mai_mai_n174_), .Y(mai_mai_n178_));
  AOI220     m0150(.A0(mai_mai_n178_), .A1(mai_mai_n156_), .B0(mai_mai_n176_), .B1(mai_mai_n173_), .Y(mai_mai_n179_));
  NO2        m0151(.A(n), .B(m), .Y(mai_mai_n180_));
  NA2        m0152(.A(mai_mai_n180_), .B(mai_mai_n50_), .Y(mai_mai_n181_));
  NAi21      m0153(.An(f), .B(e), .Y(mai_mai_n182_));
  NA2        m0154(.A(d), .B(c), .Y(mai_mai_n183_));
  NAi21      m0155(.An(d), .B(c), .Y(mai_mai_n184_));
  NAi31      m0156(.An(m), .B(n), .C(b), .Y(mai_mai_n185_));
  NA2        m0157(.A(k), .B(i), .Y(mai_mai_n186_));
  NAi21      m0158(.An(h), .B(f), .Y(mai_mai_n187_));
  NO2        m0159(.A(mai_mai_n187_), .B(mai_mai_n186_), .Y(mai_mai_n188_));
  NO2        m0160(.A(mai_mai_n185_), .B(mai_mai_n150_), .Y(mai_mai_n189_));
  NA2        m0161(.A(mai_mai_n189_), .B(mai_mai_n188_), .Y(mai_mai_n190_));
  NOi32      m0162(.An(f), .Bn(c), .C(d), .Y(mai_mai_n191_));
  NOi32      m0163(.An(f), .Bn(c), .C(e), .Y(mai_mai_n192_));
  NO2        m0164(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n193_));
  NO3        m0165(.A(n), .B(m), .C(j), .Y(mai_mai_n194_));
  NA2        m0166(.A(mai_mai_n194_), .B(mai_mai_n115_), .Y(mai_mai_n195_));
  AO210      m0167(.A0(mai_mai_n195_), .A1(mai_mai_n181_), .B0(mai_mai_n193_), .Y(mai_mai_n196_));
  NA3        m0168(.A(mai_mai_n196_), .B(mai_mai_n190_), .C(mai_mai_n179_), .Y(mai_mai_n197_));
  OR4        m0169(.A(mai_mai_n197_), .B(mai_mai_n170_), .C(mai_mai_n160_), .D(mai_mai_n153_), .Y(mai_mai_n198_));
  NO4        m0170(.A(mai_mai_n198_), .B(mai_mai_n126_), .C(mai_mai_n85_), .D(mai_mai_n55_), .Y(mai_mai_n199_));
  NA3        m0171(.A(m), .B(mai_mai_n113_), .C(j), .Y(mai_mai_n200_));
  NAi31      m0172(.An(n), .B(h), .C(g), .Y(mai_mai_n201_));
  NO2        m0173(.A(mai_mai_n201_), .B(mai_mai_n200_), .Y(mai_mai_n202_));
  NOi32      m0174(.An(m), .Bn(k), .C(l), .Y(mai_mai_n203_));
  NA3        m0175(.A(mai_mai_n203_), .B(mai_mai_n89_), .C(g), .Y(mai_mai_n204_));
  NO2        m0176(.A(mai_mai_n204_), .B(n), .Y(mai_mai_n205_));
  NOi21      m0177(.An(k), .B(j), .Y(mai_mai_n206_));
  NA4        m0178(.A(mai_mai_n206_), .B(mai_mai_n114_), .C(i), .D(g), .Y(mai_mai_n207_));
  AN2        m0179(.A(i), .B(g), .Y(mai_mai_n208_));
  NA3        m0180(.A(mai_mai_n76_), .B(mai_mai_n208_), .C(mai_mai_n114_), .Y(mai_mai_n209_));
  NA2        m0181(.A(mai_mai_n209_), .B(mai_mai_n207_), .Y(mai_mai_n210_));
  NO3        m0182(.A(mai_mai_n210_), .B(mai_mai_n205_), .C(mai_mai_n202_), .Y(mai_mai_n211_));
  NAi41      m0183(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n212_));
  INV        m0184(.A(mai_mai_n212_), .Y(mai_mai_n213_));
  INV        m0185(.A(f), .Y(mai_mai_n214_));
  INV        m0186(.A(g), .Y(mai_mai_n215_));
  NOi31      m0187(.An(i), .B(j), .C(h), .Y(mai_mai_n216_));
  NOi21      m0188(.An(l), .B(m), .Y(mai_mai_n217_));
  NA2        m0189(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  NO2        m0190(.A(mai_mai_n211_), .B(mai_mai_n32_), .Y(mai_mai_n219_));
  NOi21      m0191(.An(n), .B(m), .Y(mai_mai_n220_));
  NOi32      m0192(.An(l), .Bn(i), .C(j), .Y(mai_mai_n221_));
  NA2        m0193(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n222_));
  OA220      m0194(.A0(mai_mai_n222_), .A1(mai_mai_n106_), .B0(mai_mai_n81_), .B1(mai_mai_n80_), .Y(mai_mai_n223_));
  NAi21      m0195(.An(j), .B(h), .Y(mai_mai_n224_));
  XN2        m0196(.A(i), .B(h), .Y(mai_mai_n225_));
  NA2        m0197(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n226_));
  NOi31      m0198(.An(k), .B(n), .C(m), .Y(mai_mai_n227_));
  NOi31      m0199(.An(mai_mai_n227_), .B(mai_mai_n183_), .C(mai_mai_n182_), .Y(mai_mai_n228_));
  NA2        m0200(.A(mai_mai_n228_), .B(mai_mai_n226_), .Y(mai_mai_n229_));
  NAi31      m0201(.An(f), .B(e), .C(c), .Y(mai_mai_n230_));
  NO4        m0202(.A(mai_mai_n230_), .B(mai_mai_n175_), .C(mai_mai_n174_), .D(mai_mai_n59_), .Y(mai_mai_n231_));
  NA4        m0203(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n232_));
  NAi32      m0204(.An(m), .Bn(i), .C(k), .Y(mai_mai_n233_));
  NO3        m0205(.A(mai_mai_n233_), .B(mai_mai_n92_), .C(mai_mai_n232_), .Y(mai_mai_n234_));
  NA2        m0206(.A(k), .B(h), .Y(mai_mai_n235_));
  NO2        m0207(.A(mai_mai_n234_), .B(mai_mai_n231_), .Y(mai_mai_n236_));
  NAi21      m0208(.An(n), .B(a), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n237_), .B(mai_mai_n145_), .Y(mai_mai_n238_));
  NAi41      m0210(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n239_));
  NO2        m0211(.A(mai_mai_n239_), .B(e), .Y(mai_mai_n240_));
  NO3        m0212(.A(mai_mai_n146_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n241_));
  OAI210     m0213(.A0(mai_mai_n241_), .A1(mai_mai_n240_), .B0(mai_mai_n238_), .Y(mai_mai_n242_));
  AN4        m0214(.A(mai_mai_n242_), .B(mai_mai_n236_), .C(mai_mai_n229_), .D(mai_mai_n223_), .Y(mai_mai_n243_));
  OR2        m0215(.A(h), .B(g), .Y(mai_mai_n244_));
  NO2        m0216(.A(mai_mai_n244_), .B(mai_mai_n103_), .Y(mai_mai_n245_));
  NA2        m0217(.A(mai_mai_n245_), .B(mai_mai_n131_), .Y(mai_mai_n246_));
  NAi41      m0218(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n247_));
  NO2        m0219(.A(mai_mai_n247_), .B(mai_mai_n214_), .Y(mai_mai_n248_));
  NA2        m0220(.A(mai_mai_n158_), .B(mai_mai_n109_), .Y(mai_mai_n249_));
  NO2        m0221(.A(n), .B(a), .Y(mai_mai_n250_));
  NAi31      m0222(.An(mai_mai_n239_), .B(mai_mai_n250_), .C(mai_mai_n104_), .Y(mai_mai_n251_));
  NAi21      m0223(.An(h), .B(i), .Y(mai_mai_n252_));
  NA2        m0224(.A(mai_mai_n180_), .B(k), .Y(mai_mai_n253_));
  NO2        m0225(.A(mai_mai_n253_), .B(mai_mai_n252_), .Y(mai_mai_n254_));
  NA2        m0226(.A(mai_mai_n254_), .B(mai_mai_n191_), .Y(mai_mai_n255_));
  NA3        m0227(.A(mai_mai_n255_), .B(mai_mai_n251_), .C(mai_mai_n246_), .Y(mai_mai_n256_));
  NOi21      m0228(.An(g), .B(e), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n258_), .B(mai_mai_n257_), .Y(mai_mai_n259_));
  NOi32      m0231(.An(l), .Bn(j), .C(i), .Y(mai_mai_n260_));
  AOI210     m0232(.A0(mai_mai_n76_), .A1(mai_mai_n89_), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  NO2        m0233(.A(mai_mai_n252_), .B(mai_mai_n44_), .Y(mai_mai_n262_));
  NAi21      m0234(.An(f), .B(g), .Y(mai_mai_n263_));
  NO2        m0235(.A(mai_mai_n263_), .B(mai_mai_n65_), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n69_), .B(mai_mai_n118_), .Y(mai_mai_n265_));
  AOI220     m0237(.A0(mai_mai_n265_), .A1(mai_mai_n264_), .B0(mai_mai_n262_), .B1(mai_mai_n67_), .Y(mai_mai_n266_));
  OAI210     m0238(.A0(mai_mai_n261_), .A1(mai_mai_n259_), .B0(mai_mai_n266_), .Y(mai_mai_n267_));
  NO3        m0239(.A(mai_mai_n134_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n268_));
  NOi41      m0240(.An(mai_mai_n243_), .B(mai_mai_n267_), .C(mai_mai_n256_), .D(mai_mai_n219_), .Y(mai_mai_n269_));
  NO4        m0241(.A(mai_mai_n202_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n270_));
  NO2        m0242(.A(mai_mai_n270_), .B(mai_mai_n112_), .Y(mai_mai_n271_));
  NA3        m0243(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n272_));
  NAi21      m0244(.An(h), .B(g), .Y(mai_mai_n273_));
  OR4        m0245(.A(mai_mai_n273_), .B(mai_mai_n272_), .C(mai_mai_n222_), .D(e), .Y(mai_mai_n274_));
  NAi31      m0246(.An(g), .B(k), .C(h), .Y(mai_mai_n275_));
  NO3        m0247(.A(mai_mai_n133_), .B(mai_mai_n275_), .C(l), .Y(mai_mai_n276_));
  NAi31      m0248(.An(e), .B(d), .C(a), .Y(mai_mai_n277_));
  NA2        m0249(.A(mai_mai_n276_), .B(mai_mai_n131_), .Y(mai_mai_n278_));
  NA2        m0250(.A(mai_mai_n278_), .B(mai_mai_n274_), .Y(mai_mai_n279_));
  NA3        m0251(.A(mai_mai_n158_), .B(mai_mai_n157_), .C(mai_mai_n86_), .Y(mai_mai_n280_));
  NO2        m0252(.A(mai_mai_n280_), .B(mai_mai_n193_), .Y(mai_mai_n281_));
  INV        m0253(.A(mai_mai_n281_), .Y(mai_mai_n282_));
  NA3        m0254(.A(e), .B(c), .C(b), .Y(mai_mai_n283_));
  NO2        m0255(.A(mai_mai_n60_), .B(mai_mai_n283_), .Y(mai_mai_n284_));
  NAi32      m0256(.An(k), .Bn(i), .C(j), .Y(mai_mai_n285_));
  NAi31      m0257(.An(h), .B(l), .C(i), .Y(mai_mai_n286_));
  NA3        m0258(.A(mai_mai_n286_), .B(mai_mai_n285_), .C(mai_mai_n164_), .Y(mai_mai_n287_));
  NOi21      m0259(.An(mai_mai_n287_), .B(mai_mai_n49_), .Y(mai_mai_n288_));
  OAI210     m0260(.A0(mai_mai_n264_), .A1(mai_mai_n284_), .B0(mai_mai_n288_), .Y(mai_mai_n289_));
  NAi21      m0261(.An(l), .B(k), .Y(mai_mai_n290_));
  NO2        m0262(.A(mai_mai_n290_), .B(mai_mai_n49_), .Y(mai_mai_n291_));
  NOi21      m0263(.An(l), .B(j), .Y(mai_mai_n292_));
  NA2        m0264(.A(mai_mai_n161_), .B(mai_mai_n292_), .Y(mai_mai_n293_));
  NA3        m0265(.A(mai_mai_n119_), .B(mai_mai_n118_), .C(g), .Y(mai_mai_n294_));
  OR3        m0266(.A(mai_mai_n73_), .B(mai_mai_n75_), .C(e), .Y(mai_mai_n295_));
  AOI210     m0267(.A0(mai_mai_n294_), .A1(mai_mai_n293_), .B0(mai_mai_n295_), .Y(mai_mai_n296_));
  INV        m0268(.A(mai_mai_n296_), .Y(mai_mai_n297_));
  NAi32      m0269(.An(j), .Bn(h), .C(i), .Y(mai_mai_n298_));
  NAi21      m0270(.An(m), .B(l), .Y(mai_mai_n299_));
  NO3        m0271(.A(mai_mai_n299_), .B(mai_mai_n298_), .C(mai_mai_n86_), .Y(mai_mai_n300_));
  NA2        m0272(.A(h), .B(g), .Y(mai_mai_n301_));
  NA2        m0273(.A(mai_mai_n167_), .B(mai_mai_n45_), .Y(mai_mai_n302_));
  NO2        m0274(.A(mai_mai_n302_), .B(mai_mai_n301_), .Y(mai_mai_n303_));
  OAI210     m0275(.A0(mai_mai_n303_), .A1(mai_mai_n300_), .B0(mai_mai_n162_), .Y(mai_mai_n304_));
  NA4        m0276(.A(mai_mai_n304_), .B(mai_mai_n297_), .C(mai_mai_n289_), .D(mai_mai_n282_), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n144_), .B(d), .Y(mai_mai_n306_));
  NA2        m0278(.A(mai_mai_n306_), .B(mai_mai_n53_), .Y(mai_mai_n307_));
  NO2        m0279(.A(mai_mai_n106_), .B(mai_mai_n103_), .Y(mai_mai_n308_));
  NAi32      m0280(.An(n), .Bn(m), .C(l), .Y(mai_mai_n309_));
  NO2        m0281(.A(mai_mai_n309_), .B(mai_mai_n298_), .Y(mai_mai_n310_));
  NO2        m0282(.A(mai_mai_n123_), .B(mai_mai_n117_), .Y(mai_mai_n311_));
  NAi31      m0283(.An(k), .B(l), .C(j), .Y(mai_mai_n312_));
  OAI210     m0284(.A0(mai_mai_n290_), .A1(j), .B0(mai_mai_n312_), .Y(mai_mai_n313_));
  NOi21      m0285(.An(mai_mai_n313_), .B(mai_mai_n121_), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n314_), .B(mai_mai_n311_), .Y(mai_mai_n315_));
  NA2        m0287(.A(mai_mai_n315_), .B(mai_mai_n307_), .Y(mai_mai_n316_));
  NO4        m0288(.A(mai_mai_n316_), .B(mai_mai_n305_), .C(mai_mai_n279_), .D(mai_mai_n271_), .Y(mai_mai_n317_));
  NA2        m0289(.A(mai_mai_n254_), .B(mai_mai_n192_), .Y(mai_mai_n318_));
  NAi21      m0290(.An(m), .B(k), .Y(mai_mai_n319_));
  NO2        m0291(.A(mai_mai_n225_), .B(mai_mai_n319_), .Y(mai_mai_n320_));
  NAi41      m0292(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n321_));
  NO2        m0293(.A(mai_mai_n321_), .B(mai_mai_n149_), .Y(mai_mai_n322_));
  NA2        m0294(.A(mai_mai_n322_), .B(mai_mai_n320_), .Y(mai_mai_n323_));
  NAi31      m0295(.An(i), .B(l), .C(h), .Y(mai_mai_n324_));
  NO4        m0296(.A(mai_mai_n324_), .B(mai_mai_n149_), .C(mai_mai_n73_), .D(mai_mai_n75_), .Y(mai_mai_n325_));
  NA2        m0297(.A(e), .B(c), .Y(mai_mai_n326_));
  NO3        m0298(.A(mai_mai_n326_), .B(n), .C(d), .Y(mai_mai_n327_));
  NOi21      m0299(.An(f), .B(h), .Y(mai_mai_n328_));
  NA2        m0300(.A(mai_mai_n328_), .B(mai_mai_n119_), .Y(mai_mai_n329_));
  NO2        m0301(.A(mai_mai_n329_), .B(mai_mai_n215_), .Y(mai_mai_n330_));
  NAi31      m0302(.An(d), .B(e), .C(b), .Y(mai_mai_n331_));
  NO2        m0303(.A(mai_mai_n133_), .B(mai_mai_n331_), .Y(mai_mai_n332_));
  NA2        m0304(.A(mai_mai_n332_), .B(mai_mai_n330_), .Y(mai_mai_n333_));
  NAi41      m0305(.An(mai_mai_n325_), .B(mai_mai_n333_), .C(mai_mai_n323_), .D(mai_mai_n318_), .Y(mai_mai_n334_));
  NO4        m0306(.A(mai_mai_n321_), .B(mai_mai_n81_), .C(mai_mai_n72_), .D(mai_mai_n215_), .Y(mai_mai_n335_));
  NA2        m0307(.A(mai_mai_n250_), .B(mai_mai_n104_), .Y(mai_mai_n336_));
  OR2        m0308(.A(mai_mai_n336_), .B(mai_mai_n204_), .Y(mai_mai_n337_));
  NOi31      m0309(.An(l), .B(n), .C(m), .Y(mai_mai_n338_));
  NA2        m0310(.A(mai_mai_n338_), .B(mai_mai_n216_), .Y(mai_mai_n339_));
  NO2        m0311(.A(mai_mai_n339_), .B(mai_mai_n193_), .Y(mai_mai_n340_));
  NAi32      m0312(.An(mai_mai_n340_), .Bn(mai_mai_n335_), .C(mai_mai_n337_), .Y(mai_mai_n341_));
  NAi32      m0313(.An(m), .Bn(j), .C(k), .Y(mai_mai_n342_));
  NAi41      m0314(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n343_));
  NOi31      m0315(.An(j), .B(m), .C(k), .Y(mai_mai_n344_));
  NO2        m0316(.A(mai_mai_n127_), .B(mai_mai_n344_), .Y(mai_mai_n345_));
  AN3        m0317(.A(h), .B(g), .C(f), .Y(mai_mai_n346_));
  NOi32      m0318(.An(m), .Bn(j), .C(l), .Y(mai_mai_n347_));
  NO2        m0319(.A(mai_mai_n347_), .B(mai_mai_n98_), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n299_), .B(mai_mai_n298_), .Y(mai_mai_n349_));
  NO2        m0321(.A(mai_mai_n218_), .B(g), .Y(mai_mai_n350_));
  NA2        m0322(.A(mai_mai_n233_), .B(mai_mai_n81_), .Y(mai_mai_n351_));
  NA3        m0323(.A(mai_mai_n351_), .B(mai_mai_n346_), .C(mai_mai_n213_), .Y(mai_mai_n352_));
  INV        m0324(.A(mai_mai_n352_), .Y(mai_mai_n353_));
  NA3        m0325(.A(h), .B(g), .C(f), .Y(mai_mai_n354_));
  NO2        m0326(.A(mai_mai_n354_), .B(mai_mai_n77_), .Y(mai_mai_n355_));
  NA2        m0327(.A(mai_mai_n343_), .B(mai_mai_n212_), .Y(mai_mai_n356_));
  NA2        m0328(.A(mai_mai_n161_), .B(e), .Y(mai_mai_n357_));
  NO2        m0329(.A(mai_mai_n357_), .B(mai_mai_n41_), .Y(mai_mai_n358_));
  AOI220     m0330(.A0(mai_mai_n358_), .A1(mai_mai_n311_), .B0(mai_mai_n356_), .B1(mai_mai_n355_), .Y(mai_mai_n359_));
  NOi32      m0331(.An(j), .Bn(g), .C(i), .Y(mai_mai_n360_));
  NA3        m0332(.A(mai_mai_n360_), .B(mai_mai_n290_), .C(mai_mai_n114_), .Y(mai_mai_n361_));
  AO210      m0333(.A0(mai_mai_n112_), .A1(mai_mai_n32_), .B0(mai_mai_n361_), .Y(mai_mai_n362_));
  NOi32      m0334(.An(e), .Bn(b), .C(a), .Y(mai_mai_n363_));
  AN2        m0335(.A(l), .B(j), .Y(mai_mai_n364_));
  NO2        m0336(.A(mai_mai_n319_), .B(mai_mai_n364_), .Y(mai_mai_n365_));
  NO3        m0337(.A(mai_mai_n321_), .B(mai_mai_n72_), .C(mai_mai_n215_), .Y(mai_mai_n366_));
  NA3        m0338(.A(mai_mai_n209_), .B(mai_mai_n207_), .C(mai_mai_n35_), .Y(mai_mai_n367_));
  AOI220     m0339(.A0(mai_mai_n367_), .A1(mai_mai_n363_), .B0(mai_mai_n366_), .B1(mai_mai_n365_), .Y(mai_mai_n368_));
  NO2        m0340(.A(mai_mai_n331_), .B(n), .Y(mai_mai_n369_));
  NA2        m0341(.A(mai_mai_n208_), .B(k), .Y(mai_mai_n370_));
  NA3        m0342(.A(m), .B(mai_mai_n113_), .C(mai_mai_n214_), .Y(mai_mai_n371_));
  NA4        m0343(.A(mai_mai_n203_), .B(mai_mai_n89_), .C(g), .D(mai_mai_n214_), .Y(mai_mai_n372_));
  OAI210     m0344(.A0(mai_mai_n371_), .A1(mai_mai_n370_), .B0(mai_mai_n372_), .Y(mai_mai_n373_));
  NAi41      m0345(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n374_));
  NA2        m0346(.A(mai_mai_n51_), .B(mai_mai_n114_), .Y(mai_mai_n375_));
  NO2        m0347(.A(mai_mai_n375_), .B(mai_mai_n374_), .Y(mai_mai_n376_));
  AOI220     m0348(.A0(mai_mai_n376_), .A1(b), .B0(mai_mai_n373_), .B1(mai_mai_n369_), .Y(mai_mai_n377_));
  NA4        m0349(.A(mai_mai_n377_), .B(mai_mai_n368_), .C(mai_mai_n362_), .D(mai_mai_n359_), .Y(mai_mai_n378_));
  NO4        m0350(.A(mai_mai_n378_), .B(mai_mai_n353_), .C(mai_mai_n341_), .D(mai_mai_n334_), .Y(mai_mai_n379_));
  NA4        m0351(.A(mai_mai_n379_), .B(mai_mai_n317_), .C(mai_mai_n269_), .D(mai_mai_n199_), .Y(mai10));
  NA3        m0352(.A(m), .B(k), .C(i), .Y(mai_mai_n381_));
  NO3        m0353(.A(mai_mai_n381_), .B(j), .C(mai_mai_n215_), .Y(mai_mai_n382_));
  NOi21      m0354(.An(e), .B(f), .Y(mai_mai_n383_));
  NO4        m0355(.A(mai_mai_n150_), .B(mai_mai_n383_), .C(n), .D(mai_mai_n111_), .Y(mai_mai_n384_));
  NAi31      m0356(.An(b), .B(f), .C(c), .Y(mai_mai_n385_));
  INV        m0357(.A(mai_mai_n385_), .Y(mai_mai_n386_));
  NOi32      m0358(.An(k), .Bn(h), .C(j), .Y(mai_mai_n387_));
  NA2        m0359(.A(mai_mai_n387_), .B(mai_mai_n220_), .Y(mai_mai_n388_));
  NA2        m0360(.A(mai_mai_n159_), .B(mai_mai_n388_), .Y(mai_mai_n389_));
  AOI220     m0361(.A0(mai_mai_n389_), .A1(mai_mai_n386_), .B0(mai_mai_n384_), .B1(mai_mai_n382_), .Y(mai_mai_n390_));
  AN2        m0362(.A(j), .B(h), .Y(mai_mai_n391_));
  NO3        m0363(.A(n), .B(m), .C(k), .Y(mai_mai_n392_));
  NA2        m0364(.A(mai_mai_n392_), .B(mai_mai_n391_), .Y(mai_mai_n393_));
  NO3        m0365(.A(mai_mai_n393_), .B(mai_mai_n150_), .C(mai_mai_n214_), .Y(mai_mai_n394_));
  OR2        m0366(.A(m), .B(k), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n174_), .B(mai_mai_n395_), .Y(mai_mai_n396_));
  NA4        m0368(.A(n), .B(f), .C(c), .D(mai_mai_n117_), .Y(mai_mai_n397_));
  NOi21      m0369(.An(mai_mai_n396_), .B(mai_mai_n397_), .Y(mai_mai_n398_));
  NOi32      m0370(.An(d), .Bn(a), .C(c), .Y(mai_mai_n399_));
  NA2        m0371(.A(mai_mai_n399_), .B(mai_mai_n182_), .Y(mai_mai_n400_));
  NAi21      m0372(.An(i), .B(g), .Y(mai_mai_n401_));
  NAi31      m0373(.An(k), .B(m), .C(j), .Y(mai_mai_n402_));
  NO3        m0374(.A(mai_mai_n402_), .B(mai_mai_n401_), .C(n), .Y(mai_mai_n403_));
  NOi21      m0375(.An(mai_mai_n403_), .B(mai_mai_n400_), .Y(mai_mai_n404_));
  NO3        m0376(.A(mai_mai_n404_), .B(mai_mai_n398_), .C(mai_mai_n394_), .Y(mai_mai_n405_));
  NO2        m0377(.A(mai_mai_n397_), .B(mai_mai_n299_), .Y(mai_mai_n406_));
  NOi32      m0378(.An(f), .Bn(d), .C(c), .Y(mai_mai_n407_));
  AOI220     m0379(.A0(mai_mai_n407_), .A1(mai_mai_n310_), .B0(mai_mai_n406_), .B1(mai_mai_n216_), .Y(mai_mai_n408_));
  NA3        m0380(.A(mai_mai_n408_), .B(mai_mai_n405_), .C(mai_mai_n390_), .Y(mai_mai_n409_));
  NO2        m0381(.A(mai_mai_n59_), .B(mai_mai_n117_), .Y(mai_mai_n410_));
  NA2        m0382(.A(mai_mai_n250_), .B(mai_mai_n410_), .Y(mai_mai_n411_));
  INV        m0383(.A(e), .Y(mai_mai_n412_));
  NA2        m0384(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n413_));
  OAI220     m0385(.A0(mai_mai_n413_), .A1(mai_mai_n200_), .B0(mai_mai_n204_), .B1(mai_mai_n412_), .Y(mai_mai_n414_));
  AN2        m0386(.A(g), .B(e), .Y(mai_mai_n415_));
  NA3        m0387(.A(mai_mai_n415_), .B(mai_mai_n203_), .C(i), .Y(mai_mai_n416_));
  OAI210     m0388(.A0(mai_mai_n91_), .A1(mai_mai_n412_), .B0(mai_mai_n416_), .Y(mai_mai_n417_));
  NO2        m0389(.A(mai_mai_n101_), .B(mai_mai_n412_), .Y(mai_mai_n418_));
  NO3        m0390(.A(mai_mai_n418_), .B(mai_mai_n417_), .C(mai_mai_n414_), .Y(mai_mai_n419_));
  NOi32      m0391(.An(h), .Bn(e), .C(g), .Y(mai_mai_n420_));
  NA3        m0392(.A(mai_mai_n420_), .B(mai_mai_n292_), .C(m), .Y(mai_mai_n421_));
  NOi21      m0393(.An(g), .B(h), .Y(mai_mai_n422_));
  AN3        m0394(.A(m), .B(l), .C(i), .Y(mai_mai_n423_));
  NA3        m0395(.A(mai_mai_n423_), .B(mai_mai_n422_), .C(e), .Y(mai_mai_n424_));
  AN3        m0396(.A(h), .B(g), .C(e), .Y(mai_mai_n425_));
  NA2        m0397(.A(mai_mai_n425_), .B(mai_mai_n98_), .Y(mai_mai_n426_));
  AN3        m0398(.A(mai_mai_n426_), .B(mai_mai_n424_), .C(mai_mai_n421_), .Y(mai_mai_n427_));
  AOI210     m0399(.A0(mai_mai_n427_), .A1(mai_mai_n419_), .B0(mai_mai_n411_), .Y(mai_mai_n428_));
  NA3        m0400(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n429_));
  NO2        m0401(.A(mai_mai_n429_), .B(mai_mai_n411_), .Y(mai_mai_n430_));
  NAi31      m0402(.An(b), .B(c), .C(a), .Y(mai_mai_n431_));
  NO2        m0403(.A(mai_mai_n431_), .B(n), .Y(mai_mai_n432_));
  OAI210     m0404(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n433_));
  NO2        m0405(.A(mai_mai_n433_), .B(mai_mai_n146_), .Y(mai_mai_n434_));
  NA2        m0406(.A(mai_mai_n434_), .B(mai_mai_n432_), .Y(mai_mai_n435_));
  INV        m0407(.A(mai_mai_n435_), .Y(mai_mai_n436_));
  NO4        m0408(.A(mai_mai_n436_), .B(mai_mai_n430_), .C(mai_mai_n428_), .D(mai_mai_n409_), .Y(mai_mai_n437_));
  NA2        m0409(.A(i), .B(g), .Y(mai_mai_n438_));
  NO3        m0410(.A(mai_mai_n277_), .B(mai_mai_n438_), .C(c), .Y(mai_mai_n439_));
  NOi21      m0411(.An(a), .B(n), .Y(mai_mai_n440_));
  NOi21      m0412(.An(d), .B(c), .Y(mai_mai_n441_));
  NA2        m0413(.A(mai_mai_n441_), .B(mai_mai_n440_), .Y(mai_mai_n442_));
  NA3        m0414(.A(i), .B(g), .C(f), .Y(mai_mai_n443_));
  OR2        m0415(.A(mai_mai_n443_), .B(mai_mai_n71_), .Y(mai_mai_n444_));
  NA2        m0416(.A(mai_mai_n439_), .B(mai_mai_n291_), .Y(mai_mai_n445_));
  OR2        m0417(.A(n), .B(m), .Y(mai_mai_n446_));
  NO2        m0418(.A(mai_mai_n446_), .B(mai_mai_n151_), .Y(mai_mai_n447_));
  NO2        m0419(.A(mai_mai_n183_), .B(mai_mai_n146_), .Y(mai_mai_n448_));
  OAI210     m0420(.A0(mai_mai_n447_), .A1(mai_mai_n176_), .B0(mai_mai_n448_), .Y(mai_mai_n449_));
  INV        m0421(.A(mai_mai_n375_), .Y(mai_mai_n450_));
  NA3        m0422(.A(mai_mai_n450_), .B(mai_mai_n363_), .C(d), .Y(mai_mai_n451_));
  NAi21      m0423(.An(k), .B(j), .Y(mai_mai_n452_));
  NAi21      m0424(.An(e), .B(d), .Y(mai_mai_n453_));
  NO2        m0425(.A(mai_mai_n453_), .B(mai_mai_n56_), .Y(mai_mai_n454_));
  NO2        m0426(.A(mai_mai_n253_), .B(mai_mai_n214_), .Y(mai_mai_n455_));
  NA3        m0427(.A(mai_mai_n455_), .B(mai_mai_n454_), .C(mai_mai_n226_), .Y(mai_mai_n456_));
  NA3        m0428(.A(mai_mai_n456_), .B(mai_mai_n451_), .C(mai_mai_n449_), .Y(mai_mai_n457_));
  NO2        m0429(.A(mai_mai_n339_), .B(mai_mai_n214_), .Y(mai_mai_n458_));
  NA2        m0430(.A(mai_mai_n458_), .B(mai_mai_n454_), .Y(mai_mai_n459_));
  NOi31      m0431(.An(n), .B(m), .C(k), .Y(mai_mai_n460_));
  AOI220     m0432(.A0(mai_mai_n460_), .A1(mai_mai_n391_), .B0(mai_mai_n220_), .B1(mai_mai_n50_), .Y(mai_mai_n461_));
  NAi31      m0433(.An(g), .B(f), .C(c), .Y(mai_mai_n462_));
  OR3        m0434(.A(mai_mai_n462_), .B(mai_mai_n461_), .C(e), .Y(mai_mai_n463_));
  NA2        m0435(.A(mai_mai_n463_), .B(mai_mai_n459_), .Y(mai_mai_n464_));
  NOi41      m0436(.An(mai_mai_n445_), .B(mai_mai_n464_), .C(mai_mai_n457_), .D(mai_mai_n267_), .Y(mai_mai_n465_));
  NOi32      m0437(.An(c), .Bn(a), .C(b), .Y(mai_mai_n466_));
  NA2        m0438(.A(mai_mai_n466_), .B(mai_mai_n114_), .Y(mai_mai_n467_));
  NA2        m0439(.A(mai_mai_n275_), .B(mai_mai_n151_), .Y(mai_mai_n468_));
  AN2        m0440(.A(e), .B(d), .Y(mai_mai_n469_));
  NA2        m0441(.A(mai_mai_n469_), .B(mai_mai_n468_), .Y(mai_mai_n470_));
  INV        m0442(.A(mai_mai_n146_), .Y(mai_mai_n471_));
  NO2        m0443(.A(mai_mai_n132_), .B(mai_mai_n41_), .Y(mai_mai_n472_));
  NO2        m0444(.A(mai_mai_n66_), .B(e), .Y(mai_mai_n473_));
  NOi31      m0445(.An(j), .B(k), .C(i), .Y(mai_mai_n474_));
  NOi21      m0446(.An(mai_mai_n164_), .B(mai_mai_n474_), .Y(mai_mai_n475_));
  NA4        m0447(.A(mai_mai_n324_), .B(mai_mai_n475_), .C(mai_mai_n261_), .D(mai_mai_n120_), .Y(mai_mai_n476_));
  AOI220     m0448(.A0(mai_mai_n476_), .A1(mai_mai_n473_), .B0(mai_mai_n472_), .B1(mai_mai_n471_), .Y(mai_mai_n477_));
  AOI210     m0449(.A0(mai_mai_n477_), .A1(mai_mai_n470_), .B0(mai_mai_n467_), .Y(mai_mai_n478_));
  NO2        m0450(.A(mai_mai_n210_), .B(mai_mai_n205_), .Y(mai_mai_n479_));
  NOi21      m0451(.An(a), .B(b), .Y(mai_mai_n480_));
  NA3        m0452(.A(e), .B(d), .C(c), .Y(mai_mai_n481_));
  NAi21      m0453(.An(mai_mai_n481_), .B(mai_mai_n480_), .Y(mai_mai_n482_));
  NO2        m0454(.A(mai_mai_n479_), .B(mai_mai_n482_), .Y(mai_mai_n483_));
  NO4        m0455(.A(mai_mai_n187_), .B(mai_mai_n103_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n484_));
  NA2        m0456(.A(mai_mai_n386_), .B(mai_mai_n152_), .Y(mai_mai_n485_));
  OR2        m0457(.A(k), .B(j), .Y(mai_mai_n486_));
  NA2        m0458(.A(l), .B(k), .Y(mai_mai_n487_));
  NA3        m0459(.A(mai_mai_n487_), .B(mai_mai_n486_), .C(mai_mai_n220_), .Y(mai_mai_n488_));
  AOI210     m0460(.A0(mai_mai_n233_), .A1(mai_mai_n342_), .B0(mai_mai_n86_), .Y(mai_mai_n489_));
  NOi21      m0461(.An(mai_mai_n488_), .B(mai_mai_n489_), .Y(mai_mai_n490_));
  OR3        m0462(.A(mai_mai_n490_), .B(mai_mai_n143_), .C(mai_mai_n135_), .Y(mai_mai_n491_));
  INV        m0463(.A(mai_mai_n129_), .Y(mai_mai_n492_));
  NA2        m0464(.A(mai_mai_n399_), .B(mai_mai_n114_), .Y(mai_mai_n493_));
  NO4        m0465(.A(mai_mai_n493_), .B(mai_mai_n95_), .C(mai_mai_n113_), .D(e), .Y(mai_mai_n494_));
  NO3        m0466(.A(mai_mai_n494_), .B(mai_mai_n492_), .C(mai_mai_n325_), .Y(mai_mai_n495_));
  NA3        m0467(.A(mai_mai_n495_), .B(mai_mai_n491_), .C(mai_mai_n485_), .Y(mai_mai_n496_));
  NO4        m0468(.A(mai_mai_n496_), .B(mai_mai_n484_), .C(mai_mai_n483_), .D(mai_mai_n478_), .Y(mai_mai_n497_));
  NA2        m0469(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n498_));
  NOi21      m0470(.An(d), .B(e), .Y(mai_mai_n499_));
  NAi31      m0471(.An(j), .B(l), .C(i), .Y(mai_mai_n500_));
  OAI210     m0472(.A0(mai_mai_n500_), .A1(mai_mai_n133_), .B0(mai_mai_n103_), .Y(mai_mai_n501_));
  NO3        m0473(.A(mai_mai_n400_), .B(mai_mai_n348_), .C(mai_mai_n201_), .Y(mai_mai_n502_));
  NO2        m0474(.A(mai_mai_n400_), .B(mai_mai_n375_), .Y(mai_mai_n503_));
  NO3        m0475(.A(mai_mai_n503_), .B(mai_mai_n502_), .C(mai_mai_n308_), .Y(mai_mai_n504_));
  NA3        m0476(.A(mai_mai_n504_), .B(mai_mai_n498_), .C(mai_mai_n243_), .Y(mai_mai_n505_));
  OAI210     m0477(.A0(mai_mai_n128_), .A1(mai_mai_n127_), .B0(n), .Y(mai_mai_n506_));
  NO2        m0478(.A(mai_mai_n506_), .B(mai_mai_n132_), .Y(mai_mai_n507_));
  OA210      m0479(.A0(mai_mai_n245_), .A1(mai_mai_n507_), .B0(mai_mai_n192_), .Y(mai_mai_n508_));
  XO2        m0480(.A(i), .B(h), .Y(mai_mai_n509_));
  NA3        m0481(.A(mai_mai_n509_), .B(mai_mai_n158_), .C(n), .Y(mai_mai_n510_));
  NAi41      m0482(.An(mai_mai_n300_), .B(mai_mai_n510_), .C(mai_mai_n461_), .D(mai_mai_n388_), .Y(mai_mai_n511_));
  NOi32      m0483(.An(mai_mai_n511_), .Bn(mai_mai_n473_), .C(mai_mai_n272_), .Y(mai_mai_n512_));
  NAi31      m0484(.An(c), .B(f), .C(d), .Y(mai_mai_n513_));
  AOI210     m0485(.A0(mai_mai_n280_), .A1(mai_mai_n195_), .B0(mai_mai_n513_), .Y(mai_mai_n514_));
  NOi21      m0486(.An(mai_mai_n84_), .B(mai_mai_n514_), .Y(mai_mai_n515_));
  NA3        m0487(.A(mai_mai_n384_), .B(mai_mai_n98_), .C(mai_mai_n97_), .Y(mai_mai_n516_));
  NA2        m0488(.A(mai_mai_n227_), .B(mai_mai_n109_), .Y(mai_mai_n517_));
  AOI210     m0489(.A0(mai_mai_n517_), .A1(mai_mai_n181_), .B0(mai_mai_n513_), .Y(mai_mai_n518_));
  AOI210     m0490(.A0(mai_mai_n361_), .A1(mai_mai_n35_), .B0(mai_mai_n482_), .Y(mai_mai_n519_));
  NOi31      m0491(.An(mai_mai_n516_), .B(mai_mai_n519_), .C(mai_mai_n518_), .Y(mai_mai_n520_));
  AO220      m0492(.A0(mai_mai_n288_), .A1(mai_mai_n264_), .B0(mai_mai_n165_), .B1(mai_mai_n67_), .Y(mai_mai_n521_));
  NA3        m0493(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n522_));
  NO2        m0494(.A(mai_mai_n522_), .B(mai_mai_n442_), .Y(mai_mai_n523_));
  NO2        m0495(.A(mai_mai_n523_), .B(mai_mai_n296_), .Y(mai_mai_n524_));
  NAi41      m0496(.An(mai_mai_n521_), .B(mai_mai_n524_), .C(mai_mai_n520_), .D(mai_mai_n515_), .Y(mai_mai_n525_));
  NO4        m0497(.A(mai_mai_n525_), .B(mai_mai_n512_), .C(mai_mai_n508_), .D(mai_mai_n505_), .Y(mai_mai_n526_));
  NA4        m0498(.A(mai_mai_n526_), .B(mai_mai_n497_), .C(mai_mai_n465_), .D(mai_mai_n437_), .Y(mai11));
  NO2        m0499(.A(mai_mai_n73_), .B(f), .Y(mai_mai_n528_));
  NA2        m0500(.A(j), .B(g), .Y(mai_mai_n529_));
  NAi31      m0501(.An(i), .B(m), .C(l), .Y(mai_mai_n530_));
  NA3        m0502(.A(m), .B(k), .C(j), .Y(mai_mai_n531_));
  OAI220     m0503(.A0(mai_mai_n531_), .A1(mai_mai_n132_), .B0(mai_mai_n530_), .B1(mai_mai_n529_), .Y(mai_mai_n532_));
  NOi32      m0504(.An(e), .Bn(b), .C(f), .Y(mai_mai_n533_));
  NA2        m0505(.A(mai_mai_n260_), .B(mai_mai_n114_), .Y(mai_mai_n534_));
  NA2        m0506(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n535_));
  OAI220     m0507(.A0(mai_mai_n535_), .A1(mai_mai_n302_), .B0(mai_mai_n534_), .B1(mai_mai_n215_), .Y(mai_mai_n536_));
  NAi31      m0508(.An(d), .B(e), .C(a), .Y(mai_mai_n537_));
  NO2        m0509(.A(mai_mai_n537_), .B(n), .Y(mai_mai_n538_));
  AOI220     m0510(.A0(mai_mai_n538_), .A1(mai_mai_n102_), .B0(mai_mai_n536_), .B1(mai_mai_n533_), .Y(mai_mai_n539_));
  NAi41      m0511(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n540_));
  AN2        m0512(.A(mai_mai_n540_), .B(mai_mai_n374_), .Y(mai_mai_n541_));
  AOI210     m0513(.A0(mai_mai_n541_), .A1(mai_mai_n400_), .B0(mai_mai_n273_), .Y(mai_mai_n542_));
  NA2        m0514(.A(j), .B(i), .Y(mai_mai_n543_));
  NAi31      m0515(.An(n), .B(m), .C(k), .Y(mai_mai_n544_));
  NO3        m0516(.A(mai_mai_n544_), .B(mai_mai_n543_), .C(mai_mai_n113_), .Y(mai_mai_n545_));
  NO4        m0517(.A(n), .B(d), .C(mai_mai_n117_), .D(a), .Y(mai_mai_n546_));
  OR2        m0518(.A(n), .B(c), .Y(mai_mai_n547_));
  NO2        m0519(.A(mai_mai_n547_), .B(mai_mai_n148_), .Y(mai_mai_n548_));
  NO2        m0520(.A(mai_mai_n548_), .B(mai_mai_n546_), .Y(mai_mai_n549_));
  NOi32      m0521(.An(g), .Bn(f), .C(i), .Y(mai_mai_n550_));
  AOI220     m0522(.A0(mai_mai_n550_), .A1(mai_mai_n100_), .B0(mai_mai_n532_), .B1(f), .Y(mai_mai_n551_));
  NO2        m0523(.A(mai_mai_n275_), .B(mai_mai_n49_), .Y(mai_mai_n552_));
  NO2        m0524(.A(mai_mai_n551_), .B(mai_mai_n549_), .Y(mai_mai_n553_));
  AOI210     m0525(.A0(mai_mai_n545_), .A1(mai_mai_n542_), .B0(mai_mai_n553_), .Y(mai_mai_n554_));
  NA2        m0526(.A(mai_mai_n140_), .B(mai_mai_n34_), .Y(mai_mai_n555_));
  OAI220     m0527(.A0(mai_mai_n555_), .A1(m), .B0(mai_mai_n535_), .B1(mai_mai_n233_), .Y(mai_mai_n556_));
  NOi41      m0528(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n557_));
  NAi32      m0529(.An(e), .Bn(b), .C(c), .Y(mai_mai_n558_));
  OR2        m0530(.A(mai_mai_n558_), .B(mai_mai_n86_), .Y(mai_mai_n559_));
  AN2        m0531(.A(mai_mai_n343_), .B(mai_mai_n321_), .Y(mai_mai_n560_));
  NA2        m0532(.A(mai_mai_n560_), .B(mai_mai_n559_), .Y(mai_mai_n561_));
  OA210      m0533(.A0(mai_mai_n561_), .A1(mai_mai_n557_), .B0(mai_mai_n556_), .Y(mai_mai_n562_));
  OAI220     m0534(.A0(mai_mai_n402_), .A1(mai_mai_n401_), .B0(mai_mai_n530_), .B1(mai_mai_n529_), .Y(mai_mai_n563_));
  NAi31      m0535(.An(d), .B(c), .C(a), .Y(mai_mai_n564_));
  NO2        m0536(.A(mai_mai_n564_), .B(n), .Y(mai_mai_n565_));
  NA3        m0537(.A(mai_mai_n565_), .B(mai_mai_n563_), .C(e), .Y(mai_mai_n566_));
  NO3        m0538(.A(mai_mai_n62_), .B(mai_mai_n49_), .C(mai_mai_n215_), .Y(mai_mai_n567_));
  NO2        m0539(.A(mai_mai_n230_), .B(mai_mai_n111_), .Y(mai_mai_n568_));
  OAI210     m0540(.A0(mai_mai_n567_), .A1(mai_mai_n403_), .B0(mai_mai_n568_), .Y(mai_mai_n569_));
  NA2        m0541(.A(mai_mai_n569_), .B(mai_mai_n566_), .Y(mai_mai_n570_));
  NO2        m0542(.A(mai_mai_n277_), .B(n), .Y(mai_mai_n571_));
  NO2        m0543(.A(mai_mai_n432_), .B(mai_mai_n571_), .Y(mai_mai_n572_));
  NA2        m0544(.A(mai_mai_n563_), .B(f), .Y(mai_mai_n573_));
  NAi32      m0545(.An(d), .Bn(a), .C(b), .Y(mai_mai_n574_));
  NA2        m0546(.A(h), .B(f), .Y(mai_mai_n575_));
  NO2        m0547(.A(mai_mai_n575_), .B(mai_mai_n95_), .Y(mai_mai_n576_));
  NO2        m0548(.A(mai_mai_n573_), .B(mai_mai_n572_), .Y(mai_mai_n577_));
  NO2        m0549(.A(mai_mai_n145_), .B(c), .Y(mai_mai_n578_));
  NA3        m0550(.A(f), .B(d), .C(b), .Y(mai_mai_n579_));
  NO3        m0551(.A(mai_mai_n577_), .B(mai_mai_n570_), .C(mai_mai_n562_), .Y(mai_mai_n580_));
  AN3        m0552(.A(mai_mai_n580_), .B(mai_mai_n554_), .C(mai_mai_n539_), .Y(mai_mai_n581_));
  INV        m0553(.A(k), .Y(mai_mai_n582_));
  NA3        m0554(.A(l), .B(mai_mai_n582_), .C(i), .Y(mai_mai_n583_));
  INV        m0555(.A(mai_mai_n583_), .Y(mai_mai_n584_));
  NA4        m0556(.A(mai_mai_n399_), .B(mai_mai_n422_), .C(mai_mai_n182_), .D(mai_mai_n114_), .Y(mai_mai_n585_));
  NAi32      m0557(.An(h), .Bn(f), .C(g), .Y(mai_mai_n586_));
  NAi41      m0558(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n587_));
  OAI210     m0559(.A0(mai_mai_n537_), .A1(n), .B0(mai_mai_n587_), .Y(mai_mai_n588_));
  NA2        m0560(.A(mai_mai_n588_), .B(m), .Y(mai_mai_n589_));
  NAi31      m0561(.An(h), .B(g), .C(f), .Y(mai_mai_n590_));
  OR3        m0562(.A(mai_mai_n590_), .B(mai_mai_n277_), .C(mai_mai_n49_), .Y(mai_mai_n591_));
  NA4        m0563(.A(mai_mai_n422_), .B(mai_mai_n122_), .C(mai_mai_n114_), .D(e), .Y(mai_mai_n592_));
  AN2        m0564(.A(mai_mai_n592_), .B(mai_mai_n591_), .Y(mai_mai_n593_));
  OA210      m0565(.A0(mai_mai_n589_), .A1(mai_mai_n586_), .B0(mai_mai_n593_), .Y(mai_mai_n594_));
  NO4        m0566(.A(mai_mai_n590_), .B(mai_mai_n547_), .C(mai_mai_n148_), .D(mai_mai_n75_), .Y(mai_mai_n595_));
  NAi31      m0567(.An(mai_mai_n595_), .B(mai_mai_n594_), .C(mai_mai_n585_), .Y(mai_mai_n596_));
  NAi31      m0568(.An(f), .B(h), .C(g), .Y(mai_mai_n597_));
  NO4        m0569(.A(mai_mai_n312_), .B(mai_mai_n597_), .C(mai_mai_n73_), .D(mai_mai_n75_), .Y(mai_mai_n598_));
  NOi32      m0570(.An(b), .Bn(a), .C(c), .Y(mai_mai_n599_));
  NOi41      m0571(.An(mai_mai_n599_), .B(mai_mai_n354_), .C(mai_mai_n69_), .D(mai_mai_n118_), .Y(mai_mai_n600_));
  OR2        m0572(.A(mai_mai_n600_), .B(mai_mai_n598_), .Y(mai_mai_n601_));
  NOi32      m0573(.An(d), .Bn(a), .C(e), .Y(mai_mai_n602_));
  NA2        m0574(.A(mai_mai_n602_), .B(mai_mai_n114_), .Y(mai_mai_n603_));
  NO2        m0575(.A(n), .B(c), .Y(mai_mai_n604_));
  NA3        m0576(.A(mai_mai_n604_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n605_));
  NAi32      m0577(.An(n), .Bn(f), .C(m), .Y(mai_mai_n606_));
  NA3        m0578(.A(mai_mai_n606_), .B(mai_mai_n605_), .C(mai_mai_n603_), .Y(mai_mai_n607_));
  NOi32      m0579(.An(e), .Bn(a), .C(d), .Y(mai_mai_n608_));
  AOI210     m0580(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n608_), .Y(mai_mai_n609_));
  AOI210     m0581(.A0(mai_mai_n609_), .A1(mai_mai_n214_), .B0(mai_mai_n555_), .Y(mai_mai_n610_));
  AOI210     m0582(.A0(mai_mai_n610_), .A1(mai_mai_n607_), .B0(mai_mai_n601_), .Y(mai_mai_n611_));
  INV        m0583(.A(mai_mai_n611_), .Y(mai_mai_n612_));
  AOI210     m0584(.A0(mai_mai_n596_), .A1(mai_mai_n584_), .B0(mai_mai_n612_), .Y(mai_mai_n613_));
  NO3        m0585(.A(mai_mai_n319_), .B(mai_mai_n61_), .C(n), .Y(mai_mai_n614_));
  NA3        m0586(.A(mai_mai_n513_), .B(mai_mai_n172_), .C(mai_mai_n171_), .Y(mai_mai_n615_));
  NA2        m0587(.A(mai_mai_n462_), .B(mai_mai_n230_), .Y(mai_mai_n616_));
  OR2        m0588(.A(mai_mai_n616_), .B(mai_mai_n615_), .Y(mai_mai_n617_));
  NA2        m0589(.A(mai_mai_n76_), .B(mai_mai_n114_), .Y(mai_mai_n618_));
  NO2        m0590(.A(mai_mai_n618_), .B(mai_mai_n45_), .Y(mai_mai_n619_));
  AOI220     m0591(.A0(mai_mai_n619_), .A1(mai_mai_n542_), .B0(mai_mai_n617_), .B1(mai_mai_n614_), .Y(mai_mai_n620_));
  NO2        m0592(.A(mai_mai_n620_), .B(mai_mai_n89_), .Y(mai_mai_n621_));
  NA3        m0593(.A(mai_mai_n557_), .B(mai_mai_n344_), .C(mai_mai_n46_), .Y(mai_mai_n622_));
  NOi32      m0594(.An(e), .Bn(c), .C(f), .Y(mai_mai_n623_));
  NOi21      m0595(.An(f), .B(g), .Y(mai_mai_n624_));
  NO2        m0596(.A(mai_mai_n624_), .B(mai_mai_n212_), .Y(mai_mai_n625_));
  AOI220     m0597(.A0(mai_mai_n625_), .A1(mai_mai_n396_), .B0(mai_mai_n623_), .B1(mai_mai_n176_), .Y(mai_mai_n626_));
  NA3        m0598(.A(mai_mai_n626_), .B(mai_mai_n622_), .C(mai_mai_n179_), .Y(mai_mai_n627_));
  AOI210     m0599(.A0(mai_mai_n541_), .A1(mai_mai_n400_), .B0(mai_mai_n301_), .Y(mai_mai_n628_));
  NA2        m0600(.A(mai_mai_n628_), .B(mai_mai_n265_), .Y(mai_mai_n629_));
  NOi21      m0601(.An(j), .B(l), .Y(mai_mai_n630_));
  NAi21      m0602(.An(k), .B(h), .Y(mai_mai_n631_));
  NO2        m0603(.A(mai_mai_n631_), .B(mai_mai_n263_), .Y(mai_mai_n632_));
  NOi31      m0604(.An(m), .B(n), .C(k), .Y(mai_mai_n633_));
  NA2        m0605(.A(mai_mai_n630_), .B(mai_mai_n633_), .Y(mai_mai_n634_));
  AOI210     m0606(.A0(mai_mai_n400_), .A1(mai_mai_n374_), .B0(mai_mai_n301_), .Y(mai_mai_n635_));
  NAi21      m0607(.An(mai_mai_n634_), .B(mai_mai_n635_), .Y(mai_mai_n636_));
  NO2        m0608(.A(mai_mai_n277_), .B(mai_mai_n49_), .Y(mai_mai_n637_));
  NO2        m0609(.A(mai_mai_n537_), .B(mai_mai_n49_), .Y(mai_mai_n638_));
  NA2        m0610(.A(mai_mai_n637_), .B(mai_mai_n576_), .Y(mai_mai_n639_));
  NA3        m0611(.A(mai_mai_n639_), .B(mai_mai_n636_), .C(mai_mai_n629_), .Y(mai_mai_n640_));
  NA2        m0612(.A(mai_mai_n109_), .B(mai_mai_n36_), .Y(mai_mai_n641_));
  NO2        m0613(.A(k), .B(mai_mai_n215_), .Y(mai_mai_n642_));
  NO2        m0614(.A(mai_mai_n533_), .B(mai_mai_n363_), .Y(mai_mai_n643_));
  NO2        m0615(.A(mai_mai_n643_), .B(n), .Y(mai_mai_n644_));
  NAi31      m0616(.An(mai_mai_n641_), .B(mai_mai_n644_), .C(mai_mai_n642_), .Y(mai_mai_n645_));
  NO2        m0617(.A(mai_mai_n535_), .B(mai_mai_n177_), .Y(mai_mai_n646_));
  NA3        m0618(.A(mai_mai_n558_), .B(mai_mai_n272_), .C(mai_mai_n144_), .Y(mai_mai_n647_));
  NA2        m0619(.A(mai_mai_n509_), .B(mai_mai_n158_), .Y(mai_mai_n648_));
  NO3        m0620(.A(mai_mai_n397_), .B(mai_mai_n648_), .C(mai_mai_n89_), .Y(mai_mai_n649_));
  AOI210     m0621(.A0(mai_mai_n647_), .A1(mai_mai_n646_), .B0(mai_mai_n649_), .Y(mai_mai_n650_));
  AN3        m0622(.A(f), .B(d), .C(b), .Y(mai_mai_n651_));
  OAI210     m0623(.A0(mai_mai_n651_), .A1(mai_mai_n131_), .B0(n), .Y(mai_mai_n652_));
  NA3        m0624(.A(mai_mai_n509_), .B(mai_mai_n158_), .C(mai_mai_n215_), .Y(mai_mai_n653_));
  AOI210     m0625(.A0(mai_mai_n652_), .A1(mai_mai_n232_), .B0(mai_mai_n653_), .Y(mai_mai_n654_));
  NAi31      m0626(.An(m), .B(n), .C(k), .Y(mai_mai_n655_));
  INV        m0627(.A(mai_mai_n251_), .Y(mai_mai_n656_));
  OAI210     m0628(.A0(mai_mai_n656_), .A1(mai_mai_n654_), .B0(j), .Y(mai_mai_n657_));
  NA3        m0629(.A(mai_mai_n657_), .B(mai_mai_n650_), .C(mai_mai_n645_), .Y(mai_mai_n658_));
  NO4        m0630(.A(mai_mai_n658_), .B(mai_mai_n640_), .C(mai_mai_n627_), .D(mai_mai_n621_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n384_), .B(mai_mai_n161_), .Y(mai_mai_n660_));
  NAi31      m0632(.An(g), .B(h), .C(f), .Y(mai_mai_n661_));
  OR3        m0633(.A(mai_mai_n661_), .B(mai_mai_n277_), .C(n), .Y(mai_mai_n662_));
  OA210      m0634(.A0(mai_mai_n537_), .A1(n), .B0(mai_mai_n587_), .Y(mai_mai_n663_));
  NA3        m0635(.A(mai_mai_n420_), .B(mai_mai_n122_), .C(mai_mai_n86_), .Y(mai_mai_n664_));
  OAI210     m0636(.A0(mai_mai_n663_), .A1(mai_mai_n92_), .B0(mai_mai_n664_), .Y(mai_mai_n665_));
  NOi21      m0637(.An(mai_mai_n662_), .B(mai_mai_n665_), .Y(mai_mai_n666_));
  AOI210     m0638(.A0(mai_mai_n666_), .A1(mai_mai_n660_), .B0(mai_mai_n531_), .Y(mai_mai_n667_));
  NO3        m0639(.A(g), .B(mai_mai_n214_), .C(mai_mai_n56_), .Y(mai_mai_n668_));
  NAi21      m0640(.An(h), .B(j), .Y(mai_mai_n669_));
  NO2        m0641(.A(mai_mai_n517_), .B(mai_mai_n89_), .Y(mai_mai_n670_));
  OAI210     m0642(.A0(mai_mai_n670_), .A1(mai_mai_n396_), .B0(mai_mai_n668_), .Y(mai_mai_n671_));
  OR2        m0643(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n672_));
  NA2        m0644(.A(mai_mai_n599_), .B(mai_mai_n346_), .Y(mai_mai_n673_));
  OR2        m0645(.A(mai_mai_n634_), .B(mai_mai_n673_), .Y(mai_mai_n674_));
  NA3        m0646(.A(mai_mai_n528_), .B(mai_mai_n100_), .C(mai_mai_n99_), .Y(mai_mai_n675_));
  AN2        m0647(.A(h), .B(f), .Y(mai_mai_n676_));
  NA2        m0648(.A(mai_mai_n676_), .B(mai_mai_n37_), .Y(mai_mai_n677_));
  NA2        m0649(.A(mai_mai_n100_), .B(mai_mai_n46_), .Y(mai_mai_n678_));
  NO2        m0650(.A(mai_mai_n678_), .B(mai_mai_n336_), .Y(mai_mai_n679_));
  AOI210     m0651(.A0(mai_mai_n574_), .A1(mai_mai_n431_), .B0(mai_mai_n49_), .Y(mai_mai_n680_));
  OAI220     m0652(.A0(mai_mai_n590_), .A1(mai_mai_n583_), .B0(mai_mai_n329_), .B1(mai_mai_n529_), .Y(mai_mai_n681_));
  AOI210     m0653(.A0(mai_mai_n681_), .A1(mai_mai_n680_), .B0(mai_mai_n679_), .Y(mai_mai_n682_));
  NA4        m0654(.A(mai_mai_n682_), .B(mai_mai_n675_), .C(mai_mai_n674_), .D(mai_mai_n671_), .Y(mai_mai_n683_));
  NO2        m0655(.A(mai_mai_n252_), .B(f), .Y(mai_mai_n684_));
  NO2        m0656(.A(mai_mai_n624_), .B(mai_mai_n61_), .Y(mai_mai_n685_));
  NO3        m0657(.A(mai_mai_n685_), .B(mai_mai_n684_), .C(mai_mai_n34_), .Y(mai_mai_n686_));
  NA2        m0658(.A(mai_mai_n332_), .B(mai_mai_n140_), .Y(mai_mai_n687_));
  NA2        m0659(.A(mai_mai_n133_), .B(mai_mai_n49_), .Y(mai_mai_n688_));
  NA2        m0660(.A(mai_mai_n363_), .B(mai_mai_n114_), .Y(mai_mai_n689_));
  OA220      m0661(.A0(mai_mai_n689_), .A1(mai_mai_n555_), .B0(mai_mai_n361_), .B1(mai_mai_n112_), .Y(mai_mai_n690_));
  OAI210     m0662(.A0(mai_mai_n687_), .A1(mai_mai_n686_), .B0(mai_mai_n690_), .Y(mai_mai_n691_));
  NO3        m0663(.A(mai_mai_n407_), .B(mai_mai_n192_), .C(mai_mai_n191_), .Y(mai_mai_n692_));
  NA2        m0664(.A(mai_mai_n692_), .B(mai_mai_n230_), .Y(mai_mai_n693_));
  NA3        m0665(.A(mai_mai_n693_), .B(mai_mai_n254_), .C(j), .Y(mai_mai_n694_));
  NA2        m0666(.A(mai_mai_n466_), .B(mai_mai_n86_), .Y(mai_mai_n695_));
  NA3        m0667(.A(mai_mai_n694_), .B(mai_mai_n516_), .C(mai_mai_n405_), .Y(mai_mai_n696_));
  NO4        m0668(.A(mai_mai_n696_), .B(mai_mai_n691_), .C(mai_mai_n683_), .D(mai_mai_n667_), .Y(mai_mai_n697_));
  NA4        m0669(.A(mai_mai_n697_), .B(mai_mai_n659_), .C(mai_mai_n613_), .D(mai_mai_n581_), .Y(mai08));
  NO2        m0670(.A(k), .B(h), .Y(mai_mai_n699_));
  AO210      m0671(.A0(mai_mai_n252_), .A1(mai_mai_n452_), .B0(mai_mai_n699_), .Y(mai_mai_n700_));
  NO2        m0672(.A(mai_mai_n700_), .B(mai_mai_n299_), .Y(mai_mai_n701_));
  NA2        m0673(.A(mai_mai_n623_), .B(mai_mai_n86_), .Y(mai_mai_n702_));
  NA2        m0674(.A(mai_mai_n702_), .B(mai_mai_n462_), .Y(mai_mai_n703_));
  NA2        m0675(.A(mai_mai_n703_), .B(mai_mai_n701_), .Y(mai_mai_n704_));
  NA2        m0676(.A(mai_mai_n86_), .B(mai_mai_n111_), .Y(mai_mai_n705_));
  NO2        m0677(.A(mai_mai_n705_), .B(mai_mai_n57_), .Y(mai_mai_n706_));
  NO4        m0678(.A(mai_mai_n381_), .B(mai_mai_n113_), .C(j), .D(mai_mai_n215_), .Y(mai_mai_n707_));
  NA2        m0679(.A(mai_mai_n579_), .B(mai_mai_n232_), .Y(mai_mai_n708_));
  AOI220     m0680(.A0(mai_mai_n708_), .A1(mai_mai_n350_), .B0(mai_mai_n707_), .B1(mai_mai_n706_), .Y(mai_mai_n709_));
  AOI210     m0681(.A0(mai_mai_n579_), .A1(mai_mai_n154_), .B0(mai_mai_n86_), .Y(mai_mai_n710_));
  NA4        m0682(.A(mai_mai_n217_), .B(mai_mai_n140_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n711_));
  AN2        m0683(.A(l), .B(k), .Y(mai_mai_n712_));
  NO2        m0684(.A(mai_mai_n711_), .B(g), .Y(mai_mai_n713_));
  NA2        m0685(.A(mai_mai_n713_), .B(mai_mai_n710_), .Y(mai_mai_n714_));
  NA3        m0686(.A(mai_mai_n714_), .B(mai_mai_n709_), .C(mai_mai_n704_), .Y(mai_mai_n715_));
  INV        m0687(.A(mai_mai_n523_), .Y(mai_mai_n716_));
  NO2        m0688(.A(mai_mai_n38_), .B(mai_mai_n214_), .Y(mai_mai_n717_));
  NA2        m0689(.A(mai_mai_n717_), .B(mai_mai_n571_), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n718_), .B(mai_mai_n716_), .Y(mai_mai_n719_));
  NO2        m0691(.A(mai_mai_n541_), .B(mai_mai_n35_), .Y(mai_mai_n720_));
  INV        m0692(.A(mai_mai_n720_), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n700_), .B(mai_mai_n136_), .Y(mai_mai_n722_));
  NA2        m0694(.A(mai_mai_n722_), .B(mai_mai_n406_), .Y(mai_mai_n723_));
  OAI210     m0695(.A0(mai_mai_n721_), .A1(mai_mai_n89_), .B0(mai_mai_n723_), .Y(mai_mai_n724_));
  NA2        m0696(.A(mai_mai_n363_), .B(mai_mai_n43_), .Y(mai_mai_n725_));
  NA3        m0697(.A(mai_mai_n693_), .B(mai_mai_n338_), .C(mai_mai_n387_), .Y(mai_mai_n726_));
  NA2        m0698(.A(mai_mai_n712_), .B(mai_mai_n220_), .Y(mai_mai_n727_));
  NO2        m0699(.A(mai_mai_n727_), .B(mai_mai_n331_), .Y(mai_mai_n728_));
  AOI210     m0700(.A0(mai_mai_n728_), .A1(mai_mai_n684_), .B0(mai_mai_n494_), .Y(mai_mai_n729_));
  NA3        m0701(.A(m), .B(l), .C(k), .Y(mai_mai_n730_));
  AOI210     m0702(.A0(mai_mai_n664_), .A1(mai_mai_n662_), .B0(mai_mai_n730_), .Y(mai_mai_n731_));
  NO2        m0703(.A(mai_mai_n540_), .B(mai_mai_n273_), .Y(mai_mai_n732_));
  NOi21      m0704(.An(mai_mai_n732_), .B(mai_mai_n534_), .Y(mai_mai_n733_));
  NA4        m0705(.A(mai_mai_n114_), .B(l), .C(k), .D(mai_mai_n89_), .Y(mai_mai_n734_));
  NA3        m0706(.A(mai_mai_n122_), .B(mai_mai_n415_), .C(i), .Y(mai_mai_n735_));
  NO2        m0707(.A(mai_mai_n735_), .B(mai_mai_n734_), .Y(mai_mai_n736_));
  NO3        m0708(.A(mai_mai_n736_), .B(mai_mai_n733_), .C(mai_mai_n731_), .Y(mai_mai_n737_));
  NA4        m0709(.A(mai_mai_n737_), .B(mai_mai_n729_), .C(mai_mai_n726_), .D(mai_mai_n725_), .Y(mai_mai_n738_));
  NO4        m0710(.A(mai_mai_n738_), .B(mai_mai_n724_), .C(mai_mai_n719_), .D(mai_mai_n715_), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n625_), .B(mai_mai_n396_), .Y(mai_mai_n740_));
  NOi31      m0712(.An(g), .B(h), .C(f), .Y(mai_mai_n741_));
  NA2        m0713(.A(mai_mai_n638_), .B(mai_mai_n741_), .Y(mai_mai_n742_));
  AO210      m0714(.A0(mai_mai_n742_), .A1(mai_mai_n591_), .B0(mai_mai_n543_), .Y(mai_mai_n743_));
  INV        m0715(.A(mai_mai_n503_), .Y(mai_mai_n744_));
  NA4        m0716(.A(mai_mai_n744_), .B(mai_mai_n743_), .C(mai_mai_n740_), .D(mai_mai_n251_), .Y(mai_mai_n745_));
  NA2        m0717(.A(mai_mai_n712_), .B(mai_mai_n75_), .Y(mai_mai_n746_));
  NO4        m0718(.A(mai_mai_n692_), .B(mai_mai_n174_), .C(n), .D(i), .Y(mai_mai_n747_));
  NOi21      m0719(.An(h), .B(j), .Y(mai_mai_n748_));
  NA2        m0720(.A(mai_mai_n748_), .B(f), .Y(mai_mai_n749_));
  NO2        m0721(.A(mai_mai_n749_), .B(mai_mai_n247_), .Y(mai_mai_n750_));
  NO2        m0722(.A(mai_mai_n750_), .B(mai_mai_n747_), .Y(mai_mai_n751_));
  OAI220     m0723(.A0(mai_mai_n751_), .A1(mai_mai_n746_), .B0(mai_mai_n593_), .B1(mai_mai_n62_), .Y(mai_mai_n752_));
  AOI210     m0724(.A0(mai_mai_n745_), .A1(l), .B0(mai_mai_n752_), .Y(mai_mai_n753_));
  NO2        m0725(.A(j), .B(i), .Y(mai_mai_n754_));
  NA3        m0726(.A(mai_mai_n754_), .B(mai_mai_n82_), .C(l), .Y(mai_mai_n755_));
  NA2        m0727(.A(mai_mai_n754_), .B(mai_mai_n33_), .Y(mai_mai_n756_));
  NA2        m0728(.A(mai_mai_n425_), .B(mai_mai_n122_), .Y(mai_mai_n757_));
  OA220      m0729(.A0(mai_mai_n757_), .A1(mai_mai_n756_), .B0(mai_mai_n755_), .B1(mai_mai_n589_), .Y(mai_mai_n758_));
  NO3        m0730(.A(mai_mai_n150_), .B(mai_mai_n49_), .C(mai_mai_n111_), .Y(mai_mai_n759_));
  NO3        m0731(.A(mai_mai_n547_), .B(mai_mai_n148_), .C(mai_mai_n75_), .Y(mai_mai_n760_));
  NO3        m0732(.A(mai_mai_n487_), .B(mai_mai_n443_), .C(j), .Y(mai_mai_n761_));
  OAI210     m0733(.A0(mai_mai_n760_), .A1(mai_mai_n759_), .B0(mai_mai_n761_), .Y(mai_mai_n762_));
  OAI210     m0734(.A0(mai_mai_n742_), .A1(mai_mai_n62_), .B0(mai_mai_n762_), .Y(mai_mai_n763_));
  NA2        m0735(.A(k), .B(j), .Y(mai_mai_n764_));
  NO3        m0736(.A(mai_mai_n299_), .B(mai_mai_n764_), .C(mai_mai_n40_), .Y(mai_mai_n765_));
  AOI210     m0737(.A0(mai_mai_n533_), .A1(n), .B0(mai_mai_n557_), .Y(mai_mai_n766_));
  NA2        m0738(.A(mai_mai_n766_), .B(mai_mai_n560_), .Y(mai_mai_n767_));
  AN3        m0739(.A(mai_mai_n767_), .B(mai_mai_n765_), .C(mai_mai_n99_), .Y(mai_mai_n768_));
  NO3        m0740(.A(mai_mai_n174_), .B(mai_mai_n395_), .C(mai_mai_n113_), .Y(mai_mai_n769_));
  AOI220     m0741(.A0(mai_mai_n769_), .A1(mai_mai_n248_), .B0(mai_mai_n616_), .B1(mai_mai_n310_), .Y(mai_mai_n770_));
  INV        m0742(.A(mai_mai_n770_), .Y(mai_mai_n771_));
  NO2        m0743(.A(mai_mai_n299_), .B(mai_mai_n136_), .Y(mai_mai_n772_));
  NA2        m0744(.A(mai_mai_n772_), .B(mai_mai_n625_), .Y(mai_mai_n773_));
  NO2        m0745(.A(mai_mai_n730_), .B(mai_mai_n92_), .Y(mai_mai_n774_));
  NA2        m0746(.A(mai_mai_n774_), .B(mai_mai_n588_), .Y(mai_mai_n775_));
  NO2        m0747(.A(mai_mai_n590_), .B(mai_mai_n118_), .Y(mai_mai_n776_));
  OAI210     m0748(.A0(mai_mai_n776_), .A1(mai_mai_n761_), .B0(mai_mai_n680_), .Y(mai_mai_n777_));
  NA3        m0749(.A(mai_mai_n777_), .B(mai_mai_n775_), .C(mai_mai_n773_), .Y(mai_mai_n778_));
  OR4        m0750(.A(mai_mai_n778_), .B(mai_mai_n771_), .C(mai_mai_n768_), .D(mai_mai_n763_), .Y(mai_mai_n779_));
  NA3        m0751(.A(mai_mai_n766_), .B(mai_mai_n560_), .C(mai_mai_n559_), .Y(mai_mai_n780_));
  NA4        m0752(.A(mai_mai_n780_), .B(mai_mai_n217_), .C(mai_mai_n452_), .D(mai_mai_n34_), .Y(mai_mai_n781_));
  OAI220     m0753(.A0(mai_mai_n711_), .A1(mai_mai_n702_), .B0(mai_mai_n336_), .B1(mai_mai_n38_), .Y(mai_mai_n782_));
  INV        m0754(.A(mai_mai_n782_), .Y(mai_mai_n783_));
  NA3        m0755(.A(mai_mai_n550_), .B(mai_mai_n292_), .C(h), .Y(mai_mai_n784_));
  NOi21      m0756(.An(mai_mai_n680_), .B(mai_mai_n784_), .Y(mai_mai_n785_));
  NO2        m0757(.A(mai_mai_n93_), .B(mai_mai_n47_), .Y(mai_mai_n786_));
  OAI220     m0758(.A0(mai_mai_n784_), .A1(mai_mai_n605_), .B0(mai_mai_n755_), .B1(mai_mai_n672_), .Y(mai_mai_n787_));
  AOI210     m0759(.A0(mai_mai_n786_), .A1(mai_mai_n644_), .B0(mai_mai_n787_), .Y(mai_mai_n788_));
  NAi41      m0760(.An(mai_mai_n785_), .B(mai_mai_n788_), .C(mai_mai_n783_), .D(mai_mai_n781_), .Y(mai_mai_n789_));
  BUFFER     m0761(.A(mai_mai_n96_), .Y(mai_mai_n790_));
  AOI220     m0762(.A0(mai_mai_n790_), .A1(mai_mai_n238_), .B0(mai_mai_n761_), .B1(mai_mai_n637_), .Y(mai_mai_n791_));
  INV        m0763(.A(mai_mai_n340_), .Y(mai_mai_n792_));
  OAI210     m0764(.A0(mai_mai_n730_), .A1(mai_mai_n661_), .B0(mai_mai_n522_), .Y(mai_mai_n793_));
  NA3        m0765(.A(mai_mai_n250_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n794_));
  AOI220     m0766(.A0(mai_mai_n604_), .A1(mai_mai_n29_), .B0(mai_mai_n466_), .B1(mai_mai_n86_), .Y(mai_mai_n795_));
  NA2        m0767(.A(mai_mai_n795_), .B(mai_mai_n794_), .Y(mai_mai_n796_));
  NO2        m0768(.A(mai_mai_n784_), .B(mai_mai_n493_), .Y(mai_mai_n797_));
  AOI210     m0769(.A0(mai_mai_n796_), .A1(mai_mai_n793_), .B0(mai_mai_n797_), .Y(mai_mai_n798_));
  NA3        m0770(.A(mai_mai_n798_), .B(mai_mai_n792_), .C(mai_mai_n791_), .Y(mai_mai_n799_));
  NOi41      m0771(.An(mai_mai_n758_), .B(mai_mai_n799_), .C(mai_mai_n789_), .D(mai_mai_n779_), .Y(mai_mai_n800_));
  OR3        m0772(.A(mai_mai_n711_), .B(mai_mai_n232_), .C(g), .Y(mai_mai_n801_));
  NO3        m0773(.A(mai_mai_n345_), .B(mai_mai_n301_), .C(mai_mai_n113_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n802_), .B(mai_mai_n767_), .Y(mai_mai_n803_));
  NA2        m0775(.A(mai_mai_n46_), .B(mai_mai_n56_), .Y(mai_mai_n804_));
  NO3        m0776(.A(mai_mai_n804_), .B(mai_mai_n756_), .C(mai_mai_n277_), .Y(mai_mai_n805_));
  NO3        m0777(.A(mai_mai_n529_), .B(mai_mai_n94_), .C(h), .Y(mai_mai_n806_));
  AOI210     m0778(.A0(mai_mai_n806_), .A1(mai_mai_n706_), .B0(mai_mai_n805_), .Y(mai_mai_n807_));
  NA4        m0779(.A(mai_mai_n807_), .B(mai_mai_n803_), .C(mai_mai_n801_), .D(mai_mai_n408_), .Y(mai_mai_n808_));
  OR2        m0780(.A(mai_mai_n661_), .B(mai_mai_n93_), .Y(mai_mai_n809_));
  NOi31      m0781(.An(b), .B(d), .C(a), .Y(mai_mai_n810_));
  NO2        m0782(.A(mai_mai_n810_), .B(mai_mai_n602_), .Y(mai_mai_n811_));
  NO2        m0783(.A(mai_mai_n811_), .B(n), .Y(mai_mai_n812_));
  NOi21      m0784(.An(mai_mai_n795_), .B(mai_mai_n812_), .Y(mai_mai_n813_));
  OAI220     m0785(.A0(mai_mai_n813_), .A1(mai_mai_n809_), .B0(mai_mai_n784_), .B1(mai_mai_n603_), .Y(mai_mai_n814_));
  NO2        m0786(.A(mai_mai_n558_), .B(mai_mai_n86_), .Y(mai_mai_n815_));
  NO3        m0787(.A(mai_mai_n624_), .B(mai_mai_n331_), .C(mai_mai_n118_), .Y(mai_mai_n816_));
  NOi21      m0788(.An(mai_mai_n816_), .B(mai_mai_n159_), .Y(mai_mai_n817_));
  AOI210     m0789(.A0(mai_mai_n802_), .A1(mai_mai_n815_), .B0(mai_mai_n817_), .Y(mai_mai_n818_));
  OAI210     m0790(.A0(mai_mai_n711_), .A1(mai_mai_n397_), .B0(mai_mai_n818_), .Y(mai_mai_n819_));
  NO2        m0791(.A(mai_mai_n692_), .B(n), .Y(mai_mai_n820_));
  AOI220     m0792(.A0(mai_mai_n772_), .A1(mai_mai_n668_), .B0(mai_mai_n820_), .B1(mai_mai_n701_), .Y(mai_mai_n821_));
  NO2        m0793(.A(mai_mai_n326_), .B(mai_mai_n237_), .Y(mai_mai_n822_));
  NA2        m0794(.A(mai_mai_n122_), .B(mai_mai_n86_), .Y(mai_mai_n823_));
  AOI210     m0795(.A0(mai_mai_n429_), .A1(mai_mai_n421_), .B0(mai_mai_n823_), .Y(mai_mai_n824_));
  NA2        m0796(.A(mai_mai_n728_), .B(mai_mai_n34_), .Y(mai_mai_n825_));
  NAi21      m0797(.An(mai_mai_n734_), .B(mai_mai_n439_), .Y(mai_mai_n826_));
  NO2        m0798(.A(mai_mai_n273_), .B(i), .Y(mai_mai_n827_));
  NA2        m0799(.A(mai_mai_n595_), .B(mai_mai_n364_), .Y(mai_mai_n828_));
  AN2        m0800(.A(mai_mai_n828_), .B(mai_mai_n826_), .Y(mai_mai_n829_));
  NAi41      m0801(.An(mai_mai_n824_), .B(mai_mai_n829_), .C(mai_mai_n825_), .D(mai_mai_n821_), .Y(mai_mai_n830_));
  NO4        m0802(.A(mai_mai_n830_), .B(mai_mai_n819_), .C(mai_mai_n814_), .D(mai_mai_n808_), .Y(mai_mai_n831_));
  NA4        m0803(.A(mai_mai_n831_), .B(mai_mai_n800_), .C(mai_mai_n753_), .D(mai_mai_n739_), .Y(mai09));
  INV        m0804(.A(mai_mai_n123_), .Y(mai_mai_n833_));
  NA2        m0805(.A(f), .B(e), .Y(mai_mai_n834_));
  NO2        m0806(.A(mai_mai_n225_), .B(mai_mai_n113_), .Y(mai_mai_n835_));
  NA2        m0807(.A(mai_mai_n835_), .B(g), .Y(mai_mai_n836_));
  NA4        m0808(.A(mai_mai_n312_), .B(mai_mai_n475_), .C(mai_mai_n261_), .D(mai_mai_n120_), .Y(mai_mai_n837_));
  AOI210     m0809(.A0(mai_mai_n837_), .A1(g), .B0(mai_mai_n472_), .Y(mai_mai_n838_));
  AOI210     m0810(.A0(mai_mai_n838_), .A1(mai_mai_n836_), .B0(mai_mai_n834_), .Y(mai_mai_n839_));
  NA2        m0811(.A(mai_mai_n447_), .B(e), .Y(mai_mai_n840_));
  NO2        m0812(.A(mai_mai_n840_), .B(mai_mai_n513_), .Y(mai_mai_n841_));
  AOI210     m0813(.A0(mai_mai_n839_), .A1(mai_mai_n833_), .B0(mai_mai_n841_), .Y(mai_mai_n842_));
  NO2        m0814(.A(mai_mai_n204_), .B(mai_mai_n214_), .Y(mai_mai_n843_));
  NA3        m0815(.A(m), .B(l), .C(i), .Y(mai_mai_n844_));
  OAI220     m0816(.A0(mai_mai_n590_), .A1(mai_mai_n844_), .B0(mai_mai_n354_), .B1(mai_mai_n530_), .Y(mai_mai_n845_));
  NA4        m0817(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(g), .D(f), .Y(mai_mai_n846_));
  NAi31      m0818(.An(mai_mai_n845_), .B(mai_mai_n846_), .C(mai_mai_n444_), .Y(mai_mai_n847_));
  OA210      m0819(.A0(mai_mai_n847_), .A1(mai_mai_n843_), .B0(mai_mai_n571_), .Y(mai_mai_n848_));
  NA3        m0820(.A(mai_mai_n809_), .B(mai_mai_n573_), .C(mai_mai_n522_), .Y(mai_mai_n849_));
  OA210      m0821(.A0(mai_mai_n849_), .A1(mai_mai_n848_), .B0(mai_mai_n812_), .Y(mai_mai_n850_));
  INV        m0822(.A(mai_mai_n343_), .Y(mai_mai_n851_));
  NO2        m0823(.A(mai_mai_n128_), .B(mai_mai_n127_), .Y(mai_mai_n852_));
  INV        m0824(.A(mai_mai_n344_), .Y(mai_mai_n853_));
  AOI210     m0825(.A0(mai_mai_n853_), .A1(mai_mai_n852_), .B0(mai_mai_n597_), .Y(mai_mai_n854_));
  NA2        m0826(.A(mai_mai_n794_), .B(mai_mai_n336_), .Y(mai_mai_n855_));
  NA2        m0827(.A(mai_mai_n346_), .B(mai_mai_n347_), .Y(mai_mai_n856_));
  OAI210     m0828(.A0(mai_mai_n204_), .A1(mai_mai_n214_), .B0(mai_mai_n856_), .Y(mai_mai_n857_));
  AOI220     m0829(.A0(mai_mai_n857_), .A1(mai_mai_n855_), .B0(mai_mai_n854_), .B1(mai_mai_n851_), .Y(mai_mai_n858_));
  NA2        m0830(.A(mai_mai_n168_), .B(mai_mai_n115_), .Y(mai_mai_n859_));
  NA3        m0831(.A(mai_mai_n859_), .B(mai_mai_n700_), .C(mai_mai_n136_), .Y(mai_mai_n860_));
  NA3        m0832(.A(mai_mai_n860_), .B(mai_mai_n189_), .C(mai_mai_n31_), .Y(mai_mai_n861_));
  NA4        m0833(.A(mai_mai_n861_), .B(mai_mai_n858_), .C(mai_mai_n626_), .D(mai_mai_n84_), .Y(mai_mai_n862_));
  NO2        m0834(.A(mai_mai_n586_), .B(mai_mai_n500_), .Y(mai_mai_n863_));
  NOi21      m0835(.An(f), .B(d), .Y(mai_mai_n864_));
  NA2        m0836(.A(mai_mai_n864_), .B(m), .Y(mai_mai_n865_));
  NO2        m0837(.A(mai_mai_n865_), .B(mai_mai_n52_), .Y(mai_mai_n866_));
  NOi32      m0838(.An(g), .Bn(f), .C(d), .Y(mai_mai_n867_));
  NA4        m0839(.A(mai_mai_n867_), .B(mai_mai_n604_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n868_));
  NOi21      m0840(.An(mai_mai_n313_), .B(mai_mai_n868_), .Y(mai_mai_n869_));
  AOI210     m0841(.A0(mai_mai_n866_), .A1(mai_mai_n548_), .B0(mai_mai_n869_), .Y(mai_mai_n870_));
  NA3        m0842(.A(mai_mai_n312_), .B(mai_mai_n261_), .C(mai_mai_n120_), .Y(mai_mai_n871_));
  AN2        m0843(.A(f), .B(d), .Y(mai_mai_n872_));
  NA3        m0844(.A(mai_mai_n480_), .B(mai_mai_n872_), .C(mai_mai_n86_), .Y(mai_mai_n873_));
  NO3        m0845(.A(mai_mai_n873_), .B(mai_mai_n75_), .C(mai_mai_n215_), .Y(mai_mai_n874_));
  NO2        m0846(.A(mai_mai_n285_), .B(mai_mai_n56_), .Y(mai_mai_n875_));
  OAI210     m0847(.A0(mai_mai_n875_), .A1(mai_mai_n871_), .B0(mai_mai_n874_), .Y(mai_mai_n876_));
  NAi31      m0848(.An(mai_mai_n492_), .B(mai_mai_n876_), .C(mai_mai_n870_), .Y(mai_mai_n877_));
  NO4        m0849(.A(mai_mai_n624_), .B(mai_mai_n133_), .C(mai_mai_n331_), .D(mai_mai_n151_), .Y(mai_mai_n878_));
  NO2        m0850(.A(mai_mai_n655_), .B(mai_mai_n331_), .Y(mai_mai_n879_));
  AN2        m0851(.A(mai_mai_n879_), .B(mai_mai_n684_), .Y(mai_mai_n880_));
  NO3        m0852(.A(mai_mai_n880_), .B(mai_mai_n878_), .C(mai_mai_n234_), .Y(mai_mai_n881_));
  NA2        m0853(.A(mai_mai_n602_), .B(mai_mai_n86_), .Y(mai_mai_n882_));
  OAI220     m0854(.A0(mai_mai_n856_), .A1(mai_mai_n882_), .B0(mai_mai_n794_), .B1(mai_mai_n444_), .Y(mai_mai_n883_));
  NA3        m0855(.A(mai_mai_n158_), .B(mai_mai_n109_), .C(mai_mai_n108_), .Y(mai_mai_n884_));
  OAI220     m0856(.A0(mai_mai_n873_), .A1(mai_mai_n433_), .B0(mai_mai_n343_), .B1(mai_mai_n884_), .Y(mai_mai_n885_));
  NOi41      m0857(.An(mai_mai_n223_), .B(mai_mai_n885_), .C(mai_mai_n883_), .D(mai_mai_n308_), .Y(mai_mai_n886_));
  NA2        m0858(.A(c), .B(mai_mai_n117_), .Y(mai_mai_n887_));
  NO2        m0859(.A(mai_mai_n887_), .B(mai_mai_n412_), .Y(mai_mai_n888_));
  NA3        m0860(.A(mai_mai_n888_), .B(mai_mai_n511_), .C(f), .Y(mai_mai_n889_));
  OR2        m0861(.A(mai_mai_n661_), .B(mai_mai_n544_), .Y(mai_mai_n890_));
  INV        m0862(.A(mai_mai_n890_), .Y(mai_mai_n891_));
  NA2        m0863(.A(mai_mai_n811_), .B(mai_mai_n112_), .Y(mai_mai_n892_));
  NA2        m0864(.A(mai_mai_n892_), .B(mai_mai_n891_), .Y(mai_mai_n893_));
  NA4        m0865(.A(mai_mai_n893_), .B(mai_mai_n889_), .C(mai_mai_n886_), .D(mai_mai_n881_), .Y(mai_mai_n894_));
  NO4        m0866(.A(mai_mai_n894_), .B(mai_mai_n877_), .C(mai_mai_n862_), .D(mai_mai_n850_), .Y(mai_mai_n895_));
  NA2        m0867(.A(mai_mai_n113_), .B(j), .Y(mai_mai_n896_));
  AOI210     m0868(.A0(mai_mai_n794_), .A1(mai_mai_n336_), .B0(mai_mai_n846_), .Y(mai_mai_n897_));
  NO2        m0869(.A(mai_mai_n230_), .B(mai_mai_n224_), .Y(mai_mai_n898_));
  NA2        m0870(.A(mai_mai_n898_), .B(mai_mai_n227_), .Y(mai_mai_n899_));
  NO2        m0871(.A(mai_mai_n433_), .B(mai_mai_n834_), .Y(mai_mai_n900_));
  NA2        m0872(.A(mai_mai_n900_), .B(mai_mai_n565_), .Y(mai_mai_n901_));
  NA2        m0873(.A(mai_mai_n901_), .B(mai_mai_n899_), .Y(mai_mai_n902_));
  NA2        m0874(.A(e), .B(d), .Y(mai_mai_n903_));
  OAI220     m0875(.A0(mai_mai_n903_), .A1(c), .B0(mai_mai_n326_), .B1(d), .Y(mai_mai_n904_));
  NA3        m0876(.A(mai_mai_n904_), .B(mai_mai_n455_), .C(mai_mai_n509_), .Y(mai_mai_n905_));
  AOI210     m0877(.A0(mai_mai_n517_), .A1(mai_mai_n181_), .B0(mai_mai_n230_), .Y(mai_mai_n906_));
  INV        m0878(.A(mai_mai_n906_), .Y(mai_mai_n907_));
  NA2        m0879(.A(mai_mai_n285_), .B(mai_mai_n164_), .Y(mai_mai_n908_));
  NA2        m0880(.A(mai_mai_n874_), .B(mai_mai_n908_), .Y(mai_mai_n909_));
  NA3        m0881(.A(mai_mai_n167_), .B(mai_mai_n87_), .C(mai_mai_n34_), .Y(mai_mai_n910_));
  NA4        m0882(.A(mai_mai_n910_), .B(mai_mai_n909_), .C(mai_mai_n907_), .D(mai_mai_n905_), .Y(mai_mai_n911_));
  NO3        m0883(.A(mai_mai_n911_), .B(mai_mai_n902_), .C(mai_mai_n897_), .Y(mai_mai_n912_));
  NA2        m0884(.A(mai_mai_n851_), .B(mai_mai_n31_), .Y(mai_mai_n913_));
  AO210      m0885(.A0(mai_mai_n913_), .A1(mai_mai_n702_), .B0(mai_mai_n218_), .Y(mai_mai_n914_));
  OAI220     m0886(.A0(mai_mai_n624_), .A1(mai_mai_n61_), .B0(mai_mai_n301_), .B1(j), .Y(mai_mai_n915_));
  AOI220     m0887(.A0(mai_mai_n915_), .A1(mai_mai_n879_), .B0(mai_mai_n614_), .B1(mai_mai_n623_), .Y(mai_mai_n916_));
  OAI210     m0888(.A0(mai_mai_n840_), .A1(mai_mai_n171_), .B0(mai_mai_n916_), .Y(mai_mai_n917_));
  OAI210     m0889(.A0(mai_mai_n835_), .A1(mai_mai_n908_), .B0(mai_mai_n867_), .Y(mai_mai_n918_));
  NO2        m0890(.A(mai_mai_n918_), .B(mai_mai_n605_), .Y(mai_mai_n919_));
  AOI210     m0891(.A0(mai_mai_n119_), .A1(mai_mai_n118_), .B0(mai_mai_n260_), .Y(mai_mai_n920_));
  NO2        m0892(.A(mai_mai_n920_), .B(mai_mai_n868_), .Y(mai_mai_n921_));
  AO210      m0893(.A0(mai_mai_n855_), .A1(mai_mai_n845_), .B0(mai_mai_n921_), .Y(mai_mai_n922_));
  NOi31      m0894(.An(mai_mai_n548_), .B(mai_mai_n865_), .C(mai_mai_n293_), .Y(mai_mai_n923_));
  NO4        m0895(.A(mai_mai_n923_), .B(mai_mai_n922_), .C(mai_mai_n919_), .D(mai_mai_n917_), .Y(mai_mai_n924_));
  AO220      m0896(.A0(mai_mai_n455_), .A1(mai_mai_n748_), .B0(mai_mai_n176_), .B1(f), .Y(mai_mai_n925_));
  OAI210     m0897(.A0(mai_mai_n925_), .A1(mai_mai_n458_), .B0(mai_mai_n904_), .Y(mai_mai_n926_));
  NO2        m0898(.A(mai_mai_n443_), .B(mai_mai_n71_), .Y(mai_mai_n927_));
  OAI210     m0899(.A0(mai_mai_n849_), .A1(mai_mai_n927_), .B0(mai_mai_n706_), .Y(mai_mai_n928_));
  AN4        m0900(.A(mai_mai_n928_), .B(mai_mai_n926_), .C(mai_mai_n924_), .D(mai_mai_n914_), .Y(mai_mai_n929_));
  NA4        m0901(.A(mai_mai_n929_), .B(mai_mai_n912_), .C(mai_mai_n895_), .D(mai_mai_n842_), .Y(mai12));
  NO2        m0902(.A(mai_mai_n453_), .B(c), .Y(mai_mai_n931_));
  NO4        m0903(.A(mai_mai_n446_), .B(mai_mai_n252_), .C(mai_mai_n582_), .D(mai_mai_n215_), .Y(mai_mai_n932_));
  NA2        m0904(.A(mai_mai_n932_), .B(mai_mai_n931_), .Y(mai_mai_n933_));
  NA2        m0905(.A(mai_mai_n548_), .B(mai_mai_n927_), .Y(mai_mai_n934_));
  NO2        m0906(.A(mai_mai_n453_), .B(mai_mai_n117_), .Y(mai_mai_n935_));
  NO2        m0907(.A(mai_mai_n852_), .B(mai_mai_n354_), .Y(mai_mai_n936_));
  NO2        m0908(.A(mai_mai_n661_), .B(mai_mai_n381_), .Y(mai_mai_n937_));
  AOI220     m0909(.A0(mai_mai_n937_), .A1(mai_mai_n546_), .B0(mai_mai_n936_), .B1(mai_mai_n935_), .Y(mai_mai_n938_));
  NA4        m0910(.A(mai_mai_n938_), .B(mai_mai_n934_), .C(mai_mai_n933_), .D(mai_mai_n445_), .Y(mai_mai_n939_));
  AOI210     m0911(.A0(mai_mai_n233_), .A1(mai_mai_n342_), .B0(mai_mai_n201_), .Y(mai_mai_n940_));
  OR2        m0912(.A(mai_mai_n940_), .B(mai_mai_n932_), .Y(mai_mai_n941_));
  AOI210     m0913(.A0(mai_mai_n339_), .A1(mai_mai_n393_), .B0(mai_mai_n215_), .Y(mai_mai_n942_));
  OAI210     m0914(.A0(mai_mai_n942_), .A1(mai_mai_n941_), .B0(mai_mai_n407_), .Y(mai_mai_n943_));
  NO2        m0915(.A(mai_mai_n641_), .B(mai_mai_n263_), .Y(mai_mai_n944_));
  NO2        m0916(.A(mai_mai_n590_), .B(mai_mai_n844_), .Y(mai_mai_n945_));
  AOI220     m0917(.A0(mai_mai_n945_), .A1(mai_mai_n571_), .B0(mai_mai_n822_), .B1(mai_mai_n944_), .Y(mai_mai_n946_));
  NO2        m0918(.A(mai_mai_n150_), .B(mai_mai_n237_), .Y(mai_mai_n947_));
  NA3        m0919(.A(mai_mai_n947_), .B(mai_mai_n240_), .C(i), .Y(mai_mai_n948_));
  NA3        m0920(.A(mai_mai_n948_), .B(mai_mai_n946_), .C(mai_mai_n943_), .Y(mai_mai_n949_));
  NA4        m0921(.A(mai_mai_n447_), .B(mai_mai_n441_), .C(mai_mai_n182_), .D(g), .Y(mai_mai_n950_));
  NO3        m0922(.A(mai_mai_n666_), .B(mai_mai_n93_), .C(mai_mai_n45_), .Y(mai_mai_n951_));
  NO4        m0923(.A(mai_mai_n951_), .B(mai_mai_n1523_), .C(mai_mai_n949_), .D(mai_mai_n939_), .Y(mai_mai_n952_));
  NO2        m0924(.A(mai_mai_n371_), .B(mai_mai_n370_), .Y(mai_mai_n953_));
  NA2        m0925(.A(mai_mai_n587_), .B(mai_mai_n73_), .Y(mai_mai_n954_));
  NA2        m0926(.A(mai_mai_n558_), .B(mai_mai_n144_), .Y(mai_mai_n955_));
  NOi21      m0927(.An(mai_mai_n34_), .B(mai_mai_n655_), .Y(mai_mai_n956_));
  AOI220     m0928(.A0(mai_mai_n956_), .A1(mai_mai_n955_), .B0(mai_mai_n954_), .B1(mai_mai_n953_), .Y(mai_mai_n957_));
  OAI210     m0929(.A0(mai_mai_n251_), .A1(mai_mai_n45_), .B0(mai_mai_n957_), .Y(mai_mai_n958_));
  NA2        m0930(.A(mai_mai_n439_), .B(mai_mai_n265_), .Y(mai_mai_n959_));
  NO3        m0931(.A(mai_mai_n823_), .B(mai_mai_n91_), .C(mai_mai_n412_), .Y(mai_mai_n960_));
  NAi31      m0932(.An(mai_mai_n960_), .B(mai_mai_n959_), .C(mai_mai_n323_), .Y(mai_mai_n961_));
  NO2        m0933(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n962_));
  NO2        m0934(.A(mai_mai_n506_), .B(mai_mai_n301_), .Y(mai_mai_n963_));
  NO2        m0935(.A(mai_mai_n963_), .B(mai_mai_n367_), .Y(mai_mai_n964_));
  NO2        m0936(.A(mai_mai_n964_), .B(mai_mai_n144_), .Y(mai_mai_n965_));
  NA2        m0937(.A(mai_mai_n633_), .B(mai_mai_n364_), .Y(mai_mai_n966_));
  OAI210     m0938(.A0(mai_mai_n735_), .A1(mai_mai_n966_), .B0(mai_mai_n368_), .Y(mai_mai_n967_));
  NO4        m0939(.A(mai_mai_n967_), .B(mai_mai_n965_), .C(mai_mai_n961_), .D(mai_mai_n958_), .Y(mai_mai_n968_));
  NA2        m0940(.A(mai_mai_n349_), .B(g), .Y(mai_mai_n969_));
  NA2        m0941(.A(mai_mai_n161_), .B(i), .Y(mai_mai_n970_));
  NA2        m0942(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n971_));
  OAI220     m0943(.A0(mai_mai_n971_), .A1(mai_mai_n200_), .B0(mai_mai_n970_), .B1(mai_mai_n93_), .Y(mai_mai_n972_));
  AOI210     m0944(.A0(mai_mai_n423_), .A1(mai_mai_n37_), .B0(mai_mai_n972_), .Y(mai_mai_n973_));
  NA2        m0945(.A(mai_mai_n558_), .B(mai_mai_n385_), .Y(mai_mai_n974_));
  AOI210     m0946(.A0(mai_mai_n974_), .A1(n), .B0(mai_mai_n557_), .Y(mai_mai_n975_));
  OAI220     m0947(.A0(mai_mai_n975_), .A1(mai_mai_n969_), .B0(mai_mai_n973_), .B1(mai_mai_n336_), .Y(mai_mai_n976_));
  NO2        m0948(.A(mai_mai_n661_), .B(mai_mai_n500_), .Y(mai_mai_n977_));
  NA3        m0949(.A(mai_mai_n346_), .B(mai_mai_n630_), .C(i), .Y(mai_mai_n978_));
  OAI210     m0950(.A0(mai_mai_n443_), .A1(mai_mai_n312_), .B0(mai_mai_n978_), .Y(mai_mai_n979_));
  OAI220     m0951(.A0(mai_mai_n979_), .A1(mai_mai_n977_), .B0(mai_mai_n680_), .B1(mai_mai_n760_), .Y(mai_mai_n980_));
  NA2        m0952(.A(mai_mai_n608_), .B(mai_mai_n114_), .Y(mai_mai_n981_));
  OR3        m0953(.A(mai_mai_n312_), .B(mai_mai_n438_), .C(f), .Y(mai_mai_n982_));
  NA3        m0954(.A(mai_mai_n328_), .B(mai_mai_n119_), .C(g), .Y(mai_mai_n983_));
  AOI210     m0955(.A0(mai_mai_n677_), .A1(mai_mai_n983_), .B0(m), .Y(mai_mai_n984_));
  OAI210     m0956(.A0(mai_mai_n984_), .A1(mai_mai_n936_), .B0(mai_mai_n327_), .Y(mai_mai_n985_));
  NA2        m0957(.A(mai_mai_n695_), .B(mai_mai_n882_), .Y(mai_mai_n986_));
  NA2        m0958(.A(mai_mai_n846_), .B(mai_mai_n444_), .Y(mai_mai_n987_));
  NA2        m0959(.A(mai_mai_n221_), .B(mai_mai_n79_), .Y(mai_mai_n988_));
  NA2        m0960(.A(mai_mai_n988_), .B(mai_mai_n982_), .Y(mai_mai_n989_));
  AOI220     m0961(.A0(mai_mai_n989_), .A1(mai_mai_n258_), .B0(mai_mai_n987_), .B1(mai_mai_n986_), .Y(mai_mai_n990_));
  NA3        m0962(.A(mai_mai_n990_), .B(mai_mai_n985_), .C(mai_mai_n980_), .Y(mai_mai_n991_));
  NA2        m0963(.A(mai_mai_n665_), .B(mai_mai_n90_), .Y(mai_mai_n992_));
  NO2        m0964(.A(mai_mai_n461_), .B(mai_mai_n215_), .Y(mai_mai_n993_));
  NA2        m0965(.A(mai_mai_n993_), .B(mai_mai_n386_), .Y(mai_mai_n994_));
  NA2        m0966(.A(mai_mai_n994_), .B(mai_mai_n992_), .Y(mai_mai_n995_));
  OAI210     m0967(.A0(mai_mai_n987_), .A1(mai_mai_n945_), .B0(mai_mai_n546_), .Y(mai_mai_n996_));
  AOI210     m0968(.A0(mai_mai_n424_), .A1(mai_mai_n416_), .B0(mai_mai_n823_), .Y(mai_mai_n997_));
  OAI210     m0969(.A0(mai_mai_n371_), .A1(mai_mai_n370_), .B0(mai_mai_n110_), .Y(mai_mai_n998_));
  AOI210     m0970(.A0(mai_mai_n998_), .A1(mai_mai_n538_), .B0(mai_mai_n997_), .Y(mai_mai_n999_));
  NA2        m0971(.A(mai_mai_n984_), .B(mai_mai_n935_), .Y(mai_mai_n1000_));
  NO3        m0972(.A(mai_mai_n896_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n1001_));
  AOI220     m0973(.A0(mai_mai_n1001_), .A1(mai_mai_n628_), .B0(mai_mai_n646_), .B1(mai_mai_n533_), .Y(mai_mai_n1002_));
  NA4        m0974(.A(mai_mai_n1002_), .B(mai_mai_n1000_), .C(mai_mai_n999_), .D(mai_mai_n996_), .Y(mai_mai_n1003_));
  NO4        m0975(.A(mai_mai_n1003_), .B(mai_mai_n995_), .C(mai_mai_n991_), .D(mai_mai_n976_), .Y(mai_mai_n1004_));
  NAi31      m0976(.An(mai_mai_n141_), .B(mai_mai_n425_), .C(n), .Y(mai_mai_n1005_));
  NO2        m0977(.A(mai_mai_n127_), .B(mai_mai_n344_), .Y(mai_mai_n1006_));
  NO2        m0978(.A(mai_mai_n1006_), .B(mai_mai_n1005_), .Y(mai_mai_n1007_));
  NO3        m0979(.A(mai_mai_n273_), .B(mai_mai_n141_), .C(mai_mai_n412_), .Y(mai_mai_n1008_));
  AOI210     m0980(.A0(mai_mai_n1008_), .A1(mai_mai_n501_), .B0(mai_mai_n1007_), .Y(mai_mai_n1009_));
  INV        m0981(.A(mai_mai_n1009_), .Y(mai_mai_n1010_));
  NA2        m0982(.A(mai_mai_n230_), .B(mai_mai_n172_), .Y(mai_mai_n1011_));
  NO3        m0983(.A(mai_mai_n310_), .B(mai_mai_n447_), .C(mai_mai_n176_), .Y(mai_mai_n1012_));
  NOi31      m0984(.An(mai_mai_n1011_), .B(mai_mai_n1012_), .C(mai_mai_n215_), .Y(mai_mai_n1013_));
  NAi21      m0985(.An(mai_mai_n558_), .B(mai_mai_n993_), .Y(mai_mai_n1014_));
  NA2        m0986(.A(mai_mai_n442_), .B(mai_mai_n882_), .Y(mai_mai_n1015_));
  NO3        m0987(.A(mai_mai_n443_), .B(mai_mai_n312_), .C(mai_mai_n75_), .Y(mai_mai_n1016_));
  AOI220     m0988(.A0(mai_mai_n1016_), .A1(mai_mai_n1015_), .B0(mai_mai_n484_), .B1(g), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n1017_), .B(mai_mai_n1014_), .Y(mai_mai_n1018_));
  OAI220     m0990(.A0(mai_mai_n1005_), .A1(mai_mai_n233_), .B0(mai_mai_n978_), .B1(mai_mai_n603_), .Y(mai_mai_n1019_));
  NO2        m0991(.A(mai_mai_n662_), .B(mai_mai_n381_), .Y(mai_mai_n1020_));
  NA2        m0992(.A(mai_mai_n940_), .B(mai_mai_n931_), .Y(mai_mai_n1021_));
  NO3        m0993(.A(mai_mai_n547_), .B(mai_mai_n148_), .C(mai_mai_n214_), .Y(mai_mai_n1022_));
  OAI210     m0994(.A0(mai_mai_n1022_), .A1(mai_mai_n528_), .B0(mai_mai_n382_), .Y(mai_mai_n1023_));
  OAI220     m0995(.A0(mai_mai_n937_), .A1(mai_mai_n945_), .B0(mai_mai_n548_), .B1(mai_mai_n432_), .Y(mai_mai_n1024_));
  NA4        m0996(.A(mai_mai_n1024_), .B(mai_mai_n1023_), .C(mai_mai_n1021_), .D(mai_mai_n622_), .Y(mai_mai_n1025_));
  OAI210     m0997(.A0(mai_mai_n940_), .A1(mai_mai_n932_), .B0(mai_mai_n1011_), .Y(mai_mai_n1026_));
  NA3        m0998(.A(mai_mai_n974_), .B(mai_mai_n489_), .C(mai_mai_n46_), .Y(mai_mai_n1027_));
  AOI210     m0999(.A0(mai_mai_n384_), .A1(mai_mai_n382_), .B0(mai_mai_n335_), .Y(mai_mai_n1028_));
  NA4        m1000(.A(mai_mai_n1028_), .B(mai_mai_n1027_), .C(mai_mai_n1026_), .D(mai_mai_n274_), .Y(mai_mai_n1029_));
  OR4        m1001(.A(mai_mai_n1029_), .B(mai_mai_n1025_), .C(mai_mai_n1020_), .D(mai_mai_n1019_), .Y(mai_mai_n1030_));
  NO4        m1002(.A(mai_mai_n1030_), .B(mai_mai_n1018_), .C(mai_mai_n1013_), .D(mai_mai_n1010_), .Y(mai_mai_n1031_));
  NA4        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1004_), .C(mai_mai_n968_), .D(mai_mai_n952_), .Y(mai13));
  AN2        m1004(.A(c), .B(b), .Y(mai_mai_n1033_));
  NA3        m1005(.A(mai_mai_n250_), .B(mai_mai_n1033_), .C(m), .Y(mai_mai_n1034_));
  NA2        m1006(.A(mai_mai_n499_), .B(f), .Y(mai_mai_n1035_));
  NO4        m1007(.A(mai_mai_n1035_), .B(mai_mai_n1034_), .C(j), .D(mai_mai_n583_), .Y(mai_mai_n1036_));
  NA2        m1008(.A(mai_mai_n265_), .B(mai_mai_n1033_), .Y(mai_mai_n1037_));
  NO4        m1009(.A(mai_mai_n1037_), .B(mai_mai_n1035_), .C(mai_mai_n970_), .D(a), .Y(mai_mai_n1038_));
  NAi32      m1010(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n140_), .B(mai_mai_n45_), .Y(mai_mai_n1040_));
  NO4        m1012(.A(mai_mai_n1040_), .B(mai_mai_n1039_), .C(mai_mai_n590_), .D(mai_mai_n309_), .Y(mai_mai_n1041_));
  NA2        m1013(.A(mai_mai_n669_), .B(mai_mai_n224_), .Y(mai_mai_n1042_));
  NA2        m1014(.A(mai_mai_n415_), .B(mai_mai_n214_), .Y(mai_mai_n1043_));
  AN2        m1015(.A(d), .B(c), .Y(mai_mai_n1044_));
  NA2        m1016(.A(mai_mai_n1044_), .B(mai_mai_n117_), .Y(mai_mai_n1045_));
  NO4        m1017(.A(mai_mai_n1045_), .B(mai_mai_n1043_), .C(mai_mai_n177_), .D(mai_mai_n168_), .Y(mai_mai_n1046_));
  NA2        m1018(.A(mai_mai_n499_), .B(c), .Y(mai_mai_n1047_));
  NO4        m1019(.A(mai_mai_n1040_), .B(mai_mai_n586_), .C(mai_mai_n1047_), .D(mai_mai_n309_), .Y(mai_mai_n1048_));
  AO210      m1020(.A0(mai_mai_n1046_), .A1(mai_mai_n1042_), .B0(mai_mai_n1048_), .Y(mai_mai_n1049_));
  OR4        m1021(.A(mai_mai_n1049_), .B(mai_mai_n1041_), .C(mai_mai_n1038_), .D(mai_mai_n1036_), .Y(mai_mai_n1050_));
  NAi32      m1022(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1051_));
  NO2        m1023(.A(mai_mai_n1051_), .B(mai_mai_n145_), .Y(mai_mai_n1052_));
  NA2        m1024(.A(mai_mai_n1052_), .B(g), .Y(mai_mai_n1053_));
  OR3        m1025(.A(mai_mai_n224_), .B(mai_mai_n177_), .C(mai_mai_n168_), .Y(mai_mai_n1054_));
  NO2        m1026(.A(mai_mai_n1054_), .B(mai_mai_n1053_), .Y(mai_mai_n1055_));
  NO2        m1027(.A(mai_mai_n1047_), .B(mai_mai_n309_), .Y(mai_mai_n1056_));
  NO2        m1028(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1057_));
  NA2        m1029(.A(mai_mai_n632_), .B(mai_mai_n1057_), .Y(mai_mai_n1058_));
  NOi21      m1030(.An(mai_mai_n1056_), .B(mai_mai_n1058_), .Y(mai_mai_n1059_));
  NO2        m1031(.A(mai_mai_n764_), .B(mai_mai_n113_), .Y(mai_mai_n1060_));
  NOi41      m1032(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1061_));
  NA2        m1033(.A(mai_mai_n1061_), .B(mai_mai_n1060_), .Y(mai_mai_n1062_));
  NO2        m1034(.A(mai_mai_n1062_), .B(mai_mai_n1053_), .Y(mai_mai_n1063_));
  OR3        m1035(.A(e), .B(d), .C(c), .Y(mai_mai_n1064_));
  NA3        m1036(.A(k), .B(j), .C(i), .Y(mai_mai_n1065_));
  NO3        m1037(.A(mai_mai_n1065_), .B(mai_mai_n309_), .C(mai_mai_n92_), .Y(mai_mai_n1066_));
  NOi21      m1038(.An(mai_mai_n1066_), .B(mai_mai_n1064_), .Y(mai_mai_n1067_));
  OR4        m1039(.A(mai_mai_n1067_), .B(mai_mai_n1063_), .C(mai_mai_n1059_), .D(mai_mai_n1055_), .Y(mai_mai_n1068_));
  NA3        m1040(.A(mai_mai_n469_), .B(mai_mai_n338_), .C(mai_mai_n56_), .Y(mai_mai_n1069_));
  NO2        m1041(.A(mai_mai_n1069_), .B(mai_mai_n1058_), .Y(mai_mai_n1070_));
  NO4        m1042(.A(mai_mai_n1069_), .B(mai_mai_n586_), .C(mai_mai_n452_), .D(mai_mai_n45_), .Y(mai_mai_n1071_));
  NO2        m1043(.A(f), .B(c), .Y(mai_mai_n1072_));
  NOi21      m1044(.An(mai_mai_n1072_), .B(mai_mai_n446_), .Y(mai_mai_n1073_));
  NA2        m1045(.A(mai_mai_n1073_), .B(mai_mai_n59_), .Y(mai_mai_n1074_));
  OR2        m1046(.A(k), .B(i), .Y(mai_mai_n1075_));
  NO3        m1047(.A(mai_mai_n1075_), .B(mai_mai_n244_), .C(l), .Y(mai_mai_n1076_));
  NOi31      m1048(.An(mai_mai_n1076_), .B(mai_mai_n1074_), .C(j), .Y(mai_mai_n1077_));
  OR3        m1049(.A(mai_mai_n1077_), .B(mai_mai_n1071_), .C(mai_mai_n1070_), .Y(mai_mai_n1078_));
  OR3        m1050(.A(mai_mai_n1078_), .B(mai_mai_n1068_), .C(mai_mai_n1050_), .Y(mai02));
  OR2        m1051(.A(l), .B(k), .Y(mai_mai_n1080_));
  OR3        m1052(.A(h), .B(g), .C(f), .Y(mai_mai_n1081_));
  OR3        m1053(.A(n), .B(m), .C(i), .Y(mai_mai_n1082_));
  NO4        m1054(.A(mai_mai_n1082_), .B(mai_mai_n1081_), .C(mai_mai_n1080_), .D(mai_mai_n1064_), .Y(mai_mai_n1083_));
  NOi31      m1055(.An(e), .B(d), .C(c), .Y(mai_mai_n1084_));
  AOI210     m1056(.A0(mai_mai_n1066_), .A1(mai_mai_n1084_), .B0(mai_mai_n1041_), .Y(mai_mai_n1085_));
  AN3        m1057(.A(g), .B(f), .C(c), .Y(mai_mai_n1086_));
  NA3        m1058(.A(mai_mai_n1086_), .B(mai_mai_n469_), .C(h), .Y(mai_mai_n1087_));
  OR2        m1059(.A(mai_mai_n1065_), .B(mai_mai_n309_), .Y(mai_mai_n1088_));
  OR2        m1060(.A(mai_mai_n1088_), .B(mai_mai_n1087_), .Y(mai_mai_n1089_));
  NO3        m1061(.A(mai_mai_n1069_), .B(mai_mai_n1040_), .C(mai_mai_n586_), .Y(mai_mai_n1090_));
  NO2        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1055_), .Y(mai_mai_n1091_));
  NA3        m1063(.A(l), .B(k), .C(j), .Y(mai_mai_n1092_));
  NA2        m1064(.A(i), .B(h), .Y(mai_mai_n1093_));
  NO3        m1065(.A(mai_mai_n1093_), .B(mai_mai_n1092_), .C(mai_mai_n133_), .Y(mai_mai_n1094_));
  NO3        m1066(.A(mai_mai_n142_), .B(mai_mai_n283_), .C(mai_mai_n215_), .Y(mai_mai_n1095_));
  AOI210     m1067(.A0(mai_mai_n1095_), .A1(mai_mai_n1094_), .B0(mai_mai_n1059_), .Y(mai_mai_n1096_));
  NA3        m1068(.A(c), .B(b), .C(a), .Y(mai_mai_n1097_));
  NO3        m1069(.A(mai_mai_n1097_), .B(mai_mai_n903_), .C(mai_mai_n214_), .Y(mai_mai_n1098_));
  NO4        m1070(.A(mai_mai_n1065_), .B(mai_mai_n301_), .C(mai_mai_n49_), .D(mai_mai_n113_), .Y(mai_mai_n1099_));
  AOI210     m1071(.A0(mai_mai_n1099_), .A1(mai_mai_n1098_), .B0(mai_mai_n1070_), .Y(mai_mai_n1100_));
  AN4        m1072(.A(mai_mai_n1100_), .B(mai_mai_n1096_), .C(mai_mai_n1091_), .D(mai_mai_n1089_), .Y(mai_mai_n1101_));
  NO2        m1073(.A(mai_mai_n1045_), .B(mai_mai_n1043_), .Y(mai_mai_n1102_));
  NA2        m1074(.A(mai_mai_n1062_), .B(mai_mai_n1054_), .Y(mai_mai_n1103_));
  AOI210     m1075(.A0(mai_mai_n1103_), .A1(mai_mai_n1102_), .B0(mai_mai_n1036_), .Y(mai_mai_n1104_));
  NAi41      m1076(.An(mai_mai_n1083_), .B(mai_mai_n1104_), .C(mai_mai_n1101_), .D(mai_mai_n1085_), .Y(mai03));
  INV        m1077(.A(mai_mai_n998_), .Y(mai_mai_n1106_));
  NOi41      m1078(.An(mai_mai_n809_), .B(mai_mai_n857_), .C(mai_mai_n847_), .D(mai_mai_n717_), .Y(mai_mai_n1107_));
  OAI220     m1079(.A0(mai_mai_n1107_), .A1(mai_mai_n695_), .B0(mai_mai_n1106_), .B1(mai_mai_n587_), .Y(mai_mai_n1108_));
  NOi31      m1080(.An(i), .B(k), .C(j), .Y(mai_mai_n1109_));
  NA4        m1081(.A(mai_mai_n1109_), .B(mai_mai_n1084_), .C(mai_mai_n346_), .D(mai_mai_n338_), .Y(mai_mai_n1110_));
  OAI210     m1082(.A0(mai_mai_n823_), .A1(mai_mai_n426_), .B0(mai_mai_n1110_), .Y(mai_mai_n1111_));
  NOi31      m1083(.An(m), .B(n), .C(f), .Y(mai_mai_n1112_));
  NA2        m1084(.A(mai_mai_n1112_), .B(mai_mai_n51_), .Y(mai_mai_n1113_));
  AN2        m1085(.A(e), .B(c), .Y(mai_mai_n1114_));
  NA2        m1086(.A(mai_mai_n1114_), .B(a), .Y(mai_mai_n1115_));
  OAI220     m1087(.A0(mai_mai_n1115_), .A1(mai_mai_n1113_), .B0(mai_mai_n890_), .B1(mai_mai_n431_), .Y(mai_mai_n1116_));
  NA2        m1088(.A(mai_mai_n509_), .B(l), .Y(mai_mai_n1117_));
  NOi31      m1089(.An(mai_mai_n867_), .B(mai_mai_n1034_), .C(mai_mai_n1117_), .Y(mai_mai_n1118_));
  NO4        m1090(.A(mai_mai_n1118_), .B(mai_mai_n1116_), .C(mai_mai_n1111_), .D(mai_mai_n997_), .Y(mai_mai_n1119_));
  NO2        m1091(.A(mai_mai_n283_), .B(a), .Y(mai_mai_n1120_));
  INV        m1092(.A(mai_mai_n1041_), .Y(mai_mai_n1121_));
  NO2        m1093(.A(mai_mai_n1093_), .B(mai_mai_n487_), .Y(mai_mai_n1122_));
  NO2        m1094(.A(mai_mai_n89_), .B(g), .Y(mai_mai_n1123_));
  AOI210     m1095(.A0(mai_mai_n1123_), .A1(mai_mai_n1122_), .B0(mai_mai_n1076_), .Y(mai_mai_n1124_));
  OR2        m1096(.A(mai_mai_n1124_), .B(mai_mai_n1074_), .Y(mai_mai_n1125_));
  NA3        m1097(.A(mai_mai_n1125_), .B(mai_mai_n1121_), .C(mai_mai_n1119_), .Y(mai_mai_n1126_));
  NO4        m1098(.A(mai_mai_n1126_), .B(mai_mai_n1108_), .C(mai_mai_n824_), .D(mai_mai_n570_), .Y(mai_mai_n1127_));
  NA2        m1099(.A(c), .B(b), .Y(mai_mai_n1128_));
  NO2        m1100(.A(mai_mai_n705_), .B(mai_mai_n1128_), .Y(mai_mai_n1129_));
  OAI210     m1101(.A0(mai_mai_n865_), .A1(mai_mai_n838_), .B0(mai_mai_n419_), .Y(mai_mai_n1130_));
  OAI210     m1102(.A0(mai_mai_n1130_), .A1(mai_mai_n866_), .B0(mai_mai_n1129_), .Y(mai_mai_n1131_));
  NAi21      m1103(.An(mai_mai_n427_), .B(mai_mai_n1129_), .Y(mai_mai_n1132_));
  NA3        m1104(.A(mai_mai_n432_), .B(mai_mai_n563_), .C(f), .Y(mai_mai_n1133_));
  OAI210     m1105(.A0(mai_mai_n552_), .A1(mai_mai_n39_), .B0(mai_mai_n1120_), .Y(mai_mai_n1134_));
  NA3        m1106(.A(mai_mai_n1134_), .B(mai_mai_n1133_), .C(mai_mai_n1132_), .Y(mai_mai_n1135_));
  NA2        m1107(.A(mai_mai_n261_), .B(mai_mai_n120_), .Y(mai_mai_n1136_));
  OAI210     m1108(.A0(mai_mai_n1136_), .A1(mai_mai_n287_), .B0(g), .Y(mai_mai_n1137_));
  NAi21      m1109(.An(f), .B(d), .Y(mai_mai_n1138_));
  NO2        m1110(.A(mai_mai_n1138_), .B(mai_mai_n1097_), .Y(mai_mai_n1139_));
  INV        m1111(.A(mai_mai_n1139_), .Y(mai_mai_n1140_));
  AOI210     m1112(.A0(mai_mai_n1137_), .A1(mai_mai_n293_), .B0(mai_mai_n1140_), .Y(mai_mai_n1141_));
  AOI210     m1113(.A0(mai_mai_n1141_), .A1(mai_mai_n114_), .B0(mai_mai_n1135_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n472_), .B(mai_mai_n471_), .Y(mai_mai_n1143_));
  NO2        m1115(.A(mai_mai_n183_), .B(mai_mai_n237_), .Y(mai_mai_n1144_));
  NA2        m1116(.A(mai_mai_n1144_), .B(m), .Y(mai_mai_n1145_));
  NA3        m1117(.A(mai_mai_n920_), .B(mai_mai_n1117_), .C(mai_mai_n475_), .Y(mai_mai_n1146_));
  OAI210     m1118(.A0(mai_mai_n1146_), .A1(mai_mai_n313_), .B0(mai_mai_n473_), .Y(mai_mai_n1147_));
  AOI210     m1119(.A0(mai_mai_n1147_), .A1(mai_mai_n1143_), .B0(mai_mai_n1145_), .Y(mai_mai_n1148_));
  NA2        m1120(.A(mai_mai_n565_), .B(mai_mai_n414_), .Y(mai_mai_n1149_));
  NA2        m1121(.A(mai_mai_n157_), .B(mai_mai_n33_), .Y(mai_mai_n1150_));
  AOI210     m1122(.A0(mai_mai_n966_), .A1(mai_mai_n1150_), .B0(mai_mai_n215_), .Y(mai_mai_n1151_));
  NA2        m1123(.A(mai_mai_n1151_), .B(mai_mai_n1139_), .Y(mai_mai_n1152_));
  NO2        m1124(.A(mai_mai_n375_), .B(mai_mai_n374_), .Y(mai_mai_n1153_));
  AOI210     m1125(.A0(mai_mai_n1144_), .A1(mai_mai_n434_), .B0(mai_mai_n960_), .Y(mai_mai_n1154_));
  NAi41      m1126(.An(mai_mai_n1153_), .B(mai_mai_n1154_), .C(mai_mai_n1152_), .D(mai_mai_n1149_), .Y(mai_mai_n1155_));
  NO2        m1127(.A(mai_mai_n1155_), .B(mai_mai_n1148_), .Y(mai_mai_n1156_));
  NA4        m1128(.A(mai_mai_n1156_), .B(mai_mai_n1142_), .C(mai_mai_n1131_), .D(mai_mai_n1127_), .Y(mai00));
  AOI210     m1129(.A0(mai_mai_n300_), .A1(mai_mai_n215_), .B0(mai_mai_n276_), .Y(mai_mai_n1158_));
  NO2        m1130(.A(mai_mai_n1158_), .B(mai_mai_n579_), .Y(mai_mai_n1159_));
  AOI210     m1131(.A0(mai_mai_n900_), .A1(mai_mai_n947_), .B0(mai_mai_n1111_), .Y(mai_mai_n1160_));
  NO2        m1132(.A(mai_mai_n1090_), .B(mai_mai_n960_), .Y(mai_mai_n1161_));
  NA3        m1133(.A(mai_mai_n1161_), .B(mai_mai_n1160_), .C(mai_mai_n999_), .Y(mai_mai_n1162_));
  NA2        m1134(.A(mai_mai_n511_), .B(f), .Y(mai_mai_n1163_));
  OAI210     m1135(.A0(mai_mai_n1006_), .A1(mai_mai_n40_), .B0(mai_mai_n648_), .Y(mai_mai_n1164_));
  NA3        m1136(.A(mai_mai_n1164_), .B(mai_mai_n257_), .C(n), .Y(mai_mai_n1165_));
  AOI210     m1137(.A0(mai_mai_n1165_), .A1(mai_mai_n1163_), .B0(mai_mai_n1045_), .Y(mai_mai_n1166_));
  NO4        m1138(.A(mai_mai_n1166_), .B(mai_mai_n1162_), .C(mai_mai_n1159_), .D(mai_mai_n1068_), .Y(mai_mai_n1167_));
  NA3        m1139(.A(mai_mai_n167_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1168_));
  NA3        m1140(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1169_));
  NOi31      m1141(.An(n), .B(m), .C(i), .Y(mai_mai_n1170_));
  NA3        m1142(.A(mai_mai_n1170_), .B(mai_mai_n651_), .C(mai_mai_n51_), .Y(mai_mai_n1171_));
  OAI210     m1143(.A0(mai_mai_n1169_), .A1(mai_mai_n1168_), .B0(mai_mai_n1171_), .Y(mai_mai_n1172_));
  NO3        m1144(.A(mai_mai_n1172_), .B(mai_mai_n1153_), .C(mai_mai_n923_), .Y(mai_mai_n1173_));
  NO4        m1145(.A(mai_mai_n490_), .B(mai_mai_n357_), .C(mai_mai_n1128_), .D(mai_mai_n59_), .Y(mai_mai_n1174_));
  OR2        m1146(.A(mai_mai_n388_), .B(mai_mai_n135_), .Y(mai_mai_n1175_));
  NO2        m1147(.A(h), .B(g), .Y(mai_mai_n1176_));
  NA4        m1148(.A(mai_mai_n501_), .B(mai_mai_n469_), .C(mai_mai_n1176_), .D(mai_mai_n1033_), .Y(mai_mai_n1177_));
  AOI220     m1149(.A0(mai_mai_n320_), .A1(mai_mai_n248_), .B0(mai_mai_n178_), .B1(mai_mai_n147_), .Y(mai_mai_n1178_));
  NA3        m1150(.A(mai_mai_n1178_), .B(mai_mai_n1177_), .C(mai_mai_n1175_), .Y(mai_mai_n1179_));
  NO3        m1151(.A(mai_mai_n1179_), .B(mai_mai_n1174_), .C(mai_mai_n267_), .Y(mai_mai_n1180_));
  NO2        m1152(.A(mai_mai_n239_), .B(mai_mai_n182_), .Y(mai_mai_n1181_));
  NA2        m1153(.A(mai_mai_n1181_), .B(mai_mai_n432_), .Y(mai_mai_n1182_));
  NA3        m1154(.A(mai_mai_n180_), .B(mai_mai_n113_), .C(g), .Y(mai_mai_n1183_));
  NA3        m1155(.A(mai_mai_n469_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1184_));
  NOi31      m1156(.An(mai_mai_n875_), .B(mai_mai_n1184_), .C(mai_mai_n1183_), .Y(mai_mai_n1185_));
  NAi31      m1157(.An(mai_mai_n185_), .B(mai_mai_n863_), .C(mai_mai_n469_), .Y(mai_mai_n1186_));
  NAi31      m1158(.An(mai_mai_n1185_), .B(mai_mai_n1186_), .C(mai_mai_n1182_), .Y(mai_mai_n1187_));
  NO2        m1159(.A(mai_mai_n275_), .B(mai_mai_n75_), .Y(mai_mai_n1188_));
  NO3        m1160(.A(mai_mai_n431_), .B(mai_mai_n834_), .C(n), .Y(mai_mai_n1189_));
  AOI210     m1161(.A0(mai_mai_n1189_), .A1(mai_mai_n1188_), .B0(mai_mai_n1083_), .Y(mai_mai_n1190_));
  NAi31      m1162(.An(mai_mai_n1048_), .B(mai_mai_n1190_), .C(mai_mai_n74_), .Y(mai_mai_n1191_));
  NO4        m1163(.A(mai_mai_n1191_), .B(mai_mai_n1187_), .C(mai_mai_n325_), .D(mai_mai_n521_), .Y(mai_mai_n1192_));
  AN3        m1164(.A(mai_mai_n1192_), .B(mai_mai_n1180_), .C(mai_mai_n1173_), .Y(mai_mai_n1193_));
  NA2        m1165(.A(mai_mai_n538_), .B(mai_mai_n102_), .Y(mai_mai_n1194_));
  NA3        m1166(.A(mai_mai_n1112_), .B(mai_mai_n608_), .C(mai_mai_n468_), .Y(mai_mai_n1195_));
  NA4        m1167(.A(mai_mai_n1195_), .B(mai_mai_n566_), .C(mai_mai_n1194_), .D(mai_mai_n242_), .Y(mai_mai_n1196_));
  OAI210     m1168(.A0(mai_mai_n467_), .A1(mai_mai_n121_), .B0(mai_mai_n868_), .Y(mai_mai_n1197_));
  AOI220     m1169(.A0(mai_mai_n1197_), .A1(mai_mai_n1146_), .B0(mai_mai_n565_), .B1(mai_mai_n414_), .Y(mai_mai_n1198_));
  OR4        m1170(.A(mai_mai_n1045_), .B(mai_mai_n273_), .C(mai_mai_n222_), .D(e), .Y(mai_mai_n1199_));
  NA2        m1171(.A(n), .B(e), .Y(mai_mai_n1200_));
  NO2        m1172(.A(mai_mai_n1200_), .B(mai_mai_n145_), .Y(mai_mai_n1201_));
  NA2        m1173(.A(mai_mai_n1199_), .B(mai_mai_n1198_), .Y(mai_mai_n1202_));
  AOI210     m1174(.A0(mai_mai_n1201_), .A1(mai_mai_n854_), .B0(mai_mai_n824_), .Y(mai_mai_n1203_));
  AOI220     m1175(.A0(mai_mai_n956_), .A1(mai_mai_n578_), .B0(mai_mai_n651_), .B1(mai_mai_n245_), .Y(mai_mai_n1204_));
  NO2        m1176(.A(mai_mai_n68_), .B(h), .Y(mai_mai_n1205_));
  NO3        m1177(.A(mai_mai_n1045_), .B(mai_mai_n1043_), .C(mai_mai_n727_), .Y(mai_mai_n1206_));
  NO2        m1178(.A(mai_mai_n1080_), .B(mai_mai_n133_), .Y(mai_mai_n1207_));
  AN2        m1179(.A(mai_mai_n1207_), .B(mai_mai_n1095_), .Y(mai_mai_n1208_));
  OAI210     m1180(.A0(mai_mai_n1208_), .A1(mai_mai_n1206_), .B0(mai_mai_n1205_), .Y(mai_mai_n1209_));
  NA4        m1181(.A(mai_mai_n1209_), .B(mai_mai_n1204_), .C(mai_mai_n1203_), .D(mai_mai_n870_), .Y(mai_mai_n1210_));
  NO4        m1182(.A(mai_mai_n1210_), .B(mai_mai_n1202_), .C(mai_mai_n296_), .D(mai_mai_n1196_), .Y(mai_mai_n1211_));
  NA2        m1183(.A(mai_mai_n839_), .B(mai_mai_n759_), .Y(mai_mai_n1212_));
  NA4        m1184(.A(mai_mai_n1212_), .B(mai_mai_n1211_), .C(mai_mai_n1193_), .D(mai_mai_n1167_), .Y(mai01));
  AN2        m1185(.A(mai_mai_n1023_), .B(mai_mai_n1021_), .Y(mai_mai_n1214_));
  NO3        m1186(.A(mai_mai_n805_), .B(mai_mai_n797_), .C(mai_mai_n281_), .Y(mai_mai_n1215_));
  NO2        m1187(.A(mai_mai_n592_), .B(mai_mai_n290_), .Y(mai_mai_n1216_));
  OAI210     m1188(.A0(mai_mai_n1216_), .A1(mai_mai_n398_), .B0(i), .Y(mai_mai_n1217_));
  NA3        m1189(.A(mai_mai_n1217_), .B(mai_mai_n1215_), .C(mai_mai_n1214_), .Y(mai_mai_n1218_));
  NA2        m1190(.A(mai_mai_n558_), .B(mai_mai_n272_), .Y(mai_mai_n1219_));
  NA2        m1191(.A(mai_mai_n963_), .B(mai_mai_n1219_), .Y(mai_mai_n1220_));
  NA3        m1192(.A(mai_mai_n1220_), .B(mai_mai_n916_), .C(mai_mai_n337_), .Y(mai_mai_n1221_));
  NA2        m1193(.A(mai_mai_n45_), .B(f), .Y(mai_mai_n1222_));
  NA2        m1194(.A(mai_mai_n712_), .B(mai_mai_n97_), .Y(mai_mai_n1223_));
  OAI220     m1195(.A0(mai_mai_n1223_), .A1(mai_mai_n1222_), .B0(mai_mai_n354_), .B1(mai_mai_n285_), .Y(mai_mai_n1224_));
  NO2        m1196(.A(mai_mai_n784_), .B(mai_mai_n603_), .Y(mai_mai_n1225_));
  AOI210     m1197(.A0(mai_mai_n1224_), .A1(mai_mai_n637_), .B0(mai_mai_n1225_), .Y(mai_mai_n1226_));
  NA2        m1198(.A(mai_mai_n119_), .B(l), .Y(mai_mai_n1227_));
  NAi31      m1199(.An(mai_mai_n160_), .B(mai_mai_n1226_), .C(mai_mai_n899_), .Y(mai_mai_n1228_));
  NO3        m1200(.A(mai_mai_n785_), .B(mai_mai_n679_), .C(mai_mai_n514_), .Y(mai_mai_n1229_));
  OR2        m1201(.A(mai_mai_n195_), .B(mai_mai_n193_), .Y(mai_mai_n1230_));
  NA3        m1202(.A(mai_mai_n1230_), .B(mai_mai_n1229_), .C(mai_mai_n138_), .Y(mai_mai_n1231_));
  NO4        m1203(.A(mai_mai_n1231_), .B(mai_mai_n1228_), .C(mai_mai_n1221_), .D(mai_mai_n1218_), .Y(mai_mai_n1232_));
  INV        m1204(.A(mai_mai_n207_), .Y(mai_mai_n1233_));
  OAI210     m1205(.A0(mai_mai_n1233_), .A1(mai_mai_n303_), .B0(mai_mai_n533_), .Y(mai_mai_n1234_));
  NA2        m1206(.A(mai_mai_n541_), .B(mai_mai_n400_), .Y(mai_mai_n1235_));
  NA2        m1207(.A(mai_mai_n76_), .B(i), .Y(mai_mai_n1236_));
  AOI210     m1208(.A0(mai_mai_n591_), .A1(mai_mai_n585_), .B0(mai_mai_n1236_), .Y(mai_mai_n1237_));
  NOi21      m1209(.An(mai_mai_n567_), .B(mai_mai_n582_), .Y(mai_mai_n1238_));
  AOI210     m1210(.A0(mai_mai_n1238_), .A1(mai_mai_n1235_), .B0(mai_mai_n1237_), .Y(mai_mai_n1239_));
  AOI210     m1211(.A0(mai_mai_n204_), .A1(mai_mai_n91_), .B0(mai_mai_n214_), .Y(mai_mai_n1240_));
  OAI210     m1212(.A0(mai_mai_n812_), .A1(mai_mai_n432_), .B0(mai_mai_n1240_), .Y(mai_mai_n1241_));
  AN3        m1213(.A(m), .B(l), .C(k), .Y(mai_mai_n1242_));
  OAI210     m1214(.A0(mai_mai_n360_), .A1(mai_mai_n34_), .B0(mai_mai_n1242_), .Y(mai_mai_n1243_));
  NA2        m1215(.A(mai_mai_n203_), .B(mai_mai_n34_), .Y(mai_mai_n1244_));
  AO210      m1216(.A0(mai_mai_n1244_), .A1(mai_mai_n1243_), .B0(mai_mai_n336_), .Y(mai_mai_n1245_));
  NA4        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1241_), .C(mai_mai_n1239_), .D(mai_mai_n1234_), .Y(mai_mai_n1246_));
  AOI210     m1218(.A0(mai_mai_n595_), .A1(mai_mai_n119_), .B0(mai_mai_n601_), .Y(mai_mai_n1247_));
  OAI210     m1219(.A0(mai_mai_n1227_), .A1(mai_mai_n594_), .B0(mai_mai_n1247_), .Y(mai_mai_n1248_));
  NA2        m1220(.A(mai_mai_n280_), .B(mai_mai_n195_), .Y(mai_mai_n1249_));
  OAI210     m1221(.A0(mai_mai_n1249_), .A1(mai_mai_n389_), .B0(mai_mai_n668_), .Y(mai_mai_n1250_));
  NO3        m1222(.A(mai_mai_n823_), .B(mai_mai_n204_), .C(mai_mai_n412_), .Y(mai_mai_n1251_));
  NO2        m1223(.A(mai_mai_n1251_), .B(mai_mai_n960_), .Y(mai_mai_n1252_));
  OAI210     m1224(.A0(mai_mai_n1224_), .A1(mai_mai_n330_), .B0(mai_mai_n680_), .Y(mai_mai_n1253_));
  NA4        m1225(.A(mai_mai_n1253_), .B(mai_mai_n1252_), .C(mai_mai_n1250_), .D(mai_mai_n788_), .Y(mai_mai_n1254_));
  NO3        m1226(.A(mai_mai_n1254_), .B(mai_mai_n1248_), .C(mai_mai_n1246_), .Y(mai_mai_n1255_));
  NA3        m1227(.A(mai_mai_n604_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1256_));
  NO2        m1228(.A(mai_mai_n1256_), .B(mai_mai_n204_), .Y(mai_mai_n1257_));
  AOI210     m1229(.A0(mai_mai_n507_), .A1(mai_mai_n58_), .B0(mai_mai_n1257_), .Y(mai_mai_n1258_));
  OR3        m1230(.A(mai_mai_n1223_), .B(mai_mai_n605_), .C(mai_mai_n1222_), .Y(mai_mai_n1259_));
  NA3        m1231(.A(mai_mai_n741_), .B(mai_mai_n76_), .C(i), .Y(mai_mai_n1260_));
  NO2        m1232(.A(mai_mai_n1260_), .B(mai_mai_n981_), .Y(mai_mai_n1261_));
  NO2        m1233(.A(mai_mai_n1261_), .B(mai_mai_n1172_), .Y(mai_mai_n1262_));
  NA4        m1234(.A(mai_mai_n1262_), .B(mai_mai_n1259_), .C(mai_mai_n1258_), .D(mai_mai_n758_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(mai_mai_n970_), .B(mai_mai_n232_), .Y(mai_mai_n1264_));
  NO2        m1236(.A(mai_mai_n971_), .B(mai_mai_n560_), .Y(mai_mai_n1265_));
  OAI210     m1237(.A0(mai_mai_n1265_), .A1(mai_mai_n1264_), .B0(mai_mai_n344_), .Y(mai_mai_n1266_));
  NO3        m1238(.A(mai_mai_n81_), .B(mai_mai_n301_), .C(mai_mai_n45_), .Y(mai_mai_n1267_));
  NA2        m1239(.A(mai_mai_n1267_), .B(mai_mai_n557_), .Y(mai_mai_n1268_));
  NA2        m1240(.A(mai_mai_n1268_), .B(mai_mai_n674_), .Y(mai_mai_n1269_));
  NO2        m1241(.A(mai_mai_n372_), .B(mai_mai_n73_), .Y(mai_mai_n1270_));
  AOI210     m1242(.A0(mai_mai_n732_), .A1(mai_mai_n619_), .B0(mai_mai_n1270_), .Y(mai_mai_n1271_));
  NA2        m1243(.A(mai_mai_n1267_), .B(mai_mai_n815_), .Y(mai_mai_n1272_));
  NA3        m1244(.A(mai_mai_n1272_), .B(mai_mai_n1271_), .C(mai_mai_n390_), .Y(mai_mai_n1273_));
  NOi41      m1245(.An(mai_mai_n1266_), .B(mai_mai_n1273_), .C(mai_mai_n1269_), .D(mai_mai_n1263_), .Y(mai_mai_n1274_));
  NO2        m1246(.A(mai_mai_n132_), .B(mai_mai_n45_), .Y(mai_mai_n1275_));
  NO2        m1247(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1276_));
  AO220      m1248(.A0(mai_mai_n1276_), .A1(mai_mai_n625_), .B0(mai_mai_n1275_), .B1(mai_mai_n710_), .Y(mai_mai_n1277_));
  NA2        m1249(.A(mai_mai_n1277_), .B(mai_mai_n344_), .Y(mai_mai_n1278_));
  NO3        m1250(.A(mai_mai_n1093_), .B(mai_mai_n177_), .C(mai_mai_n89_), .Y(mai_mai_n1279_));
  INV        m1251(.A(mai_mai_n1278_), .Y(mai_mai_n1280_));
  NO2        m1252(.A(mai_mai_n616_), .B(mai_mai_n615_), .Y(mai_mai_n1281_));
  NO4        m1253(.A(mai_mai_n1093_), .B(mai_mai_n1281_), .C(mai_mai_n175_), .D(mai_mai_n89_), .Y(mai_mai_n1282_));
  NO3        m1254(.A(mai_mai_n1282_), .B(mai_mai_n1280_), .C(mai_mai_n640_), .Y(mai_mai_n1283_));
  NA4        m1255(.A(mai_mai_n1283_), .B(mai_mai_n1274_), .C(mai_mai_n1255_), .D(mai_mai_n1232_), .Y(mai06));
  NO2        m1256(.A(mai_mai_n413_), .B(mai_mai_n564_), .Y(mai_mai_n1285_));
  NO2        m1257(.A(mai_mai_n734_), .B(i), .Y(mai_mai_n1286_));
  OAI210     m1258(.A0(mai_mai_n1286_), .A1(mai_mai_n268_), .B0(mai_mai_n1285_), .Y(mai_mai_n1287_));
  NO2        m1259(.A(mai_mai_n224_), .B(mai_mai_n103_), .Y(mai_mai_n1288_));
  OAI210     m1260(.A0(mai_mai_n1288_), .A1(mai_mai_n1279_), .B0(mai_mai_n386_), .Y(mai_mai_n1289_));
  NO3        m1261(.A(mai_mai_n599_), .B(mai_mai_n810_), .C(mai_mai_n602_), .Y(mai_mai_n1290_));
  OR2        m1262(.A(mai_mai_n1290_), .B(mai_mai_n890_), .Y(mai_mai_n1291_));
  NA4        m1263(.A(mai_mai_n1291_), .B(mai_mai_n1289_), .C(mai_mai_n1287_), .D(mai_mai_n1266_), .Y(mai_mai_n1292_));
  NO3        m1264(.A(mai_mai_n1292_), .B(mai_mai_n1269_), .C(mai_mai_n256_), .Y(mai_mai_n1293_));
  NO2        m1265(.A(mai_mai_n301_), .B(mai_mai_n45_), .Y(mai_mai_n1294_));
  AOI210     m1266(.A0(mai_mai_n1294_), .A1(mai_mai_n557_), .B0(mai_mai_n1264_), .Y(mai_mai_n1295_));
  AOI210     m1267(.A0(mai_mai_n1294_), .A1(mai_mai_n561_), .B0(mai_mai_n1277_), .Y(mai_mai_n1296_));
  AOI210     m1268(.A0(mai_mai_n1296_), .A1(mai_mai_n1295_), .B0(mai_mai_n342_), .Y(mai_mai_n1297_));
  OAI210     m1269(.A0(mai_mai_n91_), .A1(mai_mai_n40_), .B0(mai_mai_n678_), .Y(mai_mai_n1298_));
  NA2        m1270(.A(mai_mai_n1298_), .B(mai_mai_n644_), .Y(mai_mai_n1299_));
  NO2        m1271(.A(mai_mai_n517_), .B(mai_mai_n172_), .Y(mai_mai_n1300_));
  NOi21      m1272(.An(mai_mai_n137_), .B(mai_mai_n45_), .Y(mai_mai_n1301_));
  NO2        m1273(.A(mai_mai_n609_), .B(mai_mai_n1113_), .Y(mai_mai_n1302_));
  OAI210     m1274(.A0(mai_mai_n462_), .A1(mai_mai_n249_), .B0(mai_mai_n910_), .Y(mai_mai_n1303_));
  NO4        m1275(.A(mai_mai_n1303_), .B(mai_mai_n1302_), .C(mai_mai_n1301_), .D(mai_mai_n1300_), .Y(mai_mai_n1304_));
  OR2        m1276(.A(mai_mai_n600_), .B(mai_mai_n598_), .Y(mai_mai_n1305_));
  NO2        m1277(.A(mai_mai_n371_), .B(mai_mai_n136_), .Y(mai_mai_n1306_));
  AOI210     m1278(.A0(mai_mai_n1306_), .A1(mai_mai_n588_), .B0(mai_mai_n1305_), .Y(mai_mai_n1307_));
  NA3        m1279(.A(mai_mai_n1307_), .B(mai_mai_n1304_), .C(mai_mai_n1299_), .Y(mai_mai_n1308_));
  NO2        m1280(.A(mai_mai_n749_), .B(mai_mai_n370_), .Y(mai_mai_n1309_));
  NO3        m1281(.A(mai_mai_n680_), .B(mai_mai_n760_), .C(mai_mai_n637_), .Y(mai_mai_n1310_));
  NOi21      m1282(.An(mai_mai_n1309_), .B(mai_mai_n1310_), .Y(mai_mai_n1311_));
  AN2        m1283(.A(mai_mai_n956_), .B(mai_mai_n647_), .Y(mai_mai_n1312_));
  NO4        m1284(.A(mai_mai_n1312_), .B(mai_mai_n1311_), .C(mai_mai_n1308_), .D(mai_mai_n1297_), .Y(mai_mai_n1313_));
  NO2        m1285(.A(mai_mai_n804_), .B(mai_mai_n277_), .Y(mai_mai_n1314_));
  OAI220     m1286(.A0(mai_mai_n734_), .A1(mai_mai_n47_), .B0(mai_mai_n224_), .B1(mai_mai_n618_), .Y(mai_mai_n1315_));
  OAI210     m1287(.A0(mai_mai_n277_), .A1(c), .B0(mai_mai_n643_), .Y(mai_mai_n1316_));
  AOI220     m1288(.A0(mai_mai_n1316_), .A1(mai_mai_n1315_), .B0(mai_mai_n1314_), .B1(mai_mai_n268_), .Y(mai_mai_n1317_));
  OAI220     m1289(.A0(mai_mai_n702_), .A1(mai_mai_n249_), .B0(mai_mai_n513_), .B1(mai_mai_n517_), .Y(mai_mai_n1318_));
  OAI210     m1290(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1319_));
  NO3        m1291(.A(mai_mai_n1319_), .B(mai_mai_n597_), .C(j), .Y(mai_mai_n1320_));
  NOi21      m1292(.An(mai_mai_n1320_), .B(mai_mai_n672_), .Y(mai_mai_n1321_));
  NO3        m1293(.A(mai_mai_n1321_), .B(mai_mai_n1318_), .C(mai_mai_n1116_), .Y(mai_mai_n1322_));
  NA4        m1294(.A(mai_mai_n795_), .B(mai_mai_n794_), .C(mai_mai_n442_), .D(mai_mai_n882_), .Y(mai_mai_n1323_));
  NAi31      m1295(.An(mai_mai_n749_), .B(mai_mai_n1323_), .C(mai_mai_n203_), .Y(mai_mai_n1324_));
  NA4        m1296(.A(mai_mai_n1324_), .B(mai_mai_n1322_), .C(mai_mai_n1317_), .D(mai_mai_n1204_), .Y(mai_mai_n1325_));
  NOi31      m1297(.An(mai_mai_n1290_), .B(mai_mai_n466_), .C(mai_mai_n399_), .Y(mai_mai_n1326_));
  OR3        m1298(.A(mai_mai_n1326_), .B(mai_mai_n784_), .C(mai_mai_n544_), .Y(mai_mai_n1327_));
  OR3        m1299(.A(mai_mai_n374_), .B(mai_mai_n224_), .C(mai_mai_n618_), .Y(mai_mai_n1328_));
  INV        m1300(.A(mai_mai_n376_), .Y(mai_mai_n1329_));
  NA3        m1301(.A(mai_mai_n1329_), .B(mai_mai_n1328_), .C(mai_mai_n1327_), .Y(mai_mai_n1330_));
  AOI220     m1302(.A0(mai_mai_n1309_), .A1(mai_mai_n759_), .B0(mai_mai_n1306_), .B1(mai_mai_n238_), .Y(mai_mai_n1331_));
  AN2        m1303(.A(mai_mai_n932_), .B(mai_mai_n931_), .Y(mai_mai_n1332_));
  NO4        m1304(.A(mai_mai_n1332_), .B(mai_mai_n880_), .C(mai_mai_n503_), .D(mai_mai_n484_), .Y(mai_mai_n1333_));
  NA3        m1305(.A(mai_mai_n1333_), .B(mai_mai_n1331_), .C(mai_mai_n1272_), .Y(mai_mai_n1334_));
  NAi21      m1306(.An(j), .B(i), .Y(mai_mai_n1335_));
  NO4        m1307(.A(mai_mai_n1281_), .B(mai_mai_n1335_), .C(mai_mai_n446_), .D(mai_mai_n235_), .Y(mai_mai_n1336_));
  NO4        m1308(.A(mai_mai_n1336_), .B(mai_mai_n1334_), .C(mai_mai_n1330_), .D(mai_mai_n1325_), .Y(mai_mai_n1337_));
  NA4        m1309(.A(mai_mai_n1337_), .B(mai_mai_n1313_), .C(mai_mai_n1293_), .D(mai_mai_n1283_), .Y(mai07));
  NAi32      m1310(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1339_));
  NO3        m1311(.A(mai_mai_n1339_), .B(g), .C(f), .Y(mai_mai_n1340_));
  OAI210     m1312(.A0(mai_mai_n324_), .A1(mai_mai_n486_), .B0(mai_mai_n1340_), .Y(mai_mai_n1341_));
  NAi21      m1313(.An(f), .B(c), .Y(mai_mai_n1342_));
  OR2        m1314(.A(e), .B(d), .Y(mai_mai_n1343_));
  OAI220     m1315(.A0(mai_mai_n1343_), .A1(mai_mai_n1342_), .B0(mai_mai_n631_), .B1(mai_mai_n326_), .Y(mai_mai_n1344_));
  NA3        m1316(.A(mai_mai_n1344_), .B(mai_mai_n1057_), .C(mai_mai_n180_), .Y(mai_mai_n1345_));
  NOi31      m1317(.An(n), .B(m), .C(b), .Y(mai_mai_n1346_));
  NO3        m1318(.A(mai_mai_n133_), .B(mai_mai_n452_), .C(h), .Y(mai_mai_n1347_));
  NA2        m1319(.A(mai_mai_n1345_), .B(mai_mai_n1341_), .Y(mai_mai_n1348_));
  NOi41      m1320(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1349_));
  NOi21      m1321(.An(h), .B(k), .Y(mai_mai_n1350_));
  NO2        m1322(.A(k), .B(i), .Y(mai_mai_n1351_));
  NA3        m1323(.A(mai_mai_n1351_), .B(mai_mai_n898_), .C(mai_mai_n180_), .Y(mai_mai_n1352_));
  NA2        m1324(.A(mai_mai_n89_), .B(mai_mai_n45_), .Y(mai_mai_n1353_));
  NO2        m1325(.A(mai_mai_n1051_), .B(mai_mai_n446_), .Y(mai_mai_n1354_));
  NA3        m1326(.A(mai_mai_n1354_), .B(mai_mai_n1353_), .C(mai_mai_n215_), .Y(mai_mai_n1355_));
  NO2        m1327(.A(mai_mai_n1065_), .B(mai_mai_n309_), .Y(mai_mai_n1356_));
  NA2        m1328(.A(mai_mai_n545_), .B(mai_mai_n82_), .Y(mai_mai_n1357_));
  NA2        m1329(.A(mai_mai_n1205_), .B(mai_mai_n291_), .Y(mai_mai_n1358_));
  NA4        m1330(.A(mai_mai_n1358_), .B(mai_mai_n1357_), .C(mai_mai_n1355_), .D(mai_mai_n1352_), .Y(mai_mai_n1359_));
  NO2        m1331(.A(mai_mai_n1359_), .B(mai_mai_n1348_), .Y(mai_mai_n1360_));
  NO3        m1332(.A(e), .B(d), .C(c), .Y(mai_mai_n1361_));
  NA2        m1333(.A(mai_mai_n1522_), .B(mai_mai_n1361_), .Y(mai_mai_n1362_));
  NO2        m1334(.A(mai_mai_n1362_), .B(mai_mai_n215_), .Y(mai_mai_n1363_));
  OR2        m1335(.A(h), .B(f), .Y(mai_mai_n1364_));
  NO3        m1336(.A(n), .B(m), .C(i), .Y(mai_mai_n1365_));
  OAI210     m1337(.A0(mai_mai_n1114_), .A1(mai_mai_n155_), .B0(mai_mai_n1365_), .Y(mai_mai_n1366_));
  NO2        m1338(.A(mai_mai_n1366_), .B(mai_mai_n1364_), .Y(mai_mai_n1367_));
  NA3        m1339(.A(mai_mai_n699_), .B(mai_mai_n688_), .C(mai_mai_n113_), .Y(mai_mai_n1368_));
  NO2        m1340(.A(mai_mai_n1368_), .B(mai_mai_n45_), .Y(mai_mai_n1369_));
  NO2        m1341(.A(l), .B(k), .Y(mai_mai_n1370_));
  NOi41      m1342(.An(mai_mai_n550_), .B(mai_mai_n1370_), .C(mai_mai_n481_), .D(mai_mai_n446_), .Y(mai_mai_n1371_));
  NO3        m1343(.A(mai_mai_n446_), .B(d), .C(c), .Y(mai_mai_n1372_));
  NO4        m1344(.A(mai_mai_n1371_), .B(mai_mai_n1369_), .C(mai_mai_n1367_), .D(mai_mai_n1363_), .Y(mai_mai_n1373_));
  NO2        m1345(.A(mai_mai_n146_), .B(h), .Y(mai_mai_n1374_));
  NO2        m1346(.A(mai_mai_n1075_), .B(l), .Y(mai_mai_n1375_));
  NO2        m1347(.A(g), .B(c), .Y(mai_mai_n1376_));
  NA3        m1348(.A(mai_mai_n1376_), .B(mai_mai_n142_), .C(mai_mai_n186_), .Y(mai_mai_n1377_));
  NO2        m1349(.A(mai_mai_n1377_), .B(mai_mai_n1375_), .Y(mai_mai_n1378_));
  NA2        m1350(.A(mai_mai_n1378_), .B(mai_mai_n180_), .Y(mai_mai_n1379_));
  OAI210     m1351(.A0(mai_mai_n1350_), .A1(mai_mai_n214_), .B0(mai_mai_n1075_), .Y(mai_mai_n1380_));
  NO2        m1352(.A(mai_mai_n453_), .B(a), .Y(mai_mai_n1381_));
  NA3        m1353(.A(mai_mai_n1381_), .B(mai_mai_n1380_), .C(mai_mai_n114_), .Y(mai_mai_n1382_));
  NO2        m1354(.A(i), .B(h), .Y(mai_mai_n1383_));
  AOI210     m1355(.A0(mai_mai_n1138_), .A1(h), .B0(mai_mai_n420_), .Y(mai_mai_n1384_));
  NA2        m1356(.A(mai_mai_n139_), .B(mai_mai_n220_), .Y(mai_mai_n1385_));
  NO2        m1357(.A(mai_mai_n1385_), .B(mai_mai_n1384_), .Y(mai_mai_n1386_));
  NO2        m1358(.A(mai_mai_n756_), .B(mai_mai_n187_), .Y(mai_mai_n1387_));
  NOi31      m1359(.An(m), .B(n), .C(b), .Y(mai_mai_n1388_));
  NOi31      m1360(.An(f), .B(d), .C(c), .Y(mai_mai_n1389_));
  NA2        m1361(.A(mai_mai_n1389_), .B(mai_mai_n1388_), .Y(mai_mai_n1390_));
  INV        m1362(.A(mai_mai_n1390_), .Y(mai_mai_n1391_));
  NO3        m1363(.A(mai_mai_n1391_), .B(mai_mai_n1387_), .C(mai_mai_n1386_), .Y(mai_mai_n1392_));
  NA2        m1364(.A(mai_mai_n1086_), .B(mai_mai_n469_), .Y(mai_mai_n1393_));
  NO4        m1365(.A(mai_mai_n1393_), .B(mai_mai_n1060_), .C(mai_mai_n446_), .D(mai_mai_n45_), .Y(mai_mai_n1394_));
  OAI210     m1366(.A0(mai_mai_n183_), .A1(mai_mai_n529_), .B0(mai_mai_n1061_), .Y(mai_mai_n1395_));
  NO3        m1367(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1396_));
  INV        m1368(.A(mai_mai_n1395_), .Y(mai_mai_n1397_));
  NO2        m1369(.A(mai_mai_n1397_), .B(mai_mai_n1394_), .Y(mai_mai_n1398_));
  AN4        m1370(.A(mai_mai_n1398_), .B(mai_mai_n1392_), .C(mai_mai_n1382_), .D(mai_mai_n1379_), .Y(mai_mai_n1399_));
  NA2        m1371(.A(mai_mai_n1346_), .B(mai_mai_n383_), .Y(mai_mai_n1400_));
  NO2        m1372(.A(mai_mai_n1400_), .B(mai_mai_n1042_), .Y(mai_mai_n1401_));
  NA2        m1373(.A(mai_mai_n1372_), .B(mai_mai_n216_), .Y(mai_mai_n1402_));
  NO2        m1374(.A(mai_mai_n187_), .B(b), .Y(mai_mai_n1403_));
  AOI220     m1375(.A0(mai_mai_n1170_), .A1(mai_mai_n1403_), .B0(mai_mai_n1094_), .B1(mai_mai_n1393_), .Y(mai_mai_n1404_));
  NAi31      m1376(.An(mai_mai_n1401_), .B(mai_mai_n1404_), .C(mai_mai_n1402_), .Y(mai_mai_n1405_));
  NO4        m1377(.A(mai_mai_n133_), .B(g), .C(f), .D(e), .Y(mai_mai_n1406_));
  NA3        m1378(.A(mai_mai_n1351_), .B(mai_mai_n292_), .C(h), .Y(mai_mai_n1407_));
  OR2        m1379(.A(e), .B(a), .Y(mai_mai_n1408_));
  NO2        m1380(.A(mai_mai_n1343_), .B(mai_mai_n1342_), .Y(mai_mai_n1409_));
  AOI210     m1381(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1409_), .Y(mai_mai_n1410_));
  NO2        m1382(.A(mai_mai_n1410_), .B(mai_mai_n1082_), .Y(mai_mai_n1411_));
  NA2        m1383(.A(mai_mai_n1349_), .B(mai_mai_n1370_), .Y(mai_mai_n1412_));
  INV        m1384(.A(mai_mai_n1412_), .Y(mai_mai_n1413_));
  OR3        m1385(.A(mai_mai_n544_), .B(mai_mai_n543_), .C(mai_mai_n113_), .Y(mai_mai_n1414_));
  NA2        m1386(.A(mai_mai_n1112_), .B(mai_mai_n412_), .Y(mai_mai_n1415_));
  NO2        m1387(.A(mai_mai_n1415_), .B(mai_mai_n441_), .Y(mai_mai_n1416_));
  AO210      m1388(.A0(mai_mai_n1416_), .A1(mai_mai_n117_), .B0(mai_mai_n1413_), .Y(mai_mai_n1417_));
  NO3        m1389(.A(mai_mai_n1417_), .B(mai_mai_n1411_), .C(mai_mai_n1405_), .Y(mai_mai_n1418_));
  NA4        m1390(.A(mai_mai_n1418_), .B(mai_mai_n1399_), .C(mai_mai_n1373_), .D(mai_mai_n1360_), .Y(mai_mai_n1419_));
  NO2        m1391(.A(mai_mai_n395_), .B(j), .Y(mai_mai_n1420_));
  NA3        m1392(.A(mai_mai_n1396_), .B(mai_mai_n1343_), .C(mai_mai_n1112_), .Y(mai_mai_n1421_));
  NAi41      m1393(.An(mai_mai_n1383_), .B(mai_mai_n1073_), .C(mai_mai_n168_), .D(mai_mai_n149_), .Y(mai_mai_n1422_));
  NA2        m1394(.A(mai_mai_n1422_), .B(mai_mai_n1421_), .Y(mai_mai_n1423_));
  NA3        m1395(.A(g), .B(mai_mai_n1420_), .C(mai_mai_n157_), .Y(mai_mai_n1424_));
  INV        m1396(.A(mai_mai_n1424_), .Y(mai_mai_n1425_));
  NO3        m1397(.A(mai_mai_n749_), .B(mai_mai_n175_), .C(mai_mai_n415_), .Y(mai_mai_n1426_));
  NO3        m1398(.A(mai_mai_n1426_), .B(mai_mai_n1425_), .C(mai_mai_n1423_), .Y(mai_mai_n1427_));
  OR2        m1399(.A(n), .B(i), .Y(mai_mai_n1428_));
  OAI210     m1400(.A0(mai_mai_n1428_), .A1(mai_mai_n1072_), .B0(mai_mai_n49_), .Y(mai_mai_n1429_));
  AOI220     m1401(.A0(mai_mai_n1429_), .A1(mai_mai_n1176_), .B0(mai_mai_n827_), .B1(mai_mai_n194_), .Y(mai_mai_n1430_));
  INV        m1402(.A(mai_mai_n1430_), .Y(mai_mai_n1431_));
  NO2        m1403(.A(mai_mai_n133_), .B(l), .Y(mai_mai_n1432_));
  NO2        m1404(.A(mai_mai_n224_), .B(k), .Y(mai_mai_n1433_));
  OAI210     m1405(.A0(mai_mai_n1433_), .A1(mai_mai_n1383_), .B0(mai_mai_n1432_), .Y(mai_mai_n1434_));
  NO2        m1406(.A(mai_mai_n1434_), .B(mai_mai_n31_), .Y(mai_mai_n1435_));
  NO3        m1407(.A(mai_mai_n1414_), .B(mai_mai_n469_), .C(mai_mai_n354_), .Y(mai_mai_n1436_));
  NO3        m1408(.A(mai_mai_n1436_), .B(mai_mai_n1435_), .C(mai_mai_n1431_), .Y(mai_mai_n1437_));
  NO3        m1409(.A(mai_mai_n1097_), .B(mai_mai_n1343_), .C(mai_mai_n49_), .Y(mai_mai_n1438_));
  NO2        m1410(.A(mai_mai_n1082_), .B(h), .Y(mai_mai_n1439_));
  NA3        m1411(.A(mai_mai_n1439_), .B(d), .C(mai_mai_n1043_), .Y(mai_mai_n1440_));
  NO2        m1412(.A(mai_mai_n1440_), .B(c), .Y(mai_mai_n1441_));
  NA2        m1413(.A(mai_mai_n180_), .B(mai_mai_n113_), .Y(mai_mai_n1442_));
  NOi21      m1414(.An(d), .B(f), .Y(mai_mai_n1443_));
  NO2        m1415(.A(mai_mai_n1343_), .B(f), .Y(mai_mai_n1444_));
  INV        m1416(.A(mai_mai_n1441_), .Y(mai_mai_n1445_));
  NA3        m1417(.A(mai_mai_n1445_), .B(mai_mai_n1437_), .C(mai_mai_n1427_), .Y(mai_mai_n1446_));
  NO3        m1418(.A(mai_mai_n1086_), .B(mai_mai_n1072_), .C(mai_mai_n40_), .Y(mai_mai_n1447_));
  NO2        m1419(.A(mai_mai_n469_), .B(mai_mai_n301_), .Y(mai_mai_n1448_));
  OAI210     m1420(.A0(mai_mai_n1448_), .A1(mai_mai_n1447_), .B0(mai_mai_n1356_), .Y(mai_mai_n1449_));
  OAI210     m1421(.A0(mai_mai_n1406_), .A1(mai_mai_n1346_), .B0(mai_mai_n887_), .Y(mai_mai_n1450_));
  OAI220     m1422(.A0(mai_mai_n1039_), .A1(mai_mai_n133_), .B0(mai_mai_n669_), .B1(mai_mai_n175_), .Y(mai_mai_n1451_));
  NA2        m1423(.A(mai_mai_n1451_), .B(mai_mai_n624_), .Y(mai_mai_n1452_));
  NA3        m1424(.A(mai_mai_n1452_), .B(mai_mai_n1450_), .C(mai_mai_n1449_), .Y(mai_mai_n1453_));
  NA2        m1425(.A(mai_mai_n1376_), .B(mai_mai_n1443_), .Y(mai_mai_n1454_));
  NO2        m1426(.A(mai_mai_n1454_), .B(m), .Y(mai_mai_n1455_));
  NO2        m1427(.A(mai_mai_n150_), .B(mai_mai_n182_), .Y(mai_mai_n1456_));
  OAI210     m1428(.A0(mai_mai_n1456_), .A1(mai_mai_n111_), .B0(mai_mai_n1388_), .Y(mai_mai_n1457_));
  INV        m1429(.A(mai_mai_n1457_), .Y(mai_mai_n1458_));
  NO3        m1430(.A(mai_mai_n1458_), .B(mai_mai_n1455_), .C(mai_mai_n1453_), .Y(mai_mai_n1459_));
  NO2        m1431(.A(mai_mai_n1342_), .B(e), .Y(mai_mai_n1460_));
  NA2        m1432(.A(mai_mai_n1460_), .B(mai_mai_n410_), .Y(mai_mai_n1461_));
  OAI210     m1433(.A0(mai_mai_n1444_), .A1(mai_mai_n1123_), .B0(mai_mai_n633_), .Y(mai_mai_n1462_));
  OR3        m1434(.A(mai_mai_n1433_), .B(mai_mai_n1205_), .C(mai_mai_n133_), .Y(mai_mai_n1463_));
  OAI220     m1435(.A0(mai_mai_n1463_), .A1(mai_mai_n1461_), .B0(mai_mai_n1462_), .B1(mai_mai_n448_), .Y(mai_mai_n1464_));
  INV        m1436(.A(mai_mai_n1464_), .Y(mai_mai_n1465_));
  NO2        m1437(.A(mai_mai_n182_), .B(c), .Y(mai_mai_n1466_));
  OAI210     m1438(.A0(mai_mai_n1466_), .A1(mai_mai_n1460_), .B0(mai_mai_n180_), .Y(mai_mai_n1467_));
  AOI220     m1439(.A0(mai_mai_n1467_), .A1(mai_mai_n1074_), .B0(mai_mai_n535_), .B1(mai_mai_n370_), .Y(mai_mai_n1468_));
  NA2        m1440(.A(mai_mai_n543_), .B(g), .Y(mai_mai_n1469_));
  AOI210     m1441(.A0(mai_mai_n1469_), .A1(mai_mai_n1372_), .B0(mai_mai_n1438_), .Y(mai_mai_n1470_));
  NO2        m1442(.A(mai_mai_n1408_), .B(f), .Y(mai_mai_n1471_));
  NA2        m1443(.A(mai_mai_n1123_), .B(a), .Y(mai_mai_n1472_));
  OAI220     m1444(.A0(mai_mai_n1472_), .A1(mai_mai_n69_), .B0(mai_mai_n1470_), .B1(mai_mai_n214_), .Y(mai_mai_n1473_));
  AOI210     m1445(.A0(mai_mai_n903_), .A1(mai_mai_n422_), .B0(mai_mai_n105_), .Y(mai_mai_n1474_));
  OR2        m1446(.A(mai_mai_n1474_), .B(mai_mai_n543_), .Y(mai_mai_n1475_));
  NA2        m1447(.A(mai_mai_n1471_), .B(mai_mai_n1353_), .Y(mai_mai_n1476_));
  OAI220     m1448(.A0(mai_mai_n1476_), .A1(mai_mai_n49_), .B0(mai_mai_n1475_), .B1(mai_mai_n175_), .Y(mai_mai_n1477_));
  NA4        m1449(.A(mai_mai_n1095_), .B(mai_mai_n1092_), .C(mai_mai_n220_), .D(mai_mai_n68_), .Y(mai_mai_n1478_));
  NA2        m1450(.A(mai_mai_n1347_), .B(mai_mai_n183_), .Y(mai_mai_n1479_));
  NO2        m1451(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1480_));
  OAI210     m1452(.A0(mai_mai_n1408_), .A1(mai_mai_n864_), .B0(mai_mai_n486_), .Y(mai_mai_n1481_));
  OAI210     m1453(.A0(mai_mai_n1481_), .A1(mai_mai_n1098_), .B0(mai_mai_n1480_), .Y(mai_mai_n1482_));
  NO2        m1454(.A(mai_mai_n252_), .B(g), .Y(mai_mai_n1483_));
  NO2        m1455(.A(m), .B(i), .Y(mai_mai_n1484_));
  BUFFER     m1456(.A(mai_mai_n1484_), .Y(mai_mai_n1485_));
  AOI220     m1457(.A0(mai_mai_n1485_), .A1(mai_mai_n1374_), .B0(mai_mai_n1073_), .B1(mai_mai_n1483_), .Y(mai_mai_n1486_));
  NA4        m1458(.A(mai_mai_n1486_), .B(mai_mai_n1482_), .C(mai_mai_n1479_), .D(mai_mai_n1478_), .Y(mai_mai_n1487_));
  NO4        m1459(.A(mai_mai_n1487_), .B(mai_mai_n1477_), .C(mai_mai_n1473_), .D(mai_mai_n1468_), .Y(mai_mai_n1488_));
  NA3        m1460(.A(mai_mai_n1488_), .B(mai_mai_n1465_), .C(mai_mai_n1459_), .Y(mai_mai_n1489_));
  NA3        m1461(.A(mai_mai_n962_), .B(mai_mai_n139_), .C(mai_mai_n46_), .Y(mai_mai_n1490_));
  AOI210     m1462(.A0(mai_mai_n147_), .A1(c), .B0(mai_mai_n1490_), .Y(mai_mai_n1491_));
  INV        m1463(.A(mai_mai_n184_), .Y(mai_mai_n1492_));
  NA2        m1464(.A(mai_mai_n1492_), .B(mai_mai_n1439_), .Y(mai_mai_n1493_));
  AO210      m1465(.A0(mai_mai_n134_), .A1(l), .B0(mai_mai_n1400_), .Y(mai_mai_n1494_));
  NA2        m1466(.A(mai_mai_n1494_), .B(mai_mai_n1493_), .Y(mai_mai_n1495_));
  NO2        m1467(.A(mai_mai_n1495_), .B(mai_mai_n1491_), .Y(mai_mai_n1496_));
  AOI210     m1468(.A0(mai_mai_n155_), .A1(mai_mai_n56_), .B0(mai_mai_n1460_), .Y(mai_mai_n1497_));
  NO2        m1469(.A(mai_mai_n1497_), .B(mai_mai_n1442_), .Y(mai_mai_n1498_));
  NOi21      m1470(.An(mai_mai_n1347_), .B(e), .Y(mai_mai_n1499_));
  NO2        m1471(.A(mai_mai_n1499_), .B(mai_mai_n1498_), .Y(mai_mai_n1500_));
  AN2        m1472(.A(mai_mai_n1095_), .B(mai_mai_n1080_), .Y(mai_mai_n1501_));
  AOI220     m1473(.A0(mai_mai_n1484_), .A1(mai_mai_n642_), .B0(mai_mai_n1057_), .B1(mai_mai_n158_), .Y(mai_mai_n1502_));
  NOi31      m1474(.An(mai_mai_n30_), .B(mai_mai_n1502_), .C(n), .Y(mai_mai_n1503_));
  AOI210     m1475(.A0(mai_mai_n1501_), .A1(mai_mai_n1170_), .B0(mai_mai_n1503_), .Y(mai_mai_n1504_));
  NA2        m1476(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1505_));
  NO2        m1477(.A(mai_mai_n1351_), .B(mai_mai_n119_), .Y(mai_mai_n1506_));
  OAI220     m1478(.A0(mai_mai_n1506_), .A1(mai_mai_n1400_), .B0(mai_mai_n1415_), .B1(mai_mai_n1505_), .Y(mai_mai_n1507_));
  INV        m1479(.A(mai_mai_n1507_), .Y(mai_mai_n1508_));
  NA4        m1480(.A(mai_mai_n1508_), .B(mai_mai_n1504_), .C(mai_mai_n1500_), .D(mai_mai_n1496_), .Y(mai_mai_n1509_));
  OR4        m1481(.A(mai_mai_n1509_), .B(mai_mai_n1489_), .C(mai_mai_n1446_), .D(mai_mai_n1419_), .Y(mai04));
  NOi31      m1482(.An(mai_mai_n1406_), .B(mai_mai_n1407_), .C(mai_mai_n1045_), .Y(mai_mai_n1511_));
  NA2        m1483(.A(mai_mai_n1444_), .B(mai_mai_n827_), .Y(mai_mai_n1512_));
  NO4        m1484(.A(mai_mai_n1512_), .B(mai_mai_n1034_), .C(mai_mai_n487_), .D(j), .Y(mai_mai_n1513_));
  OR3        m1485(.A(mai_mai_n1513_), .B(mai_mai_n1511_), .C(mai_mai_n1063_), .Y(mai_mai_n1514_));
  NO3        m1486(.A(mai_mai_n1353_), .B(mai_mai_n92_), .C(k), .Y(mai_mai_n1515_));
  AOI210     m1487(.A0(mai_mai_n1515_), .A1(mai_mai_n1056_), .B0(mai_mai_n1185_), .Y(mai_mai_n1516_));
  NA2        m1488(.A(mai_mai_n1516_), .B(mai_mai_n1209_), .Y(mai_mai_n1517_));
  NO4        m1489(.A(mai_mai_n1517_), .B(mai_mai_n1514_), .C(mai_mai_n1071_), .D(mai_mai_n1050_), .Y(mai_mai_n1518_));
  NA4        m1490(.A(mai_mai_n1518_), .B(mai_mai_n1125_), .C(mai_mai_n1110_), .D(mai_mai_n1101_), .Y(mai05));
  INV        m1491(.A(m), .Y(mai_mai_n1522_));
  INV        m1492(.A(mai_mai_n950_), .Y(mai_mai_n1523_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(g), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(g), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(g), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(g), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n74_), .B(men_men_n64_), .Y(men_men_n83_));
  INV        u0055(.A(n), .Y(men_men_n84_));
  NOi32      u0056(.An(e), .Bn(b), .C(d), .Y(men_men_n85_));
  NA2        u0057(.A(men_men_n85_), .B(men_men_n84_), .Y(men_men_n86_));
  INV        u0058(.A(j), .Y(men_men_n87_));
  AN3        u0059(.A(m), .B(k), .C(i), .Y(men_men_n88_));
  NA3        u0060(.A(men_men_n88_), .B(men_men_n87_), .C(g), .Y(men_men_n89_));
  NO2        u0061(.A(men_men_n89_), .B(f), .Y(men_men_n90_));
  NAi32      u0062(.An(g), .Bn(f), .C(h), .Y(men_men_n91_));
  NAi31      u0063(.An(j), .B(m), .C(l), .Y(men_men_n92_));
  NO2        u0064(.A(men_men_n92_), .B(men_men_n91_), .Y(men_men_n93_));
  NA2        u0065(.A(m), .B(l), .Y(men_men_n94_));
  NAi31      u0066(.An(k), .B(j), .C(g), .Y(men_men_n95_));
  NO3        u0067(.A(men_men_n95_), .B(men_men_n94_), .C(f), .Y(men_men_n96_));
  AN2        u0068(.A(j), .B(g), .Y(men_men_n97_));
  NOi32      u0069(.An(m), .Bn(l), .C(i), .Y(men_men_n98_));
  NOi21      u0070(.An(g), .B(i), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(j), .C(k), .Y(men_men_n100_));
  AOI220     u0072(.A0(men_men_n100_), .A1(men_men_n99_), .B0(men_men_n98_), .B1(men_men_n97_), .Y(men_men_n101_));
  NO2        u0073(.A(men_men_n101_), .B(f), .Y(men_men_n102_));
  NO4        u0074(.A(men_men_n102_), .B(men_men_n96_), .C(men_men_n93_), .D(men_men_n90_), .Y(men_men_n103_));
  NAi41      u0075(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n104_));
  AN2        u0076(.A(e), .B(b), .Y(men_men_n105_));
  NOi31      u0077(.An(c), .B(h), .C(f), .Y(men_men_n106_));
  NA2        u0078(.A(men_men_n106_), .B(men_men_n105_), .Y(men_men_n107_));
  NOi21      u0079(.An(g), .B(f), .Y(men_men_n108_));
  NOi21      u0080(.An(i), .B(h), .Y(men_men_n109_));
  NA3        u0081(.A(men_men_n109_), .B(men_men_n108_), .C(men_men_n36_), .Y(men_men_n110_));
  INV        u0082(.A(a), .Y(men_men_n111_));
  NA2        u0083(.A(men_men_n105_), .B(men_men_n111_), .Y(men_men_n112_));
  INV        u0084(.A(l), .Y(men_men_n113_));
  NOi21      u0085(.An(m), .B(n), .Y(men_men_n114_));
  AN2        u0086(.A(k), .B(h), .Y(men_men_n115_));
  NO2        u0087(.A(men_men_n110_), .B(men_men_n86_), .Y(men_men_n116_));
  INV        u0088(.A(b), .Y(men_men_n117_));
  NA2        u0089(.A(l), .B(j), .Y(men_men_n118_));
  AN2        u0090(.A(k), .B(i), .Y(men_men_n119_));
  NA2        u0091(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NA2        u0092(.A(g), .B(e), .Y(men_men_n121_));
  NOi32      u0093(.An(c), .Bn(a), .C(d), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n114_), .Y(men_men_n123_));
  NO4        u0095(.A(men_men_n123_), .B(men_men_n121_), .C(men_men_n120_), .D(men_men_n117_), .Y(men_men_n124_));
  NO2        u0096(.A(men_men_n124_), .B(men_men_n116_), .Y(men_men_n125_));
  OAI210     u0097(.A0(men_men_n103_), .A1(men_men_n86_), .B0(men_men_n125_), .Y(men_men_n126_));
  NOi31      u0098(.An(k), .B(m), .C(j), .Y(men_men_n127_));
  NA3        u0099(.A(men_men_n127_), .B(men_men_n79_), .C(men_men_n78_), .Y(men_men_n128_));
  NOi31      u0100(.An(k), .B(m), .C(i), .Y(men_men_n129_));
  NA3        u0101(.A(men_men_n129_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n130_));
  NA2        u0102(.A(men_men_n130_), .B(men_men_n128_), .Y(men_men_n131_));
  NOi32      u0103(.An(f), .Bn(b), .C(e), .Y(men_men_n132_));
  NAi21      u0104(.An(g), .B(h), .Y(men_men_n133_));
  NAi21      u0105(.An(m), .B(n), .Y(men_men_n134_));
  NAi21      u0106(.An(j), .B(k), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n133_), .Y(men_men_n136_));
  NAi41      u0108(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n137_));
  NAi31      u0109(.An(j), .B(k), .C(h), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n134_), .Y(men_men_n139_));
  AOI210     u0111(.A0(men_men_n136_), .A1(men_men_n132_), .B0(men_men_n139_), .Y(men_men_n140_));
  NO2        u0112(.A(k), .B(j), .Y(men_men_n141_));
  NO2        u0113(.A(men_men_n141_), .B(men_men_n134_), .Y(men_men_n142_));
  AN2        u0114(.A(k), .B(j), .Y(men_men_n143_));
  NAi21      u0115(.An(c), .B(b), .Y(men_men_n144_));
  NA2        u0116(.A(f), .B(d), .Y(men_men_n145_));
  NO4        u0117(.A(men_men_n145_), .B(men_men_n144_), .C(men_men_n143_), .D(men_men_n133_), .Y(men_men_n146_));
  NA2        u0118(.A(h), .B(c), .Y(men_men_n147_));
  NAi31      u0119(.An(f), .B(e), .C(b), .Y(men_men_n148_));
  NA2        u0120(.A(men_men_n146_), .B(men_men_n142_), .Y(men_men_n149_));
  NA2        u0121(.A(d), .B(b), .Y(men_men_n150_));
  NAi21      u0122(.An(e), .B(f), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n151_), .B(men_men_n150_), .Y(men_men_n152_));
  NA2        u0124(.A(b), .B(a), .Y(men_men_n153_));
  NAi21      u0125(.An(e), .B(g), .Y(men_men_n154_));
  NAi21      u0126(.An(c), .B(d), .Y(men_men_n155_));
  NAi31      u0127(.An(l), .B(k), .C(h), .Y(men_men_n156_));
  NO2        u0128(.A(men_men_n134_), .B(men_men_n156_), .Y(men_men_n157_));
  NA2        u0129(.A(men_men_n157_), .B(men_men_n152_), .Y(men_men_n158_));
  NAi41      u0130(.An(men_men_n131_), .B(men_men_n158_), .C(men_men_n149_), .D(men_men_n140_), .Y(men_men_n159_));
  NAi31      u0131(.An(e), .B(f), .C(b), .Y(men_men_n160_));
  NOi21      u0132(.An(g), .B(d), .Y(men_men_n161_));
  NO2        u0133(.A(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  NOi21      u0134(.An(h), .B(i), .Y(men_men_n163_));
  NOi21      u0135(.An(k), .B(m), .Y(men_men_n164_));
  NA3        u0136(.A(men_men_n164_), .B(men_men_n163_), .C(n), .Y(men_men_n165_));
  NOi21      u0137(.An(h), .B(g), .Y(men_men_n166_));
  NO2        u0138(.A(men_men_n145_), .B(men_men_n144_), .Y(men_men_n167_));
  NA2        u0139(.A(men_men_n167_), .B(men_men_n166_), .Y(men_men_n168_));
  NAi31      u0140(.An(l), .B(j), .C(h), .Y(men_men_n169_));
  NO2        u0141(.A(men_men_n169_), .B(men_men_n49_), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n67_), .Y(men_men_n171_));
  NOi32      u0143(.An(n), .Bn(k), .C(m), .Y(men_men_n172_));
  NA2        u0144(.A(l), .B(i), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  OAI210     u0146(.A0(men_men_n174_), .A1(men_men_n168_), .B0(men_men_n171_), .Y(men_men_n175_));
  NAi31      u0147(.An(d), .B(f), .C(c), .Y(men_men_n176_));
  NAi31      u0148(.An(e), .B(f), .C(c), .Y(men_men_n177_));
  NA2        u0149(.A(men_men_n177_), .B(men_men_n176_), .Y(men_men_n178_));
  NA2        u0150(.A(j), .B(h), .Y(men_men_n179_));
  OR3        u0151(.A(n), .B(m), .C(k), .Y(men_men_n180_));
  NO2        u0152(.A(men_men_n180_), .B(men_men_n179_), .Y(men_men_n181_));
  NAi32      u0153(.An(m), .Bn(k), .C(n), .Y(men_men_n182_));
  NO2        u0154(.A(men_men_n182_), .B(men_men_n179_), .Y(men_men_n183_));
  AOI220     u0155(.A0(men_men_n183_), .A1(men_men_n162_), .B0(men_men_n181_), .B1(men_men_n178_), .Y(men_men_n184_));
  NO2        u0156(.A(n), .B(m), .Y(men_men_n185_));
  NA2        u0157(.A(men_men_n185_), .B(men_men_n50_), .Y(men_men_n186_));
  NAi21      u0158(.An(f), .B(e), .Y(men_men_n187_));
  NA2        u0159(.A(d), .B(c), .Y(men_men_n188_));
  NO2        u0160(.A(men_men_n188_), .B(men_men_n187_), .Y(men_men_n189_));
  NOi21      u0161(.An(men_men_n189_), .B(men_men_n186_), .Y(men_men_n190_));
  NAi21      u0162(.An(d), .B(c), .Y(men_men_n191_));
  NAi31      u0163(.An(m), .B(n), .C(b), .Y(men_men_n192_));
  NA2        u0164(.A(k), .B(i), .Y(men_men_n193_));
  NAi21      u0165(.An(h), .B(f), .Y(men_men_n194_));
  NO2        u0166(.A(men_men_n194_), .B(men_men_n193_), .Y(men_men_n195_));
  NO2        u0167(.A(men_men_n192_), .B(men_men_n155_), .Y(men_men_n196_));
  NA2        u0168(.A(men_men_n196_), .B(men_men_n195_), .Y(men_men_n197_));
  NOi32      u0169(.An(f), .Bn(c), .C(d), .Y(men_men_n198_));
  NOi32      u0170(.An(f), .Bn(c), .C(e), .Y(men_men_n199_));
  NO2        u0171(.A(men_men_n199_), .B(men_men_n198_), .Y(men_men_n200_));
  NO3        u0172(.A(n), .B(m), .C(j), .Y(men_men_n201_));
  NA2        u0173(.A(men_men_n201_), .B(men_men_n115_), .Y(men_men_n202_));
  AO210      u0174(.A0(men_men_n202_), .A1(men_men_n186_), .B0(men_men_n200_), .Y(men_men_n203_));
  NAi41      u0175(.An(men_men_n190_), .B(men_men_n203_), .C(men_men_n197_), .D(men_men_n184_), .Y(men_men_n204_));
  OR3        u0176(.A(men_men_n204_), .B(men_men_n175_), .C(men_men_n159_), .Y(men_men_n205_));
  NO4        u0177(.A(men_men_n205_), .B(men_men_n126_), .C(men_men_n83_), .D(men_men_n55_), .Y(men_men_n206_));
  NA3        u0178(.A(m), .B(men_men_n113_), .C(j), .Y(men_men_n207_));
  NAi31      u0179(.An(n), .B(h), .C(g), .Y(men_men_n208_));
  NO2        u0180(.A(men_men_n208_), .B(men_men_n207_), .Y(men_men_n209_));
  NOi32      u0181(.An(m), .Bn(k), .C(l), .Y(men_men_n210_));
  NA3        u0182(.A(men_men_n210_), .B(men_men_n87_), .C(g), .Y(men_men_n211_));
  NO2        u0183(.A(men_men_n211_), .B(n), .Y(men_men_n212_));
  NOi21      u0184(.An(k), .B(j), .Y(men_men_n213_));
  NA4        u0185(.A(men_men_n213_), .B(men_men_n114_), .C(i), .D(g), .Y(men_men_n214_));
  AN2        u0186(.A(i), .B(g), .Y(men_men_n215_));
  NA3        u0187(.A(men_men_n76_), .B(men_men_n215_), .C(men_men_n114_), .Y(men_men_n216_));
  NA2        u0188(.A(men_men_n216_), .B(men_men_n214_), .Y(men_men_n217_));
  NO3        u0189(.A(men_men_n217_), .B(men_men_n212_), .C(men_men_n209_), .Y(men_men_n218_));
  NAi41      u0190(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n219_));
  INV        u0191(.A(men_men_n219_), .Y(men_men_n220_));
  INV        u0192(.A(f), .Y(men_men_n221_));
  INV        u0193(.A(g), .Y(men_men_n222_));
  NOi31      u0194(.An(i), .B(j), .C(h), .Y(men_men_n223_));
  NOi21      u0195(.An(l), .B(m), .Y(men_men_n224_));
  NA2        u0196(.A(men_men_n224_), .B(men_men_n223_), .Y(men_men_n225_));
  NO3        u0197(.A(men_men_n225_), .B(men_men_n222_), .C(men_men_n221_), .Y(men_men_n226_));
  NA2        u0198(.A(men_men_n226_), .B(men_men_n220_), .Y(men_men_n227_));
  OAI210     u0199(.A0(men_men_n218_), .A1(men_men_n32_), .B0(men_men_n227_), .Y(men_men_n228_));
  NOi21      u0200(.An(n), .B(m), .Y(men_men_n229_));
  NOi32      u0201(.An(l), .Bn(i), .C(j), .Y(men_men_n230_));
  NA2        u0202(.A(men_men_n230_), .B(men_men_n229_), .Y(men_men_n231_));
  OA220      u0203(.A0(men_men_n231_), .A1(men_men_n107_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n232_));
  NAi21      u0204(.An(j), .B(h), .Y(men_men_n233_));
  XN2        u0205(.A(i), .B(h), .Y(men_men_n234_));
  NA2        u0206(.A(men_men_n234_), .B(men_men_n233_), .Y(men_men_n235_));
  NOi31      u0207(.An(k), .B(n), .C(m), .Y(men_men_n236_));
  NOi31      u0208(.An(men_men_n236_), .B(men_men_n188_), .C(men_men_n187_), .Y(men_men_n237_));
  NA2        u0209(.A(men_men_n237_), .B(men_men_n235_), .Y(men_men_n238_));
  NAi31      u0210(.An(f), .B(e), .C(c), .Y(men_men_n239_));
  NO4        u0211(.A(men_men_n239_), .B(men_men_n180_), .C(men_men_n179_), .D(men_men_n59_), .Y(men_men_n240_));
  NA4        u0212(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n241_));
  NAi32      u0213(.An(m), .Bn(i), .C(k), .Y(men_men_n242_));
  NO3        u0214(.A(men_men_n242_), .B(men_men_n91_), .C(men_men_n241_), .Y(men_men_n243_));
  NA2        u0215(.A(k), .B(h), .Y(men_men_n244_));
  NO2        u0216(.A(men_men_n243_), .B(men_men_n240_), .Y(men_men_n245_));
  NAi21      u0217(.An(n), .B(a), .Y(men_men_n246_));
  NO2        u0218(.A(men_men_n246_), .B(men_men_n150_), .Y(men_men_n247_));
  NAi41      u0219(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n248_));
  NO2        u0220(.A(men_men_n248_), .B(e), .Y(men_men_n249_));
  NO3        u0221(.A(men_men_n151_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n250_));
  OAI210     u0222(.A0(men_men_n250_), .A1(men_men_n249_), .B0(men_men_n247_), .Y(men_men_n251_));
  AN4        u0223(.A(men_men_n251_), .B(men_men_n245_), .C(men_men_n238_), .D(men_men_n232_), .Y(men_men_n252_));
  OR2        u0224(.A(h), .B(g), .Y(men_men_n253_));
  NO2        u0225(.A(men_men_n253_), .B(men_men_n104_), .Y(men_men_n254_));
  NA2        u0226(.A(men_men_n254_), .B(men_men_n132_), .Y(men_men_n255_));
  NAi41      u0227(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n256_));
  NO2        u0228(.A(men_men_n256_), .B(men_men_n221_), .Y(men_men_n257_));
  NA2        u0229(.A(men_men_n164_), .B(men_men_n109_), .Y(men_men_n258_));
  NAi21      u0230(.An(men_men_n258_), .B(men_men_n257_), .Y(men_men_n259_));
  NO2        u0231(.A(n), .B(a), .Y(men_men_n260_));
  NAi31      u0232(.An(men_men_n248_), .B(men_men_n260_), .C(men_men_n105_), .Y(men_men_n261_));
  AN2        u0233(.A(men_men_n261_), .B(men_men_n259_), .Y(men_men_n262_));
  NAi21      u0234(.An(h), .B(i), .Y(men_men_n263_));
  NA2        u0235(.A(men_men_n185_), .B(k), .Y(men_men_n264_));
  NO2        u0236(.A(men_men_n264_), .B(men_men_n263_), .Y(men_men_n265_));
  NA2        u0237(.A(men_men_n265_), .B(men_men_n198_), .Y(men_men_n266_));
  NA3        u0238(.A(men_men_n266_), .B(men_men_n262_), .C(men_men_n255_), .Y(men_men_n267_));
  NOi21      u0239(.An(g), .B(e), .Y(men_men_n268_));
  NO2        u0240(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n269_));
  NA2        u0241(.A(men_men_n269_), .B(men_men_n268_), .Y(men_men_n270_));
  NOi32      u0242(.An(l), .Bn(j), .C(i), .Y(men_men_n271_));
  AOI210     u0243(.A0(men_men_n76_), .A1(men_men_n87_), .B0(men_men_n271_), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n263_), .B(men_men_n44_), .Y(men_men_n273_));
  NAi21      u0245(.An(f), .B(g), .Y(men_men_n274_));
  NO2        u0246(.A(men_men_n274_), .B(men_men_n65_), .Y(men_men_n275_));
  NO2        u0247(.A(men_men_n69_), .B(men_men_n118_), .Y(men_men_n276_));
  AOI220     u0248(.A0(men_men_n276_), .A1(men_men_n275_), .B0(men_men_n273_), .B1(men_men_n67_), .Y(men_men_n277_));
  OAI210     u0249(.A0(men_men_n272_), .A1(men_men_n270_), .B0(men_men_n277_), .Y(men_men_n278_));
  NO3        u0250(.A(men_men_n135_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n279_));
  NOi41      u0251(.An(men_men_n252_), .B(men_men_n278_), .C(men_men_n267_), .D(men_men_n228_), .Y(men_men_n280_));
  NO4        u0252(.A(men_men_n209_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n281_));
  NO2        u0253(.A(men_men_n281_), .B(men_men_n112_), .Y(men_men_n282_));
  NA3        u0254(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n283_));
  NAi21      u0255(.An(h), .B(g), .Y(men_men_n284_));
  OR4        u0256(.A(men_men_n284_), .B(men_men_n283_), .C(men_men_n231_), .D(e), .Y(men_men_n285_));
  NO2        u0257(.A(men_men_n258_), .B(men_men_n274_), .Y(men_men_n286_));
  NA2        u0258(.A(men_men_n286_), .B(men_men_n78_), .Y(men_men_n287_));
  NAi31      u0259(.An(g), .B(k), .C(h), .Y(men_men_n288_));
  NO3        u0260(.A(men_men_n134_), .B(men_men_n288_), .C(l), .Y(men_men_n289_));
  NAi31      u0261(.An(e), .B(d), .C(a), .Y(men_men_n290_));
  NA2        u0262(.A(men_men_n289_), .B(men_men_n132_), .Y(men_men_n291_));
  NA3        u0263(.A(men_men_n291_), .B(men_men_n287_), .C(men_men_n285_), .Y(men_men_n292_));
  NA4        u0264(.A(men_men_n164_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n118_), .Y(men_men_n293_));
  NA3        u0265(.A(men_men_n164_), .B(men_men_n163_), .C(men_men_n84_), .Y(men_men_n294_));
  NO2        u0266(.A(men_men_n294_), .B(men_men_n200_), .Y(men_men_n295_));
  NOi21      u0267(.An(men_men_n293_), .B(men_men_n295_), .Y(men_men_n296_));
  NA3        u0268(.A(e), .B(c), .C(b), .Y(men_men_n297_));
  NO2        u0269(.A(men_men_n60_), .B(men_men_n297_), .Y(men_men_n298_));
  NAi32      u0270(.An(k), .Bn(i), .C(j), .Y(men_men_n299_));
  NAi31      u0271(.An(h), .B(l), .C(i), .Y(men_men_n300_));
  NA3        u0272(.A(men_men_n300_), .B(men_men_n299_), .C(men_men_n169_), .Y(men_men_n301_));
  NOi21      u0273(.An(men_men_n301_), .B(men_men_n49_), .Y(men_men_n302_));
  OAI210     u0274(.A0(men_men_n275_), .A1(men_men_n298_), .B0(men_men_n302_), .Y(men_men_n303_));
  NAi21      u0275(.An(l), .B(k), .Y(men_men_n304_));
  NO2        u0276(.A(men_men_n304_), .B(men_men_n49_), .Y(men_men_n305_));
  NOi21      u0277(.An(l), .B(j), .Y(men_men_n306_));
  NA2        u0278(.A(men_men_n166_), .B(men_men_n306_), .Y(men_men_n307_));
  NA3        u0279(.A(men_men_n119_), .B(men_men_n118_), .C(g), .Y(men_men_n308_));
  OR3        u0280(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n309_));
  AOI210     u0281(.A0(men_men_n308_), .A1(men_men_n307_), .B0(men_men_n309_), .Y(men_men_n310_));
  INV        u0282(.A(men_men_n310_), .Y(men_men_n311_));
  NAi32      u0283(.An(j), .Bn(h), .C(i), .Y(men_men_n312_));
  NAi21      u0284(.An(m), .B(l), .Y(men_men_n313_));
  NO3        u0285(.A(men_men_n313_), .B(men_men_n312_), .C(men_men_n84_), .Y(men_men_n314_));
  NA2        u0286(.A(h), .B(g), .Y(men_men_n315_));
  NA2        u0287(.A(men_men_n172_), .B(men_men_n45_), .Y(men_men_n316_));
  NO2        u0288(.A(men_men_n316_), .B(men_men_n315_), .Y(men_men_n317_));
  OAI210     u0289(.A0(men_men_n317_), .A1(men_men_n314_), .B0(men_men_n167_), .Y(men_men_n318_));
  NA4        u0290(.A(men_men_n318_), .B(men_men_n311_), .C(men_men_n303_), .D(men_men_n296_), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n148_), .B(d), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n107_), .B(men_men_n104_), .Y(men_men_n321_));
  NAi32      u0293(.An(n), .Bn(m), .C(l), .Y(men_men_n322_));
  NO2        u0294(.A(men_men_n322_), .B(men_men_n312_), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n323_), .B(men_men_n189_), .Y(men_men_n324_));
  NO2        u0296(.A(men_men_n123_), .B(men_men_n117_), .Y(men_men_n325_));
  NAi31      u0297(.An(k), .B(l), .C(j), .Y(men_men_n326_));
  OAI210     u0298(.A0(men_men_n304_), .A1(j), .B0(men_men_n326_), .Y(men_men_n327_));
  NOi21      u0299(.An(men_men_n327_), .B(men_men_n121_), .Y(men_men_n328_));
  NA2        u0300(.A(men_men_n328_), .B(men_men_n325_), .Y(men_men_n329_));
  NA2        u0301(.A(men_men_n329_), .B(men_men_n324_), .Y(men_men_n330_));
  NO4        u0302(.A(men_men_n330_), .B(men_men_n319_), .C(men_men_n292_), .D(men_men_n282_), .Y(men_men_n331_));
  NA2        u0303(.A(men_men_n265_), .B(men_men_n199_), .Y(men_men_n332_));
  NAi21      u0304(.An(m), .B(k), .Y(men_men_n333_));
  NO2        u0305(.A(men_men_n234_), .B(men_men_n333_), .Y(men_men_n334_));
  NAi41      u0306(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n335_));
  NO2        u0307(.A(men_men_n335_), .B(men_men_n154_), .Y(men_men_n336_));
  NA2        u0308(.A(men_men_n336_), .B(men_men_n334_), .Y(men_men_n337_));
  NAi31      u0309(.An(i), .B(l), .C(h), .Y(men_men_n338_));
  NO4        u0310(.A(men_men_n338_), .B(men_men_n154_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n339_));
  NA2        u0311(.A(e), .B(c), .Y(men_men_n340_));
  NO3        u0312(.A(men_men_n340_), .B(n), .C(d), .Y(men_men_n341_));
  NOi21      u0313(.An(f), .B(h), .Y(men_men_n342_));
  NAi31      u0314(.An(d), .B(e), .C(b), .Y(men_men_n343_));
  NO2        u0315(.A(men_men_n134_), .B(men_men_n343_), .Y(men_men_n344_));
  NAi31      u0316(.An(men_men_n339_), .B(men_men_n337_), .C(men_men_n332_), .Y(men_men_n345_));
  NO4        u0317(.A(men_men_n335_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n222_), .Y(men_men_n346_));
  NA2        u0318(.A(men_men_n260_), .B(men_men_n105_), .Y(men_men_n347_));
  OR2        u0319(.A(men_men_n347_), .B(men_men_n211_), .Y(men_men_n348_));
  NOi31      u0320(.An(l), .B(n), .C(m), .Y(men_men_n349_));
  NA2        u0321(.A(men_men_n349_), .B(men_men_n223_), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n350_), .B(men_men_n200_), .Y(men_men_n351_));
  NAi32      u0323(.An(men_men_n351_), .Bn(men_men_n346_), .C(men_men_n348_), .Y(men_men_n352_));
  NAi32      u0324(.An(m), .Bn(j), .C(k), .Y(men_men_n353_));
  NAi41      u0325(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n354_));
  OAI210     u0326(.A0(men_men_n219_), .A1(men_men_n353_), .B0(men_men_n354_), .Y(men_men_n355_));
  NOi31      u0327(.An(j), .B(m), .C(k), .Y(men_men_n356_));
  NO2        u0328(.A(men_men_n127_), .B(men_men_n356_), .Y(men_men_n357_));
  AN3        u0329(.A(h), .B(g), .C(f), .Y(men_men_n358_));
  NAi31      u0330(.An(men_men_n357_), .B(men_men_n358_), .C(men_men_n355_), .Y(men_men_n359_));
  NOi32      u0331(.An(m), .Bn(j), .C(l), .Y(men_men_n360_));
  NO2        u0332(.A(men_men_n360_), .B(men_men_n98_), .Y(men_men_n361_));
  NAi32      u0333(.An(men_men_n361_), .Bn(men_men_n208_), .C(men_men_n320_), .Y(men_men_n362_));
  NO2        u0334(.A(men_men_n313_), .B(men_men_n312_), .Y(men_men_n363_));
  NO2        u0335(.A(men_men_n225_), .B(g), .Y(men_men_n364_));
  NO2        u0336(.A(men_men_n160_), .B(men_men_n84_), .Y(men_men_n365_));
  AOI220     u0337(.A0(men_men_n365_), .A1(men_men_n364_), .B0(men_men_n257_), .B1(men_men_n363_), .Y(men_men_n366_));
  NA2        u0338(.A(men_men_n242_), .B(men_men_n81_), .Y(men_men_n367_));
  NA3        u0339(.A(men_men_n367_), .B(men_men_n358_), .C(men_men_n220_), .Y(men_men_n368_));
  NA4        u0340(.A(men_men_n368_), .B(men_men_n366_), .C(men_men_n362_), .D(men_men_n359_), .Y(men_men_n369_));
  NA3        u0341(.A(h), .B(g), .C(f), .Y(men_men_n370_));
  NO2        u0342(.A(men_men_n370_), .B(men_men_n77_), .Y(men_men_n371_));
  NA2        u0343(.A(men_men_n354_), .B(men_men_n219_), .Y(men_men_n372_));
  NA2        u0344(.A(men_men_n166_), .B(e), .Y(men_men_n373_));
  NO2        u0345(.A(men_men_n373_), .B(men_men_n41_), .Y(men_men_n374_));
  AOI220     u0346(.A0(men_men_n374_), .A1(men_men_n325_), .B0(men_men_n372_), .B1(men_men_n371_), .Y(men_men_n375_));
  NOi32      u0347(.An(j), .Bn(g), .C(i), .Y(men_men_n376_));
  NA3        u0348(.A(men_men_n376_), .B(men_men_n304_), .C(men_men_n114_), .Y(men_men_n377_));
  AO210      u0349(.A0(men_men_n112_), .A1(men_men_n32_), .B0(men_men_n377_), .Y(men_men_n378_));
  NOi32      u0350(.An(e), .Bn(b), .C(a), .Y(men_men_n379_));
  AN2        u0351(.A(l), .B(j), .Y(men_men_n380_));
  NA3        u0352(.A(men_men_n216_), .B(men_men_n214_), .C(men_men_n35_), .Y(men_men_n381_));
  NA2        u0353(.A(men_men_n381_), .B(men_men_n379_), .Y(men_men_n382_));
  NO2        u0354(.A(men_men_n343_), .B(n), .Y(men_men_n383_));
  NA2        u0355(.A(men_men_n215_), .B(k), .Y(men_men_n384_));
  NA3        u0356(.A(m), .B(men_men_n113_), .C(men_men_n221_), .Y(men_men_n385_));
  NA4        u0357(.A(men_men_n210_), .B(men_men_n87_), .C(g), .D(men_men_n221_), .Y(men_men_n386_));
  OAI210     u0358(.A0(men_men_n385_), .A1(men_men_n384_), .B0(men_men_n386_), .Y(men_men_n387_));
  NAi41      u0359(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n388_));
  NA2        u0360(.A(men_men_n51_), .B(men_men_n114_), .Y(men_men_n389_));
  NO2        u0361(.A(men_men_n389_), .B(men_men_n388_), .Y(men_men_n390_));
  AOI220     u0362(.A0(men_men_n390_), .A1(b), .B0(men_men_n387_), .B1(men_men_n383_), .Y(men_men_n391_));
  NA4        u0363(.A(men_men_n391_), .B(men_men_n382_), .C(men_men_n378_), .D(men_men_n375_), .Y(men_men_n392_));
  NO4        u0364(.A(men_men_n392_), .B(men_men_n369_), .C(men_men_n352_), .D(men_men_n345_), .Y(men_men_n393_));
  NA4        u0365(.A(men_men_n393_), .B(men_men_n331_), .C(men_men_n280_), .D(men_men_n206_), .Y(men10));
  NA3        u0366(.A(m), .B(k), .C(i), .Y(men_men_n395_));
  NO3        u0367(.A(men_men_n395_), .B(j), .C(men_men_n222_), .Y(men_men_n396_));
  NOi21      u0368(.An(e), .B(f), .Y(men_men_n397_));
  NO4        u0369(.A(men_men_n155_), .B(men_men_n397_), .C(n), .D(men_men_n111_), .Y(men_men_n398_));
  NAi31      u0370(.An(b), .B(f), .C(c), .Y(men_men_n399_));
  INV        u0371(.A(men_men_n399_), .Y(men_men_n400_));
  NOi32      u0372(.An(k), .Bn(h), .C(j), .Y(men_men_n401_));
  NA2        u0373(.A(men_men_n401_), .B(men_men_n229_), .Y(men_men_n402_));
  NA2        u0374(.A(men_men_n165_), .B(men_men_n402_), .Y(men_men_n403_));
  AOI220     u0375(.A0(men_men_n403_), .A1(men_men_n400_), .B0(men_men_n398_), .B1(men_men_n396_), .Y(men_men_n404_));
  AN2        u0376(.A(j), .B(h), .Y(men_men_n405_));
  NO3        u0377(.A(n), .B(m), .C(k), .Y(men_men_n406_));
  NA2        u0378(.A(men_men_n406_), .B(men_men_n405_), .Y(men_men_n407_));
  NO3        u0379(.A(men_men_n407_), .B(men_men_n155_), .C(men_men_n221_), .Y(men_men_n408_));
  OR2        u0380(.A(m), .B(k), .Y(men_men_n409_));
  NO2        u0381(.A(men_men_n179_), .B(men_men_n409_), .Y(men_men_n410_));
  NA4        u0382(.A(n), .B(f), .C(c), .D(men_men_n117_), .Y(men_men_n411_));
  NOi21      u0383(.An(men_men_n410_), .B(men_men_n411_), .Y(men_men_n412_));
  NOi32      u0384(.An(d), .Bn(a), .C(c), .Y(men_men_n413_));
  NA2        u0385(.A(men_men_n413_), .B(men_men_n187_), .Y(men_men_n414_));
  NAi21      u0386(.An(i), .B(g), .Y(men_men_n415_));
  NAi31      u0387(.An(k), .B(m), .C(j), .Y(men_men_n416_));
  NO3        u0388(.A(men_men_n416_), .B(men_men_n415_), .C(n), .Y(men_men_n417_));
  NOi21      u0389(.An(men_men_n417_), .B(men_men_n414_), .Y(men_men_n418_));
  NO3        u0390(.A(men_men_n418_), .B(men_men_n412_), .C(men_men_n408_), .Y(men_men_n419_));
  NO2        u0391(.A(men_men_n411_), .B(men_men_n313_), .Y(men_men_n420_));
  NOi32      u0392(.An(f), .Bn(d), .C(c), .Y(men_men_n421_));
  AOI220     u0393(.A0(men_men_n421_), .A1(men_men_n323_), .B0(men_men_n420_), .B1(men_men_n223_), .Y(men_men_n422_));
  NA3        u0394(.A(men_men_n422_), .B(men_men_n419_), .C(men_men_n404_), .Y(men_men_n423_));
  NO2        u0395(.A(men_men_n59_), .B(men_men_n117_), .Y(men_men_n424_));
  NA2        u0396(.A(men_men_n260_), .B(men_men_n424_), .Y(men_men_n425_));
  INV        u0397(.A(e), .Y(men_men_n426_));
  NA2        u0398(.A(men_men_n46_), .B(e), .Y(men_men_n427_));
  OAI220     u0399(.A0(men_men_n427_), .A1(men_men_n207_), .B0(men_men_n211_), .B1(men_men_n426_), .Y(men_men_n428_));
  AN2        u0400(.A(g), .B(e), .Y(men_men_n429_));
  NA3        u0401(.A(men_men_n429_), .B(men_men_n210_), .C(i), .Y(men_men_n430_));
  OAI210     u0402(.A0(men_men_n89_), .A1(men_men_n426_), .B0(men_men_n430_), .Y(men_men_n431_));
  NO2        u0403(.A(men_men_n431_), .B(men_men_n428_), .Y(men_men_n432_));
  NOi32      u0404(.An(h), .Bn(e), .C(g), .Y(men_men_n433_));
  NA3        u0405(.A(men_men_n433_), .B(men_men_n306_), .C(m), .Y(men_men_n434_));
  NOi21      u0406(.An(g), .B(h), .Y(men_men_n435_));
  AN3        u0407(.A(m), .B(l), .C(i), .Y(men_men_n436_));
  NA3        u0408(.A(men_men_n436_), .B(men_men_n435_), .C(e), .Y(men_men_n437_));
  AN3        u0409(.A(h), .B(g), .C(e), .Y(men_men_n438_));
  NA2        u0410(.A(men_men_n438_), .B(men_men_n98_), .Y(men_men_n439_));
  NO2        u0411(.A(men_men_n432_), .B(men_men_n425_), .Y(men_men_n440_));
  NA3        u0412(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n441_));
  NO2        u0413(.A(men_men_n441_), .B(men_men_n425_), .Y(men_men_n442_));
  NA3        u0414(.A(men_men_n413_), .B(men_men_n187_), .C(men_men_n84_), .Y(men_men_n443_));
  NAi31      u0415(.An(b), .B(c), .C(a), .Y(men_men_n444_));
  NO2        u0416(.A(men_men_n444_), .B(n), .Y(men_men_n445_));
  OAI210     u0417(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n446_));
  NO2        u0418(.A(men_men_n446_), .B(men_men_n151_), .Y(men_men_n447_));
  NA2        u0419(.A(men_men_n447_), .B(men_men_n445_), .Y(men_men_n448_));
  INV        u0420(.A(men_men_n448_), .Y(men_men_n449_));
  NO4        u0421(.A(men_men_n449_), .B(men_men_n442_), .C(men_men_n440_), .D(men_men_n423_), .Y(men_men_n450_));
  NA2        u0422(.A(i), .B(g), .Y(men_men_n451_));
  NO3        u0423(.A(men_men_n290_), .B(men_men_n451_), .C(c), .Y(men_men_n452_));
  NOi21      u0424(.An(a), .B(n), .Y(men_men_n453_));
  NOi21      u0425(.An(d), .B(c), .Y(men_men_n454_));
  NA2        u0426(.A(men_men_n454_), .B(men_men_n453_), .Y(men_men_n455_));
  NA3        u0427(.A(i), .B(g), .C(f), .Y(men_men_n456_));
  OR2        u0428(.A(men_men_n456_), .B(men_men_n71_), .Y(men_men_n457_));
  NA3        u0429(.A(men_men_n436_), .B(men_men_n435_), .C(men_men_n187_), .Y(men_men_n458_));
  AOI210     u0430(.A0(men_men_n458_), .A1(men_men_n457_), .B0(men_men_n455_), .Y(men_men_n459_));
  AOI210     u0431(.A0(men_men_n452_), .A1(men_men_n305_), .B0(men_men_n459_), .Y(men_men_n460_));
  OR2        u0432(.A(n), .B(m), .Y(men_men_n461_));
  NO2        u0433(.A(men_men_n461_), .B(men_men_n156_), .Y(men_men_n462_));
  NO2        u0434(.A(men_men_n188_), .B(men_men_n151_), .Y(men_men_n463_));
  OAI210     u0435(.A0(men_men_n462_), .A1(men_men_n181_), .B0(men_men_n463_), .Y(men_men_n464_));
  INV        u0436(.A(men_men_n389_), .Y(men_men_n465_));
  NA3        u0437(.A(men_men_n465_), .B(men_men_n379_), .C(d), .Y(men_men_n466_));
  NO2        u0438(.A(men_men_n444_), .B(men_men_n49_), .Y(men_men_n467_));
  NO3        u0439(.A(men_men_n66_), .B(men_men_n113_), .C(e), .Y(men_men_n468_));
  NAi21      u0440(.An(k), .B(j), .Y(men_men_n469_));
  NA3        u0441(.A(i), .B(men_men_n468_), .C(men_men_n467_), .Y(men_men_n470_));
  NAi21      u0442(.An(e), .B(d), .Y(men_men_n471_));
  NO2        u0443(.A(men_men_n471_), .B(men_men_n56_), .Y(men_men_n472_));
  NO2        u0444(.A(men_men_n264_), .B(men_men_n221_), .Y(men_men_n473_));
  NA3        u0445(.A(men_men_n473_), .B(men_men_n472_), .C(men_men_n235_), .Y(men_men_n474_));
  NA4        u0446(.A(men_men_n474_), .B(men_men_n470_), .C(men_men_n466_), .D(men_men_n464_), .Y(men_men_n475_));
  NO2        u0447(.A(men_men_n350_), .B(men_men_n221_), .Y(men_men_n476_));
  NA2        u0448(.A(men_men_n476_), .B(men_men_n472_), .Y(men_men_n477_));
  NOi31      u0449(.An(n), .B(m), .C(k), .Y(men_men_n478_));
  AOI220     u0450(.A0(men_men_n478_), .A1(men_men_n405_), .B0(men_men_n229_), .B1(men_men_n50_), .Y(men_men_n479_));
  NAi31      u0451(.An(g), .B(f), .C(c), .Y(men_men_n480_));
  NA2        u0452(.A(men_men_n477_), .B(men_men_n324_), .Y(men_men_n481_));
  NOi41      u0453(.An(men_men_n460_), .B(men_men_n481_), .C(men_men_n475_), .D(men_men_n278_), .Y(men_men_n482_));
  NOi32      u0454(.An(c), .Bn(a), .C(b), .Y(men_men_n483_));
  NA2        u0455(.A(men_men_n483_), .B(men_men_n114_), .Y(men_men_n484_));
  AN2        u0456(.A(e), .B(d), .Y(men_men_n485_));
  INV        u0457(.A(men_men_n151_), .Y(men_men_n486_));
  NO2        u0458(.A(men_men_n133_), .B(men_men_n41_), .Y(men_men_n487_));
  NO2        u0459(.A(men_men_n66_), .B(e), .Y(men_men_n488_));
  NOi31      u0460(.An(j), .B(k), .C(i), .Y(men_men_n489_));
  NOi21      u0461(.An(men_men_n169_), .B(men_men_n489_), .Y(men_men_n490_));
  NA4        u0462(.A(men_men_n338_), .B(men_men_n490_), .C(men_men_n272_), .D(men_men_n120_), .Y(men_men_n491_));
  NA2        u0463(.A(men_men_n491_), .B(men_men_n488_), .Y(men_men_n492_));
  NO2        u0464(.A(men_men_n492_), .B(men_men_n484_), .Y(men_men_n493_));
  NO2        u0465(.A(men_men_n217_), .B(men_men_n212_), .Y(men_men_n494_));
  NOi21      u0466(.An(a), .B(b), .Y(men_men_n495_));
  NA3        u0467(.A(e), .B(d), .C(c), .Y(men_men_n496_));
  NAi21      u0468(.An(men_men_n496_), .B(men_men_n495_), .Y(men_men_n497_));
  NO2        u0469(.A(men_men_n443_), .B(men_men_n211_), .Y(men_men_n498_));
  NOi21      u0470(.An(men_men_n497_), .B(men_men_n498_), .Y(men_men_n499_));
  AOI210     u0471(.A0(men_men_n281_), .A1(men_men_n494_), .B0(men_men_n499_), .Y(men_men_n500_));
  NO4        u0472(.A(men_men_n194_), .B(men_men_n104_), .C(men_men_n56_), .D(b), .Y(men_men_n501_));
  NA2        u0473(.A(men_men_n400_), .B(men_men_n157_), .Y(men_men_n502_));
  OR2        u0474(.A(k), .B(j), .Y(men_men_n503_));
  NA2        u0475(.A(l), .B(k), .Y(men_men_n504_));
  NA3        u0476(.A(men_men_n504_), .B(men_men_n503_), .C(men_men_n229_), .Y(men_men_n505_));
  AOI210     u0477(.A0(men_men_n242_), .A1(men_men_n353_), .B0(men_men_n84_), .Y(men_men_n506_));
  NOi21      u0478(.An(men_men_n505_), .B(men_men_n506_), .Y(men_men_n507_));
  OR3        u0479(.A(men_men_n507_), .B(men_men_n147_), .C(men_men_n137_), .Y(men_men_n508_));
  NA3        u0480(.A(men_men_n293_), .B(men_men_n130_), .C(men_men_n128_), .Y(men_men_n509_));
  NA2        u0481(.A(men_men_n413_), .B(men_men_n114_), .Y(men_men_n510_));
  NO4        u0482(.A(men_men_n510_), .B(men_men_n95_), .C(men_men_n113_), .D(e), .Y(men_men_n511_));
  NO3        u0483(.A(men_men_n443_), .B(men_men_n92_), .C(men_men_n133_), .Y(men_men_n512_));
  NO4        u0484(.A(men_men_n512_), .B(men_men_n511_), .C(men_men_n509_), .D(men_men_n339_), .Y(men_men_n513_));
  NA3        u0485(.A(men_men_n513_), .B(men_men_n508_), .C(men_men_n502_), .Y(men_men_n514_));
  NO4        u0486(.A(men_men_n514_), .B(men_men_n501_), .C(men_men_n500_), .D(men_men_n493_), .Y(men_men_n515_));
  NA2        u0487(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n516_));
  NOi21      u0488(.An(d), .B(e), .Y(men_men_n517_));
  NO2        u0489(.A(men_men_n194_), .B(men_men_n56_), .Y(men_men_n518_));
  NAi31      u0490(.An(j), .B(l), .C(i), .Y(men_men_n519_));
  OAI210     u0491(.A0(men_men_n519_), .A1(men_men_n134_), .B0(men_men_n104_), .Y(men_men_n520_));
  NA4        u0492(.A(men_men_n520_), .B(men_men_n518_), .C(men_men_n517_), .D(b), .Y(men_men_n521_));
  NO3        u0493(.A(men_men_n414_), .B(men_men_n361_), .C(men_men_n208_), .Y(men_men_n522_));
  NO2        u0494(.A(men_men_n414_), .B(men_men_n389_), .Y(men_men_n523_));
  NO4        u0495(.A(men_men_n523_), .B(men_men_n522_), .C(men_men_n190_), .D(men_men_n321_), .Y(men_men_n524_));
  NA4        u0496(.A(men_men_n524_), .B(men_men_n521_), .C(men_men_n516_), .D(men_men_n252_), .Y(men_men_n525_));
  OAI210     u0497(.A0(men_men_n129_), .A1(men_men_n127_), .B0(n), .Y(men_men_n526_));
  NO2        u0498(.A(men_men_n526_), .B(men_men_n133_), .Y(men_men_n527_));
  OA210      u0499(.A0(men_men_n314_), .A1(men_men_n527_), .B0(men_men_n199_), .Y(men_men_n528_));
  XO2        u0500(.A(i), .B(h), .Y(men_men_n529_));
  NA3        u0501(.A(men_men_n529_), .B(men_men_n164_), .C(n), .Y(men_men_n530_));
  NAi41      u0502(.An(men_men_n314_), .B(men_men_n530_), .C(men_men_n479_), .D(men_men_n402_), .Y(men_men_n531_));
  NOi32      u0503(.An(men_men_n531_), .Bn(men_men_n488_), .C(men_men_n283_), .Y(men_men_n532_));
  NAi31      u0504(.An(c), .B(f), .C(d), .Y(men_men_n533_));
  AOI210     u0505(.A0(men_men_n294_), .A1(men_men_n202_), .B0(men_men_n533_), .Y(men_men_n534_));
  INV        u0506(.A(men_men_n534_), .Y(men_men_n535_));
  NA3        u0507(.A(men_men_n398_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n536_));
  NA2        u0508(.A(men_men_n236_), .B(men_men_n109_), .Y(men_men_n537_));
  AOI210     u0509(.A0(men_men_n537_), .A1(men_men_n186_), .B0(men_men_n533_), .Y(men_men_n538_));
  NOi21      u0510(.An(men_men_n536_), .B(men_men_n538_), .Y(men_men_n539_));
  AO220      u0511(.A0(men_men_n302_), .A1(men_men_n275_), .B0(men_men_n170_), .B1(men_men_n67_), .Y(men_men_n540_));
  NA3        u0512(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n541_), .B(men_men_n455_), .Y(men_men_n542_));
  NO2        u0514(.A(men_men_n542_), .B(men_men_n310_), .Y(men_men_n543_));
  NAi41      u0515(.An(men_men_n540_), .B(men_men_n543_), .C(men_men_n539_), .D(men_men_n535_), .Y(men_men_n544_));
  NO4        u0516(.A(men_men_n544_), .B(men_men_n532_), .C(men_men_n528_), .D(men_men_n525_), .Y(men_men_n545_));
  NA4        u0517(.A(men_men_n545_), .B(men_men_n515_), .C(men_men_n482_), .D(men_men_n450_), .Y(men11));
  NO2        u0518(.A(men_men_n73_), .B(f), .Y(men_men_n547_));
  NA2        u0519(.A(j), .B(g), .Y(men_men_n548_));
  NAi31      u0520(.An(i), .B(m), .C(l), .Y(men_men_n549_));
  NA3        u0521(.A(m), .B(k), .C(j), .Y(men_men_n550_));
  OAI220     u0522(.A0(men_men_n550_), .A1(men_men_n133_), .B0(men_men_n549_), .B1(men_men_n548_), .Y(men_men_n551_));
  NA2        u0523(.A(men_men_n551_), .B(men_men_n547_), .Y(men_men_n552_));
  NOi32      u0524(.An(e), .Bn(b), .C(f), .Y(men_men_n553_));
  NA2        u0525(.A(men_men_n271_), .B(men_men_n114_), .Y(men_men_n554_));
  NA2        u0526(.A(men_men_n46_), .B(j), .Y(men_men_n555_));
  OAI220     u0527(.A0(men_men_n555_), .A1(men_men_n316_), .B0(men_men_n554_), .B1(men_men_n222_), .Y(men_men_n556_));
  NAi31      u0528(.An(d), .B(e), .C(a), .Y(men_men_n557_));
  NO2        u0529(.A(men_men_n557_), .B(n), .Y(men_men_n558_));
  AOI220     u0530(.A0(men_men_n558_), .A1(men_men_n102_), .B0(men_men_n556_), .B1(men_men_n553_), .Y(men_men_n559_));
  NAi41      u0531(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n560_));
  AN2        u0532(.A(men_men_n560_), .B(men_men_n388_), .Y(men_men_n561_));
  AOI210     u0533(.A0(men_men_n561_), .A1(men_men_n414_), .B0(men_men_n284_), .Y(men_men_n562_));
  NA2        u0534(.A(j), .B(i), .Y(men_men_n563_));
  NAi31      u0535(.An(n), .B(m), .C(k), .Y(men_men_n564_));
  NO3        u0536(.A(men_men_n564_), .B(men_men_n563_), .C(men_men_n113_), .Y(men_men_n565_));
  NO4        u0537(.A(n), .B(d), .C(men_men_n117_), .D(a), .Y(men_men_n566_));
  OR2        u0538(.A(n), .B(c), .Y(men_men_n567_));
  NO2        u0539(.A(men_men_n567_), .B(men_men_n153_), .Y(men_men_n568_));
  NO2        u0540(.A(men_men_n568_), .B(men_men_n566_), .Y(men_men_n569_));
  NOi32      u0541(.An(g), .Bn(f), .C(i), .Y(men_men_n570_));
  AOI220     u0542(.A0(men_men_n570_), .A1(men_men_n100_), .B0(men_men_n551_), .B1(f), .Y(men_men_n571_));
  NO2        u0543(.A(men_men_n288_), .B(men_men_n49_), .Y(men_men_n572_));
  NO2        u0544(.A(men_men_n571_), .B(men_men_n569_), .Y(men_men_n573_));
  AOI210     u0545(.A0(men_men_n565_), .A1(men_men_n562_), .B0(men_men_n573_), .Y(men_men_n574_));
  NA2        u0546(.A(men_men_n143_), .B(men_men_n34_), .Y(men_men_n575_));
  OAI220     u0547(.A0(men_men_n575_), .A1(m), .B0(men_men_n555_), .B1(men_men_n242_), .Y(men_men_n576_));
  NOi41      u0548(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n577_));
  NAi32      u0549(.An(e), .Bn(b), .C(c), .Y(men_men_n578_));
  OR2        u0550(.A(men_men_n578_), .B(men_men_n84_), .Y(men_men_n579_));
  AN2        u0551(.A(men_men_n354_), .B(men_men_n335_), .Y(men_men_n580_));
  NA2        u0552(.A(men_men_n580_), .B(men_men_n579_), .Y(men_men_n581_));
  OA210      u0553(.A0(men_men_n581_), .A1(men_men_n577_), .B0(men_men_n576_), .Y(men_men_n582_));
  OAI220     u0554(.A0(men_men_n416_), .A1(men_men_n415_), .B0(men_men_n549_), .B1(men_men_n548_), .Y(men_men_n583_));
  NAi31      u0555(.An(d), .B(c), .C(a), .Y(men_men_n584_));
  NO2        u0556(.A(men_men_n584_), .B(n), .Y(men_men_n585_));
  NA3        u0557(.A(men_men_n585_), .B(men_men_n583_), .C(e), .Y(men_men_n586_));
  NO3        u0558(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n222_), .Y(men_men_n587_));
  NO2        u0559(.A(men_men_n239_), .B(men_men_n111_), .Y(men_men_n588_));
  OAI210     u0560(.A0(men_men_n587_), .A1(men_men_n417_), .B0(men_men_n588_), .Y(men_men_n589_));
  NA2        u0561(.A(men_men_n589_), .B(men_men_n586_), .Y(men_men_n590_));
  NO2        u0562(.A(men_men_n290_), .B(n), .Y(men_men_n591_));
  NO2        u0563(.A(men_men_n445_), .B(men_men_n591_), .Y(men_men_n592_));
  NA2        u0564(.A(men_men_n583_), .B(f), .Y(men_men_n593_));
  NAi32      u0565(.An(d), .Bn(a), .C(b), .Y(men_men_n594_));
  NO2        u0566(.A(men_men_n594_), .B(men_men_n49_), .Y(men_men_n595_));
  NA2        u0567(.A(h), .B(f), .Y(men_men_n596_));
  NO2        u0568(.A(men_men_n596_), .B(men_men_n95_), .Y(men_men_n597_));
  NO3        u0569(.A(men_men_n182_), .B(men_men_n179_), .C(g), .Y(men_men_n598_));
  AOI220     u0570(.A0(men_men_n598_), .A1(men_men_n58_), .B0(men_men_n597_), .B1(men_men_n595_), .Y(men_men_n599_));
  OAI210     u0571(.A0(men_men_n593_), .A1(men_men_n592_), .B0(men_men_n599_), .Y(men_men_n600_));
  AN3        u0572(.A(j), .B(h), .C(g), .Y(men_men_n601_));
  NO2        u0573(.A(men_men_n150_), .B(c), .Y(men_men_n602_));
  NA3        u0574(.A(men_men_n602_), .B(men_men_n601_), .C(men_men_n478_), .Y(men_men_n603_));
  NA3        u0575(.A(f), .B(d), .C(b), .Y(men_men_n604_));
  NO4        u0576(.A(men_men_n604_), .B(men_men_n182_), .C(men_men_n179_), .D(g), .Y(men_men_n605_));
  NAi21      u0577(.An(men_men_n605_), .B(men_men_n603_), .Y(men_men_n606_));
  NO4        u0578(.A(men_men_n606_), .B(men_men_n600_), .C(men_men_n590_), .D(men_men_n582_), .Y(men_men_n607_));
  AN4        u0579(.A(men_men_n607_), .B(men_men_n574_), .C(men_men_n559_), .D(men_men_n552_), .Y(men_men_n608_));
  INV        u0580(.A(k), .Y(men_men_n609_));
  NA3        u0581(.A(l), .B(men_men_n609_), .C(i), .Y(men_men_n610_));
  INV        u0582(.A(men_men_n610_), .Y(men_men_n611_));
  NA4        u0583(.A(men_men_n413_), .B(men_men_n435_), .C(men_men_n187_), .D(men_men_n114_), .Y(men_men_n612_));
  NAi32      u0584(.An(h), .Bn(f), .C(g), .Y(men_men_n613_));
  NAi41      u0585(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n614_));
  OAI210     u0586(.A0(men_men_n557_), .A1(n), .B0(men_men_n614_), .Y(men_men_n615_));
  NA2        u0587(.A(men_men_n615_), .B(m), .Y(men_men_n616_));
  NAi31      u0588(.An(h), .B(g), .C(f), .Y(men_men_n617_));
  OR3        u0589(.A(men_men_n617_), .B(men_men_n290_), .C(men_men_n49_), .Y(men_men_n618_));
  NA4        u0590(.A(men_men_n435_), .B(men_men_n122_), .C(men_men_n114_), .D(e), .Y(men_men_n619_));
  AN2        u0591(.A(men_men_n619_), .B(men_men_n618_), .Y(men_men_n620_));
  OA210      u0592(.A0(men_men_n616_), .A1(men_men_n613_), .B0(men_men_n620_), .Y(men_men_n621_));
  NO3        u0593(.A(men_men_n613_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n622_));
  NO4        u0594(.A(men_men_n617_), .B(men_men_n567_), .C(men_men_n153_), .D(men_men_n75_), .Y(men_men_n623_));
  OR2        u0595(.A(men_men_n623_), .B(men_men_n622_), .Y(men_men_n624_));
  NAi31      u0596(.An(men_men_n624_), .B(men_men_n621_), .C(men_men_n612_), .Y(men_men_n625_));
  NAi31      u0597(.An(f), .B(h), .C(g), .Y(men_men_n626_));
  NO4        u0598(.A(men_men_n326_), .B(men_men_n626_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n627_));
  NOi32      u0599(.An(b), .Bn(a), .C(c), .Y(men_men_n628_));
  NOi41      u0600(.An(men_men_n628_), .B(men_men_n370_), .C(men_men_n69_), .D(men_men_n118_), .Y(men_men_n629_));
  OR2        u0601(.A(men_men_n629_), .B(men_men_n627_), .Y(men_men_n630_));
  NOi32      u0602(.An(d), .Bn(a), .C(e), .Y(men_men_n631_));
  NA2        u0603(.A(men_men_n631_), .B(men_men_n114_), .Y(men_men_n632_));
  NO2        u0604(.A(n), .B(c), .Y(men_men_n633_));
  NA3        u0605(.A(men_men_n633_), .B(men_men_n29_), .C(m), .Y(men_men_n634_));
  NAi32      u0606(.An(n), .Bn(f), .C(m), .Y(men_men_n635_));
  NA3        u0607(.A(men_men_n635_), .B(men_men_n634_), .C(men_men_n632_), .Y(men_men_n636_));
  NOi32      u0608(.An(e), .Bn(a), .C(d), .Y(men_men_n637_));
  AOI210     u0609(.A0(men_men_n29_), .A1(d), .B0(men_men_n637_), .Y(men_men_n638_));
  AOI210     u0610(.A0(men_men_n638_), .A1(men_men_n221_), .B0(men_men_n575_), .Y(men_men_n639_));
  AOI210     u0611(.A0(men_men_n639_), .A1(men_men_n636_), .B0(men_men_n630_), .Y(men_men_n640_));
  OAI210     u0612(.A0(men_men_n259_), .A1(men_men_n87_), .B0(men_men_n640_), .Y(men_men_n641_));
  AOI210     u0613(.A0(men_men_n625_), .A1(men_men_n611_), .B0(men_men_n641_), .Y(men_men_n642_));
  NO3        u0614(.A(men_men_n333_), .B(men_men_n61_), .C(n), .Y(men_men_n643_));
  NA3        u0615(.A(men_men_n533_), .B(men_men_n177_), .C(men_men_n176_), .Y(men_men_n644_));
  NA2        u0616(.A(men_men_n480_), .B(men_men_n239_), .Y(men_men_n645_));
  OR2        u0617(.A(men_men_n645_), .B(men_men_n644_), .Y(men_men_n646_));
  NA2        u0618(.A(men_men_n76_), .B(men_men_n114_), .Y(men_men_n647_));
  NO2        u0619(.A(men_men_n647_), .B(men_men_n45_), .Y(men_men_n648_));
  AOI220     u0620(.A0(men_men_n648_), .A1(men_men_n562_), .B0(men_men_n646_), .B1(men_men_n643_), .Y(men_men_n649_));
  NO2        u0621(.A(men_men_n649_), .B(men_men_n87_), .Y(men_men_n650_));
  NA3        u0622(.A(men_men_n577_), .B(men_men_n356_), .C(men_men_n46_), .Y(men_men_n651_));
  NOi32      u0623(.An(e), .Bn(c), .C(f), .Y(men_men_n652_));
  NOi21      u0624(.An(f), .B(g), .Y(men_men_n653_));
  NO2        u0625(.A(men_men_n653_), .B(men_men_n219_), .Y(men_men_n654_));
  AOI220     u0626(.A0(men_men_n654_), .A1(men_men_n410_), .B0(men_men_n652_), .B1(men_men_n181_), .Y(men_men_n655_));
  NA3        u0627(.A(men_men_n655_), .B(men_men_n651_), .C(men_men_n184_), .Y(men_men_n656_));
  AOI210     u0628(.A0(men_men_n561_), .A1(men_men_n414_), .B0(men_men_n315_), .Y(men_men_n657_));
  NA2        u0629(.A(men_men_n657_), .B(men_men_n276_), .Y(men_men_n658_));
  NOi21      u0630(.An(j), .B(l), .Y(men_men_n659_));
  NAi21      u0631(.An(k), .B(h), .Y(men_men_n660_));
  NO2        u0632(.A(men_men_n660_), .B(men_men_n274_), .Y(men_men_n661_));
  NA2        u0633(.A(men_men_n661_), .B(men_men_n659_), .Y(men_men_n662_));
  OR2        u0634(.A(men_men_n662_), .B(men_men_n616_), .Y(men_men_n663_));
  NOi31      u0635(.An(m), .B(n), .C(k), .Y(men_men_n664_));
  NA2        u0636(.A(men_men_n659_), .B(men_men_n664_), .Y(men_men_n665_));
  AOI210     u0637(.A0(men_men_n414_), .A1(men_men_n388_), .B0(men_men_n315_), .Y(men_men_n666_));
  NAi21      u0638(.An(men_men_n665_), .B(men_men_n666_), .Y(men_men_n667_));
  NO2        u0639(.A(men_men_n290_), .B(men_men_n49_), .Y(men_men_n668_));
  NO2        u0640(.A(men_men_n326_), .B(men_men_n626_), .Y(men_men_n669_));
  NO2        u0641(.A(men_men_n557_), .B(men_men_n49_), .Y(men_men_n670_));
  AOI220     u0642(.A0(men_men_n670_), .A1(men_men_n669_), .B0(men_men_n668_), .B1(men_men_n597_), .Y(men_men_n671_));
  NA4        u0643(.A(men_men_n671_), .B(men_men_n667_), .C(men_men_n663_), .D(men_men_n658_), .Y(men_men_n672_));
  NA2        u0644(.A(men_men_n109_), .B(men_men_n36_), .Y(men_men_n673_));
  NO2        u0645(.A(k), .B(men_men_n222_), .Y(men_men_n674_));
  NO2        u0646(.A(men_men_n553_), .B(men_men_n379_), .Y(men_men_n675_));
  NO2        u0647(.A(men_men_n555_), .B(men_men_n182_), .Y(men_men_n676_));
  NA3        u0648(.A(men_men_n578_), .B(men_men_n283_), .C(men_men_n148_), .Y(men_men_n677_));
  NA2        u0649(.A(men_men_n529_), .B(men_men_n164_), .Y(men_men_n678_));
  NO3        u0650(.A(men_men_n411_), .B(men_men_n678_), .C(men_men_n87_), .Y(men_men_n679_));
  AOI210     u0651(.A0(men_men_n677_), .A1(men_men_n676_), .B0(men_men_n679_), .Y(men_men_n680_));
  AN3        u0652(.A(f), .B(d), .C(b), .Y(men_men_n681_));
  OAI210     u0653(.A0(men_men_n681_), .A1(men_men_n132_), .B0(n), .Y(men_men_n682_));
  NA3        u0654(.A(men_men_n529_), .B(men_men_n164_), .C(men_men_n222_), .Y(men_men_n683_));
  AOI210     u0655(.A0(men_men_n682_), .A1(men_men_n241_), .B0(men_men_n683_), .Y(men_men_n684_));
  NAi31      u0656(.An(m), .B(n), .C(k), .Y(men_men_n685_));
  OR2        u0657(.A(men_men_n137_), .B(men_men_n61_), .Y(men_men_n686_));
  OAI210     u0658(.A0(men_men_n686_), .A1(men_men_n685_), .B0(men_men_n261_), .Y(men_men_n687_));
  OAI210     u0659(.A0(men_men_n687_), .A1(men_men_n684_), .B0(j), .Y(men_men_n688_));
  NA2        u0660(.A(men_men_n688_), .B(men_men_n680_), .Y(men_men_n689_));
  NO4        u0661(.A(men_men_n689_), .B(men_men_n672_), .C(men_men_n656_), .D(men_men_n650_), .Y(men_men_n690_));
  NA2        u0662(.A(men_men_n398_), .B(men_men_n166_), .Y(men_men_n691_));
  NAi31      u0663(.An(g), .B(h), .C(f), .Y(men_men_n692_));
  OR3        u0664(.A(men_men_n692_), .B(men_men_n290_), .C(n), .Y(men_men_n693_));
  OA210      u0665(.A0(men_men_n557_), .A1(n), .B0(men_men_n614_), .Y(men_men_n694_));
  NA3        u0666(.A(men_men_n433_), .B(men_men_n122_), .C(men_men_n84_), .Y(men_men_n695_));
  OAI210     u0667(.A0(men_men_n694_), .A1(men_men_n91_), .B0(men_men_n695_), .Y(men_men_n696_));
  NOi21      u0668(.An(men_men_n693_), .B(men_men_n696_), .Y(men_men_n697_));
  AOI210     u0669(.A0(men_men_n697_), .A1(men_men_n691_), .B0(men_men_n550_), .Y(men_men_n698_));
  NO3        u0670(.A(g), .B(men_men_n221_), .C(men_men_n56_), .Y(men_men_n699_));
  NAi21      u0671(.An(h), .B(j), .Y(men_men_n700_));
  NA2        u0672(.A(men_men_n410_), .B(men_men_n699_), .Y(men_men_n701_));
  OR2        u0673(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n628_), .B(men_men_n358_), .Y(men_men_n703_));
  OA220      u0675(.A0(men_men_n665_), .A1(men_men_n703_), .B0(men_men_n662_), .B1(men_men_n702_), .Y(men_men_n704_));
  NA3        u0676(.A(men_men_n547_), .B(men_men_n100_), .C(men_men_n99_), .Y(men_men_n705_));
  AN2        u0677(.A(h), .B(f), .Y(men_men_n706_));
  NA2        u0678(.A(men_men_n706_), .B(men_men_n37_), .Y(men_men_n707_));
  NO2        u0679(.A(men_men_n707_), .B(men_men_n484_), .Y(men_men_n708_));
  AOI210     u0680(.A0(men_men_n594_), .A1(men_men_n444_), .B0(men_men_n49_), .Y(men_men_n709_));
  INV        u0681(.A(men_men_n708_), .Y(men_men_n710_));
  NA4        u0682(.A(men_men_n710_), .B(men_men_n705_), .C(men_men_n704_), .D(men_men_n701_), .Y(men_men_n711_));
  NO2        u0683(.A(men_men_n263_), .B(f), .Y(men_men_n712_));
  INV        u0684(.A(men_men_n61_), .Y(men_men_n713_));
  NO3        u0685(.A(men_men_n713_), .B(men_men_n712_), .C(men_men_n34_), .Y(men_men_n714_));
  NA2        u0686(.A(men_men_n344_), .B(men_men_n143_), .Y(men_men_n715_));
  NA2        u0687(.A(men_men_n134_), .B(men_men_n49_), .Y(men_men_n716_));
  AOI220     u0688(.A0(men_men_n716_), .A1(men_men_n553_), .B0(men_men_n379_), .B1(men_men_n114_), .Y(men_men_n717_));
  OA220      u0689(.A0(men_men_n717_), .A1(men_men_n575_), .B0(men_men_n377_), .B1(men_men_n112_), .Y(men_men_n718_));
  OAI210     u0690(.A0(men_men_n715_), .A1(men_men_n714_), .B0(men_men_n718_), .Y(men_men_n719_));
  NO3        u0691(.A(men_men_n421_), .B(men_men_n199_), .C(men_men_n198_), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n720_), .B(men_men_n239_), .Y(men_men_n721_));
  NA3        u0693(.A(men_men_n721_), .B(men_men_n265_), .C(j), .Y(men_men_n722_));
  NO3        u0694(.A(men_men_n480_), .B(men_men_n179_), .C(i), .Y(men_men_n723_));
  NA2        u0695(.A(men_men_n483_), .B(men_men_n84_), .Y(men_men_n724_));
  NO4        u0696(.A(men_men_n550_), .B(men_men_n724_), .C(men_men_n133_), .D(men_men_n221_), .Y(men_men_n725_));
  INV        u0697(.A(men_men_n725_), .Y(men_men_n726_));
  NA4        u0698(.A(men_men_n726_), .B(men_men_n722_), .C(men_men_n536_), .D(men_men_n419_), .Y(men_men_n727_));
  NO4        u0699(.A(men_men_n727_), .B(men_men_n719_), .C(men_men_n711_), .D(men_men_n698_), .Y(men_men_n728_));
  NA4        u0700(.A(men_men_n728_), .B(men_men_n690_), .C(men_men_n642_), .D(men_men_n608_), .Y(men08));
  NO2        u0701(.A(k), .B(h), .Y(men_men_n730_));
  AO210      u0702(.A0(men_men_n263_), .A1(men_men_n469_), .B0(men_men_n730_), .Y(men_men_n731_));
  NO2        u0703(.A(men_men_n731_), .B(men_men_n313_), .Y(men_men_n732_));
  NA2        u0704(.A(men_men_n652_), .B(men_men_n84_), .Y(men_men_n733_));
  NA2        u0705(.A(men_men_n733_), .B(men_men_n480_), .Y(men_men_n734_));
  AOI210     u0706(.A0(men_men_n734_), .A1(men_men_n732_), .B0(men_men_n512_), .Y(men_men_n735_));
  NA2        u0707(.A(men_men_n84_), .B(men_men_n111_), .Y(men_men_n736_));
  NO2        u0708(.A(men_men_n736_), .B(men_men_n57_), .Y(men_men_n737_));
  NA2        u0709(.A(men_men_n604_), .B(men_men_n241_), .Y(men_men_n738_));
  AOI210     u0710(.A0(men_men_n604_), .A1(men_men_n160_), .B0(men_men_n84_), .Y(men_men_n739_));
  NA4        u0711(.A(men_men_n224_), .B(men_men_n143_), .C(men_men_n45_), .D(h), .Y(men_men_n740_));
  AN2        u0712(.A(l), .B(k), .Y(men_men_n741_));
  NA4        u0713(.A(men_men_n741_), .B(men_men_n109_), .C(men_men_n75_), .D(men_men_n222_), .Y(men_men_n742_));
  INV        u0714(.A(men_men_n742_), .Y(men_men_n743_));
  NA2        u0715(.A(men_men_n743_), .B(men_men_n739_), .Y(men_men_n744_));
  NA3        u0716(.A(men_men_n744_), .B(men_men_n735_), .C(men_men_n366_), .Y(men_men_n745_));
  AN2        u0717(.A(men_men_n558_), .B(men_men_n96_), .Y(men_men_n746_));
  NO4        u0718(.A(men_men_n179_), .B(men_men_n409_), .C(men_men_n113_), .D(g), .Y(men_men_n747_));
  AOI210     u0719(.A0(men_men_n747_), .A1(men_men_n738_), .B0(men_men_n542_), .Y(men_men_n748_));
  NO2        u0720(.A(men_men_n38_), .B(men_men_n221_), .Y(men_men_n749_));
  AOI220     u0721(.A0(men_men_n654_), .A1(men_men_n363_), .B0(men_men_n749_), .B1(men_men_n591_), .Y(men_men_n750_));
  NAi31      u0722(.An(men_men_n746_), .B(men_men_n750_), .C(men_men_n748_), .Y(men_men_n751_));
  NO2        u0723(.A(men_men_n561_), .B(men_men_n35_), .Y(men_men_n752_));
  OAI210     u0724(.A0(men_men_n578_), .A1(men_men_n47_), .B0(men_men_n686_), .Y(men_men_n753_));
  NO2        u0725(.A(men_men_n504_), .B(men_men_n134_), .Y(men_men_n754_));
  AOI210     u0726(.A0(men_men_n754_), .A1(men_men_n753_), .B0(men_men_n752_), .Y(men_men_n755_));
  NO3        u0727(.A(men_men_n333_), .B(men_men_n133_), .C(men_men_n41_), .Y(men_men_n756_));
  NAi21      u0728(.An(men_men_n756_), .B(men_men_n742_), .Y(men_men_n757_));
  NA2        u0729(.A(men_men_n731_), .B(men_men_n138_), .Y(men_men_n758_));
  AOI220     u0730(.A0(men_men_n758_), .A1(men_men_n420_), .B0(men_men_n757_), .B1(men_men_n78_), .Y(men_men_n759_));
  OAI210     u0731(.A0(men_men_n755_), .A1(men_men_n87_), .B0(men_men_n759_), .Y(men_men_n760_));
  NA3        u0732(.A(men_men_n721_), .B(men_men_n349_), .C(men_men_n401_), .Y(men_men_n761_));
  NA2        u0733(.A(men_men_n741_), .B(men_men_n229_), .Y(men_men_n762_));
  NO2        u0734(.A(men_men_n762_), .B(men_men_n343_), .Y(men_men_n763_));
  AOI210     u0735(.A0(men_men_n763_), .A1(men_men_n712_), .B0(men_men_n511_), .Y(men_men_n764_));
  NA3        u0736(.A(m), .B(l), .C(k), .Y(men_men_n765_));
  AOI210     u0737(.A0(men_men_n695_), .A1(men_men_n693_), .B0(men_men_n765_), .Y(men_men_n766_));
  NO2        u0738(.A(men_men_n560_), .B(men_men_n284_), .Y(men_men_n767_));
  NOi21      u0739(.An(men_men_n767_), .B(men_men_n554_), .Y(men_men_n768_));
  NA4        u0740(.A(men_men_n114_), .B(l), .C(k), .D(men_men_n87_), .Y(men_men_n769_));
  NA3        u0741(.A(men_men_n122_), .B(men_men_n429_), .C(i), .Y(men_men_n770_));
  NO2        u0742(.A(men_men_n770_), .B(men_men_n769_), .Y(men_men_n771_));
  NO3        u0743(.A(men_men_n771_), .B(men_men_n768_), .C(men_men_n766_), .Y(men_men_n772_));
  NA3        u0744(.A(men_men_n772_), .B(men_men_n764_), .C(men_men_n761_), .Y(men_men_n773_));
  NO4        u0745(.A(men_men_n773_), .B(men_men_n760_), .C(men_men_n751_), .D(men_men_n745_), .Y(men_men_n774_));
  NA2        u0746(.A(men_men_n654_), .B(men_men_n410_), .Y(men_men_n775_));
  NOi31      u0747(.An(g), .B(h), .C(f), .Y(men_men_n776_));
  NA2        u0748(.A(men_men_n670_), .B(men_men_n776_), .Y(men_men_n777_));
  AO210      u0749(.A0(men_men_n777_), .A1(men_men_n618_), .B0(men_men_n563_), .Y(men_men_n778_));
  NO3        u0750(.A(men_men_n414_), .B(men_men_n548_), .C(h), .Y(men_men_n779_));
  AOI210     u0751(.A0(men_men_n779_), .A1(men_men_n114_), .B0(men_men_n523_), .Y(men_men_n780_));
  NA4        u0752(.A(men_men_n780_), .B(men_men_n778_), .C(men_men_n775_), .D(men_men_n262_), .Y(men_men_n781_));
  NA2        u0753(.A(men_men_n741_), .B(men_men_n75_), .Y(men_men_n782_));
  NO4        u0754(.A(men_men_n720_), .B(men_men_n179_), .C(n), .D(i), .Y(men_men_n783_));
  NOi21      u0755(.An(h), .B(j), .Y(men_men_n784_));
  NA2        u0756(.A(men_men_n784_), .B(f), .Y(men_men_n785_));
  NO2        u0757(.A(men_men_n785_), .B(men_men_n256_), .Y(men_men_n786_));
  NO3        u0758(.A(men_men_n786_), .B(men_men_n783_), .C(men_men_n723_), .Y(men_men_n787_));
  OAI220     u0759(.A0(men_men_n787_), .A1(men_men_n782_), .B0(men_men_n620_), .B1(men_men_n62_), .Y(men_men_n788_));
  AOI210     u0760(.A0(men_men_n781_), .A1(l), .B0(men_men_n788_), .Y(men_men_n789_));
  NO2        u0761(.A(j), .B(i), .Y(men_men_n790_));
  NA3        u0762(.A(men_men_n790_), .B(men_men_n82_), .C(l), .Y(men_men_n791_));
  NA2        u0763(.A(men_men_n790_), .B(men_men_n33_), .Y(men_men_n792_));
  NA2        u0764(.A(men_men_n438_), .B(men_men_n122_), .Y(men_men_n793_));
  OA220      u0765(.A0(men_men_n793_), .A1(men_men_n792_), .B0(men_men_n791_), .B1(men_men_n616_), .Y(men_men_n794_));
  NO3        u0766(.A(men_men_n155_), .B(men_men_n49_), .C(men_men_n111_), .Y(men_men_n795_));
  NO3        u0767(.A(men_men_n567_), .B(men_men_n153_), .C(men_men_n75_), .Y(men_men_n796_));
  NO3        u0768(.A(men_men_n504_), .B(men_men_n456_), .C(j), .Y(men_men_n797_));
  OAI210     u0769(.A0(men_men_n796_), .A1(men_men_n795_), .B0(men_men_n797_), .Y(men_men_n798_));
  OAI210     u0770(.A0(men_men_n777_), .A1(men_men_n62_), .B0(men_men_n798_), .Y(men_men_n799_));
  NA2        u0771(.A(k), .B(j), .Y(men_men_n800_));
  AOI210     u0772(.A0(men_men_n553_), .A1(n), .B0(men_men_n577_), .Y(men_men_n801_));
  NA2        u0773(.A(men_men_n801_), .B(men_men_n580_), .Y(men_men_n802_));
  NO3        u0774(.A(men_men_n179_), .B(men_men_n409_), .C(men_men_n113_), .Y(men_men_n803_));
  AOI220     u0775(.A0(men_men_n803_), .A1(men_men_n257_), .B0(men_men_n645_), .B1(men_men_n323_), .Y(men_men_n804_));
  NAi31      u0776(.An(men_men_n638_), .B(men_men_n93_), .C(men_men_n84_), .Y(men_men_n805_));
  NA2        u0777(.A(men_men_n805_), .B(men_men_n804_), .Y(men_men_n806_));
  NO2        u0778(.A(men_men_n313_), .B(men_men_n138_), .Y(men_men_n807_));
  AOI220     u0779(.A0(men_men_n807_), .A1(men_men_n654_), .B0(men_men_n756_), .B1(men_men_n739_), .Y(men_men_n808_));
  NO2        u0780(.A(men_men_n765_), .B(men_men_n91_), .Y(men_men_n809_));
  NA2        u0781(.A(men_men_n797_), .B(men_men_n709_), .Y(men_men_n810_));
  NA2        u0782(.A(men_men_n810_), .B(men_men_n808_), .Y(men_men_n811_));
  OR3        u0783(.A(men_men_n811_), .B(men_men_n806_), .C(men_men_n799_), .Y(men_men_n812_));
  NA3        u0784(.A(men_men_n801_), .B(men_men_n580_), .C(men_men_n579_), .Y(men_men_n813_));
  NA4        u0785(.A(men_men_n813_), .B(men_men_n224_), .C(men_men_n469_), .D(men_men_n34_), .Y(men_men_n814_));
  NO4        u0786(.A(men_men_n504_), .B(men_men_n451_), .C(j), .D(f), .Y(men_men_n815_));
  OAI220     u0787(.A0(men_men_n740_), .A1(men_men_n733_), .B0(men_men_n347_), .B1(men_men_n38_), .Y(men_men_n816_));
  AOI210     u0788(.A0(men_men_n815_), .A1(men_men_n269_), .B0(men_men_n816_), .Y(men_men_n817_));
  NA3        u0789(.A(men_men_n570_), .B(men_men_n306_), .C(h), .Y(men_men_n818_));
  NOi21      u0790(.An(men_men_n709_), .B(men_men_n818_), .Y(men_men_n819_));
  OAI220     u0791(.A0(men_men_n818_), .A1(men_men_n634_), .B0(men_men_n791_), .B1(men_men_n702_), .Y(men_men_n820_));
  INV        u0792(.A(men_men_n820_), .Y(men_men_n821_));
  NAi41      u0793(.An(men_men_n819_), .B(men_men_n821_), .C(men_men_n817_), .D(men_men_n814_), .Y(men_men_n822_));
  OR2        u0794(.A(men_men_n809_), .B(men_men_n96_), .Y(men_men_n823_));
  AOI220     u0795(.A0(men_men_n823_), .A1(men_men_n247_), .B0(men_men_n797_), .B1(men_men_n668_), .Y(men_men_n824_));
  NO2        u0796(.A(men_men_n694_), .B(men_men_n75_), .Y(men_men_n825_));
  AOI210     u0797(.A0(men_men_n815_), .A1(men_men_n825_), .B0(men_men_n351_), .Y(men_men_n826_));
  OAI210     u0798(.A0(men_men_n765_), .A1(men_men_n692_), .B0(men_men_n541_), .Y(men_men_n827_));
  NA3        u0799(.A(men_men_n260_), .B(men_men_n59_), .C(b), .Y(men_men_n828_));
  AOI220     u0800(.A0(men_men_n633_), .A1(men_men_n29_), .B0(men_men_n483_), .B1(men_men_n84_), .Y(men_men_n829_));
  NA2        u0801(.A(men_men_n829_), .B(men_men_n828_), .Y(men_men_n830_));
  NO2        u0802(.A(men_men_n818_), .B(men_men_n510_), .Y(men_men_n831_));
  AOI210     u0803(.A0(men_men_n830_), .A1(men_men_n827_), .B0(men_men_n831_), .Y(men_men_n832_));
  NA3        u0804(.A(men_men_n832_), .B(men_men_n826_), .C(men_men_n824_), .Y(men_men_n833_));
  NOi41      u0805(.An(men_men_n794_), .B(men_men_n833_), .C(men_men_n822_), .D(men_men_n812_), .Y(men_men_n834_));
  OR3        u0806(.A(men_men_n740_), .B(men_men_n241_), .C(g), .Y(men_men_n835_));
  NO3        u0807(.A(men_men_n357_), .B(men_men_n315_), .C(men_men_n113_), .Y(men_men_n836_));
  NA2        u0808(.A(men_men_n836_), .B(men_men_n802_), .Y(men_men_n837_));
  NA2        u0809(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n838_));
  NO3        u0810(.A(men_men_n838_), .B(men_men_n792_), .C(men_men_n290_), .Y(men_men_n839_));
  INV        u0811(.A(men_men_n839_), .Y(men_men_n840_));
  NA4        u0812(.A(men_men_n840_), .B(men_men_n837_), .C(men_men_n835_), .D(men_men_n422_), .Y(men_men_n841_));
  OR2        u0813(.A(men_men_n692_), .B(men_men_n92_), .Y(men_men_n842_));
  NOi31      u0814(.An(b), .B(d), .C(a), .Y(men_men_n843_));
  NO2        u0815(.A(men_men_n843_), .B(men_men_n631_), .Y(men_men_n844_));
  NO2        u0816(.A(men_men_n844_), .B(n), .Y(men_men_n845_));
  NOi21      u0817(.An(men_men_n829_), .B(men_men_n845_), .Y(men_men_n846_));
  OAI220     u0818(.A0(men_men_n846_), .A1(men_men_n842_), .B0(men_men_n818_), .B1(men_men_n632_), .Y(men_men_n847_));
  NO2        u0819(.A(men_men_n343_), .B(men_men_n118_), .Y(men_men_n848_));
  NOi21      u0820(.An(men_men_n848_), .B(men_men_n165_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n720_), .B(n), .Y(men_men_n850_));
  AOI220     u0822(.A0(men_men_n807_), .A1(men_men_n699_), .B0(men_men_n850_), .B1(men_men_n732_), .Y(men_men_n851_));
  NO2        u0823(.A(men_men_n340_), .B(men_men_n246_), .Y(men_men_n852_));
  OAI210     u0824(.A0(men_men_n96_), .A1(men_men_n93_), .B0(men_men_n852_), .Y(men_men_n853_));
  NA2        u0825(.A(men_men_n122_), .B(men_men_n84_), .Y(men_men_n854_));
  AOI210     u0826(.A0(men_men_n441_), .A1(men_men_n434_), .B0(men_men_n854_), .Y(men_men_n855_));
  NAi21      u0827(.An(men_men_n855_), .B(men_men_n853_), .Y(men_men_n856_));
  NA2        u0828(.A(men_men_n763_), .B(men_men_n34_), .Y(men_men_n857_));
  NAi21      u0829(.An(men_men_n769_), .B(men_men_n452_), .Y(men_men_n858_));
  NO2        u0830(.A(men_men_n284_), .B(i), .Y(men_men_n859_));
  NA2        u0831(.A(men_men_n747_), .B(men_men_n365_), .Y(men_men_n860_));
  OAI210     u0832(.A0(men_men_n623_), .A1(men_men_n622_), .B0(men_men_n380_), .Y(men_men_n861_));
  AN3        u0833(.A(men_men_n861_), .B(men_men_n860_), .C(men_men_n858_), .Y(men_men_n862_));
  NAi41      u0834(.An(men_men_n856_), .B(men_men_n862_), .C(men_men_n857_), .D(men_men_n851_), .Y(men_men_n863_));
  NO4        u0835(.A(men_men_n863_), .B(men_men_n849_), .C(men_men_n847_), .D(men_men_n841_), .Y(men_men_n864_));
  NA4        u0836(.A(men_men_n864_), .B(men_men_n834_), .C(men_men_n789_), .D(men_men_n774_), .Y(men09));
  INV        u0837(.A(men_men_n123_), .Y(men_men_n866_));
  NA2        u0838(.A(f), .B(e), .Y(men_men_n867_));
  NO2        u0839(.A(men_men_n234_), .B(men_men_n113_), .Y(men_men_n868_));
  NA2        u0840(.A(men_men_n868_), .B(g), .Y(men_men_n869_));
  NA4        u0841(.A(men_men_n326_), .B(men_men_n490_), .C(men_men_n272_), .D(men_men_n120_), .Y(men_men_n870_));
  AOI210     u0842(.A0(men_men_n870_), .A1(g), .B0(men_men_n487_), .Y(men_men_n871_));
  AOI210     u0843(.A0(men_men_n871_), .A1(men_men_n869_), .B0(men_men_n867_), .Y(men_men_n872_));
  NA2        u0844(.A(men_men_n872_), .B(men_men_n866_), .Y(men_men_n873_));
  NO2        u0845(.A(men_men_n211_), .B(men_men_n221_), .Y(men_men_n874_));
  NA3        u0846(.A(m), .B(l), .C(i), .Y(men_men_n875_));
  NA4        u0847(.A(men_men_n88_), .B(men_men_n87_), .C(g), .D(f), .Y(men_men_n876_));
  NA2        u0848(.A(men_men_n876_), .B(men_men_n457_), .Y(men_men_n877_));
  OA210      u0849(.A0(men_men_n877_), .A1(men_men_n874_), .B0(men_men_n591_), .Y(men_men_n878_));
  NA3        u0850(.A(men_men_n842_), .B(men_men_n593_), .C(men_men_n541_), .Y(men_men_n879_));
  OA210      u0851(.A0(men_men_n879_), .A1(men_men_n878_), .B0(men_men_n845_), .Y(men_men_n880_));
  INV        u0852(.A(men_men_n354_), .Y(men_men_n881_));
  NO2        u0853(.A(men_men_n129_), .B(men_men_n127_), .Y(men_men_n882_));
  NOi31      u0854(.An(k), .B(m), .C(l), .Y(men_men_n883_));
  NO2        u0855(.A(men_men_n356_), .B(men_men_n883_), .Y(men_men_n884_));
  AOI210     u0856(.A0(men_men_n884_), .A1(men_men_n882_), .B0(men_men_n626_), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n828_), .B(men_men_n347_), .Y(men_men_n886_));
  NA2        u0858(.A(men_men_n358_), .B(men_men_n360_), .Y(men_men_n887_));
  OAI210     u0859(.A0(men_men_n211_), .A1(men_men_n221_), .B0(men_men_n887_), .Y(men_men_n888_));
  AOI220     u0860(.A0(men_men_n888_), .A1(men_men_n886_), .B0(men_men_n885_), .B1(men_men_n881_), .Y(men_men_n889_));
  NA2        u0861(.A(men_men_n173_), .B(men_men_n115_), .Y(men_men_n890_));
  NA3        u0862(.A(men_men_n890_), .B(men_men_n731_), .C(men_men_n138_), .Y(men_men_n891_));
  NA3        u0863(.A(men_men_n891_), .B(men_men_n196_), .C(men_men_n31_), .Y(men_men_n892_));
  NA3        u0864(.A(men_men_n892_), .B(men_men_n889_), .C(men_men_n655_), .Y(men_men_n893_));
  NO2        u0865(.A(men_men_n613_), .B(men_men_n519_), .Y(men_men_n894_));
  NA2        u0866(.A(men_men_n894_), .B(men_men_n196_), .Y(men_men_n895_));
  NOi21      u0867(.An(f), .B(d), .Y(men_men_n896_));
  NA2        u0868(.A(men_men_n896_), .B(m), .Y(men_men_n897_));
  NO2        u0869(.A(men_men_n897_), .B(men_men_n52_), .Y(men_men_n898_));
  NOi32      u0870(.An(g), .Bn(f), .C(d), .Y(men_men_n899_));
  NA4        u0871(.A(men_men_n899_), .B(men_men_n633_), .C(men_men_n29_), .D(m), .Y(men_men_n900_));
  NOi21      u0872(.An(men_men_n327_), .B(men_men_n900_), .Y(men_men_n901_));
  AOI210     u0873(.A0(men_men_n898_), .A1(men_men_n568_), .B0(men_men_n901_), .Y(men_men_n902_));
  NA3        u0874(.A(men_men_n326_), .B(men_men_n272_), .C(men_men_n120_), .Y(men_men_n903_));
  AN2        u0875(.A(f), .B(d), .Y(men_men_n904_));
  NA3        u0876(.A(men_men_n495_), .B(men_men_n904_), .C(men_men_n84_), .Y(men_men_n905_));
  NO3        u0877(.A(men_men_n905_), .B(men_men_n75_), .C(men_men_n222_), .Y(men_men_n906_));
  NO2        u0878(.A(men_men_n299_), .B(men_men_n56_), .Y(men_men_n907_));
  OAI210     u0879(.A0(men_men_n907_), .A1(men_men_n903_), .B0(men_men_n906_), .Y(men_men_n908_));
  NAi41      u0880(.An(men_men_n509_), .B(men_men_n908_), .C(men_men_n902_), .D(men_men_n895_), .Y(men_men_n909_));
  NO4        u0881(.A(men_men_n653_), .B(men_men_n134_), .C(men_men_n343_), .D(men_men_n156_), .Y(men_men_n910_));
  NO2        u0882(.A(men_men_n685_), .B(men_men_n343_), .Y(men_men_n911_));
  AN2        u0883(.A(men_men_n911_), .B(men_men_n712_), .Y(men_men_n912_));
  NO3        u0884(.A(men_men_n912_), .B(men_men_n910_), .C(men_men_n243_), .Y(men_men_n913_));
  NA2        u0885(.A(men_men_n631_), .B(men_men_n84_), .Y(men_men_n914_));
  OAI220     u0886(.A0(men_men_n887_), .A1(men_men_n914_), .B0(men_men_n828_), .B1(men_men_n457_), .Y(men_men_n915_));
  NA3        u0887(.A(men_men_n164_), .B(men_men_n109_), .C(men_men_n108_), .Y(men_men_n916_));
  OAI220     u0888(.A0(men_men_n905_), .A1(men_men_n446_), .B0(men_men_n354_), .B1(men_men_n916_), .Y(men_men_n917_));
  NOi41      u0889(.An(men_men_n232_), .B(men_men_n917_), .C(men_men_n915_), .D(men_men_n321_), .Y(men_men_n918_));
  NA2        u0890(.A(c), .B(men_men_n117_), .Y(men_men_n919_));
  NO2        u0891(.A(men_men_n919_), .B(men_men_n426_), .Y(men_men_n920_));
  NA3        u0892(.A(men_men_n920_), .B(men_men_n531_), .C(f), .Y(men_men_n921_));
  OR2        u0893(.A(men_men_n692_), .B(men_men_n564_), .Y(men_men_n922_));
  INV        u0894(.A(men_men_n922_), .Y(men_men_n923_));
  NA2        u0895(.A(men_men_n844_), .B(men_men_n112_), .Y(men_men_n924_));
  NA2        u0896(.A(men_men_n924_), .B(men_men_n923_), .Y(men_men_n925_));
  NA4        u0897(.A(men_men_n925_), .B(men_men_n921_), .C(men_men_n918_), .D(men_men_n913_), .Y(men_men_n926_));
  NO4        u0898(.A(men_men_n926_), .B(men_men_n909_), .C(men_men_n893_), .D(men_men_n880_), .Y(men_men_n927_));
  OR2        u0899(.A(men_men_n905_), .B(men_men_n75_), .Y(men_men_n928_));
  NA2        u0900(.A(men_men_n113_), .B(j), .Y(men_men_n929_));
  NA2        u0901(.A(men_men_n868_), .B(g), .Y(men_men_n930_));
  AOI210     u0902(.A0(men_men_n930_), .A1(men_men_n307_), .B0(men_men_n928_), .Y(men_men_n931_));
  AOI210     u0903(.A0(men_men_n828_), .A1(men_men_n347_), .B0(men_men_n876_), .Y(men_men_n932_));
  NO2        u0904(.A(men_men_n138_), .B(men_men_n134_), .Y(men_men_n933_));
  NO2        u0905(.A(men_men_n239_), .B(men_men_n233_), .Y(men_men_n934_));
  AOI220     u0906(.A0(men_men_n934_), .A1(men_men_n236_), .B0(men_men_n320_), .B1(men_men_n933_), .Y(men_men_n935_));
  NO2        u0907(.A(men_men_n446_), .B(men_men_n867_), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n936_), .B(men_men_n585_), .Y(men_men_n937_));
  NA2        u0909(.A(men_men_n937_), .B(men_men_n935_), .Y(men_men_n938_));
  NA2        u0910(.A(e), .B(d), .Y(men_men_n939_));
  OAI220     u0911(.A0(men_men_n939_), .A1(c), .B0(men_men_n340_), .B1(d), .Y(men_men_n940_));
  NA3        u0912(.A(men_men_n940_), .B(men_men_n473_), .C(men_men_n529_), .Y(men_men_n941_));
  AOI210     u0913(.A0(men_men_n537_), .A1(men_men_n186_), .B0(men_men_n239_), .Y(men_men_n942_));
  AOI210     u0914(.A0(men_men_n654_), .A1(men_men_n363_), .B0(men_men_n942_), .Y(men_men_n943_));
  NA2        u0915(.A(men_men_n299_), .B(men_men_n169_), .Y(men_men_n944_));
  NA2        u0916(.A(men_men_n906_), .B(men_men_n944_), .Y(men_men_n945_));
  NA3        u0917(.A(men_men_n945_), .B(men_men_n943_), .C(men_men_n941_), .Y(men_men_n946_));
  NO4        u0918(.A(men_men_n946_), .B(men_men_n938_), .C(men_men_n932_), .D(men_men_n931_), .Y(men_men_n947_));
  NA2        u0919(.A(men_men_n881_), .B(men_men_n31_), .Y(men_men_n948_));
  AO210      u0920(.A0(men_men_n948_), .A1(men_men_n733_), .B0(men_men_n225_), .Y(men_men_n949_));
  OAI220     u0921(.A0(men_men_n653_), .A1(men_men_n61_), .B0(men_men_n315_), .B1(j), .Y(men_men_n950_));
  AOI220     u0922(.A0(men_men_n950_), .A1(men_men_n911_), .B0(men_men_n643_), .B1(men_men_n652_), .Y(men_men_n951_));
  INV        u0923(.A(men_men_n951_), .Y(men_men_n952_));
  OAI210     u0924(.A0(men_men_n868_), .A1(men_men_n944_), .B0(men_men_n899_), .Y(men_men_n953_));
  NO2        u0925(.A(men_men_n953_), .B(men_men_n634_), .Y(men_men_n954_));
  AOI210     u0926(.A0(men_men_n119_), .A1(men_men_n118_), .B0(men_men_n271_), .Y(men_men_n955_));
  NO2        u0927(.A(men_men_n955_), .B(men_men_n900_), .Y(men_men_n956_));
  NOi31      u0928(.An(men_men_n568_), .B(men_men_n897_), .C(men_men_n307_), .Y(men_men_n957_));
  NO4        u0929(.A(men_men_n957_), .B(men_men_n956_), .C(men_men_n954_), .D(men_men_n952_), .Y(men_men_n958_));
  AO220      u0930(.A0(men_men_n473_), .A1(men_men_n784_), .B0(men_men_n181_), .B1(f), .Y(men_men_n959_));
  OAI210     u0931(.A0(men_men_n959_), .A1(men_men_n476_), .B0(men_men_n940_), .Y(men_men_n960_));
  NO2        u0932(.A(men_men_n456_), .B(men_men_n71_), .Y(men_men_n961_));
  OAI210     u0933(.A0(men_men_n879_), .A1(men_men_n961_), .B0(men_men_n737_), .Y(men_men_n962_));
  AN4        u0934(.A(men_men_n962_), .B(men_men_n960_), .C(men_men_n958_), .D(men_men_n949_), .Y(men_men_n963_));
  NA4        u0935(.A(men_men_n963_), .B(men_men_n947_), .C(men_men_n927_), .D(men_men_n873_), .Y(men12));
  NO2        u0936(.A(men_men_n471_), .B(c), .Y(men_men_n965_));
  NO4        u0937(.A(men_men_n461_), .B(men_men_n263_), .C(men_men_n609_), .D(men_men_n222_), .Y(men_men_n966_));
  NA2        u0938(.A(men_men_n966_), .B(men_men_n965_), .Y(men_men_n967_));
  NA2        u0939(.A(men_men_n568_), .B(men_men_n961_), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n471_), .B(men_men_n117_), .Y(men_men_n969_));
  NO2        u0941(.A(men_men_n882_), .B(men_men_n370_), .Y(men_men_n970_));
  NO2        u0942(.A(men_men_n692_), .B(men_men_n395_), .Y(men_men_n971_));
  AOI220     u0943(.A0(men_men_n971_), .A1(men_men_n566_), .B0(men_men_n970_), .B1(men_men_n969_), .Y(men_men_n972_));
  NA4        u0944(.A(men_men_n972_), .B(men_men_n968_), .C(men_men_n967_), .D(men_men_n460_), .Y(men_men_n973_));
  AOI210     u0945(.A0(men_men_n242_), .A1(men_men_n353_), .B0(men_men_n208_), .Y(men_men_n974_));
  OR2        u0946(.A(men_men_n974_), .B(men_men_n966_), .Y(men_men_n975_));
  AOI210     u0947(.A0(men_men_n350_), .A1(men_men_n407_), .B0(men_men_n222_), .Y(men_men_n976_));
  OAI210     u0948(.A0(men_men_n976_), .A1(men_men_n975_), .B0(men_men_n421_), .Y(men_men_n977_));
  NO2        u0949(.A(men_men_n673_), .B(men_men_n274_), .Y(men_men_n978_));
  NO2        u0950(.A(men_men_n617_), .B(men_men_n875_), .Y(men_men_n979_));
  AOI220     u0951(.A0(men_men_n979_), .A1(men_men_n591_), .B0(men_men_n852_), .B1(men_men_n978_), .Y(men_men_n980_));
  NO2        u0952(.A(men_men_n155_), .B(men_men_n246_), .Y(men_men_n981_));
  NA3        u0953(.A(men_men_n981_), .B(men_men_n249_), .C(i), .Y(men_men_n982_));
  NA3        u0954(.A(men_men_n982_), .B(men_men_n980_), .C(men_men_n977_), .Y(men_men_n983_));
  OR2        u0955(.A(men_men_n341_), .B(men_men_n969_), .Y(men_men_n984_));
  NA2        u0956(.A(men_men_n984_), .B(men_men_n371_), .Y(men_men_n985_));
  NO3        u0957(.A(men_men_n134_), .B(men_men_n156_), .C(men_men_n222_), .Y(men_men_n986_));
  NA2        u0958(.A(men_men_n986_), .B(men_men_n553_), .Y(men_men_n987_));
  NA2        u0959(.A(men_men_n987_), .B(men_men_n985_), .Y(men_men_n988_));
  NO3        u0960(.A(men_men_n697_), .B(men_men_n92_), .C(men_men_n45_), .Y(men_men_n989_));
  NO4        u0961(.A(men_men_n989_), .B(men_men_n988_), .C(men_men_n983_), .D(men_men_n973_), .Y(men_men_n990_));
  NO2        u0962(.A(men_men_n385_), .B(men_men_n384_), .Y(men_men_n991_));
  NA2        u0963(.A(men_men_n614_), .B(men_men_n73_), .Y(men_men_n992_));
  NA2        u0964(.A(men_men_n578_), .B(men_men_n148_), .Y(men_men_n993_));
  NOi21      u0965(.An(men_men_n34_), .B(men_men_n685_), .Y(men_men_n994_));
  AOI220     u0966(.A0(men_men_n994_), .A1(men_men_n993_), .B0(men_men_n992_), .B1(men_men_n991_), .Y(men_men_n995_));
  OAI210     u0967(.A0(men_men_n261_), .A1(men_men_n45_), .B0(men_men_n995_), .Y(men_men_n996_));
  NA2        u0968(.A(men_men_n452_), .B(men_men_n276_), .Y(men_men_n997_));
  NO3        u0969(.A(men_men_n854_), .B(men_men_n89_), .C(men_men_n426_), .Y(men_men_n998_));
  NAi31      u0970(.An(men_men_n998_), .B(men_men_n997_), .C(men_men_n337_), .Y(men_men_n999_));
  NO2        u0971(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n1000_));
  NO2        u0972(.A(men_men_n526_), .B(men_men_n315_), .Y(men_men_n1001_));
  NA2        u0973(.A(men_men_n664_), .B(men_men_n380_), .Y(men_men_n1002_));
  OAI210     u0974(.A0(men_men_n770_), .A1(men_men_n1002_), .B0(men_men_n382_), .Y(men_men_n1003_));
  NO3        u0975(.A(men_men_n1003_), .B(men_men_n999_), .C(men_men_n996_), .Y(men_men_n1004_));
  NA2        u0976(.A(men_men_n363_), .B(g), .Y(men_men_n1005_));
  NA2        u0977(.A(men_men_n166_), .B(i), .Y(men_men_n1006_));
  NA2        u0978(.A(men_men_n46_), .B(i), .Y(men_men_n1007_));
  NO2        u0979(.A(men_men_n148_), .B(men_men_n84_), .Y(men_men_n1008_));
  OR2        u0980(.A(men_men_n1008_), .B(men_men_n577_), .Y(men_men_n1009_));
  NA2        u0981(.A(men_men_n578_), .B(men_men_n399_), .Y(men_men_n1010_));
  AOI210     u0982(.A0(men_men_n1010_), .A1(n), .B0(men_men_n1009_), .Y(men_men_n1011_));
  NO2        u0983(.A(men_men_n1011_), .B(men_men_n1005_), .Y(men_men_n1012_));
  NO2        u0984(.A(men_men_n692_), .B(men_men_n519_), .Y(men_men_n1013_));
  NA3        u0985(.A(men_men_n358_), .B(men_men_n659_), .C(i), .Y(men_men_n1014_));
  OAI210     u0986(.A0(men_men_n456_), .A1(men_men_n326_), .B0(men_men_n1014_), .Y(men_men_n1015_));
  OAI220     u0987(.A0(men_men_n1015_), .A1(men_men_n1013_), .B0(men_men_n709_), .B1(men_men_n796_), .Y(men_men_n1016_));
  NA2        u0988(.A(men_men_n637_), .B(men_men_n114_), .Y(men_men_n1017_));
  OR3        u0989(.A(men_men_n326_), .B(men_men_n451_), .C(f), .Y(men_men_n1018_));
  NA3        u0990(.A(men_men_n659_), .B(men_men_n82_), .C(i), .Y(men_men_n1019_));
  OA220      u0991(.A0(men_men_n1019_), .A1(men_men_n1017_), .B0(men_men_n1018_), .B1(men_men_n616_), .Y(men_men_n1020_));
  NA3        u0992(.A(men_men_n342_), .B(men_men_n119_), .C(g), .Y(men_men_n1021_));
  AOI210     u0993(.A0(men_men_n707_), .A1(men_men_n1021_), .B0(m), .Y(men_men_n1022_));
  OAI210     u0994(.A0(men_men_n1022_), .A1(men_men_n970_), .B0(men_men_n341_), .Y(men_men_n1023_));
  NA2        u0995(.A(men_men_n724_), .B(men_men_n914_), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n876_), .B(men_men_n457_), .Y(men_men_n1025_));
  NA2        u0997(.A(men_men_n230_), .B(men_men_n79_), .Y(men_men_n1026_));
  NA3        u0998(.A(men_men_n1026_), .B(men_men_n1019_), .C(men_men_n1018_), .Y(men_men_n1027_));
  AOI220     u0999(.A0(men_men_n1027_), .A1(men_men_n269_), .B0(men_men_n1025_), .B1(men_men_n1024_), .Y(men_men_n1028_));
  NA4        u1000(.A(men_men_n1028_), .B(men_men_n1023_), .C(men_men_n1020_), .D(men_men_n1016_), .Y(men_men_n1029_));
  NO2        u1001(.A(men_men_n395_), .B(men_men_n91_), .Y(men_men_n1030_));
  OAI210     u1002(.A0(men_men_n1030_), .A1(men_men_n978_), .B0(men_men_n247_), .Y(men_men_n1031_));
  NA2        u1003(.A(men_men_n696_), .B(men_men_n88_), .Y(men_men_n1032_));
  NO2        u1004(.A(men_men_n479_), .B(men_men_n222_), .Y(men_men_n1033_));
  AOI220     u1005(.A0(men_men_n1033_), .A1(men_men_n400_), .B0(men_men_n984_), .B1(men_men_n226_), .Y(men_men_n1034_));
  AOI220     u1006(.A0(men_men_n971_), .A1(men_men_n981_), .B0(men_men_n615_), .B1(men_men_n90_), .Y(men_men_n1035_));
  NA4        u1007(.A(men_men_n1035_), .B(men_men_n1034_), .C(men_men_n1032_), .D(men_men_n1031_), .Y(men_men_n1036_));
  OAI210     u1008(.A0(men_men_n1025_), .A1(men_men_n979_), .B0(men_men_n566_), .Y(men_men_n1037_));
  AOI210     u1009(.A0(men_men_n437_), .A1(men_men_n430_), .B0(men_men_n854_), .Y(men_men_n1038_));
  OAI210     u1010(.A0(men_men_n385_), .A1(men_men_n384_), .B0(men_men_n110_), .Y(men_men_n1039_));
  AOI210     u1011(.A0(men_men_n1039_), .A1(men_men_n558_), .B0(men_men_n1038_), .Y(men_men_n1040_));
  NA2        u1012(.A(men_men_n1022_), .B(men_men_n969_), .Y(men_men_n1041_));
  NO3        u1013(.A(men_men_n929_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1042_));
  NA2        u1014(.A(men_men_n1042_), .B(men_men_n657_), .Y(men_men_n1043_));
  NA4        u1015(.A(men_men_n1043_), .B(men_men_n1041_), .C(men_men_n1040_), .D(men_men_n1037_), .Y(men_men_n1044_));
  NO4        u1016(.A(men_men_n1044_), .B(men_men_n1036_), .C(men_men_n1029_), .D(men_men_n1012_), .Y(men_men_n1045_));
  NAi31      u1017(.An(men_men_n144_), .B(men_men_n438_), .C(n), .Y(men_men_n1046_));
  NO3        u1018(.A(men_men_n127_), .B(men_men_n356_), .C(men_men_n883_), .Y(men_men_n1047_));
  NO2        u1019(.A(men_men_n1047_), .B(men_men_n1046_), .Y(men_men_n1048_));
  NO3        u1020(.A(men_men_n284_), .B(men_men_n144_), .C(men_men_n426_), .Y(men_men_n1049_));
  AOI210     u1021(.A0(men_men_n1049_), .A1(men_men_n520_), .B0(men_men_n1048_), .Y(men_men_n1050_));
  NA2        u1022(.A(men_men_n512_), .B(i), .Y(men_men_n1051_));
  NA2        u1023(.A(men_men_n1051_), .B(men_men_n1050_), .Y(men_men_n1052_));
  NA2        u1024(.A(men_men_n239_), .B(men_men_n177_), .Y(men_men_n1053_));
  NO3        u1025(.A(men_men_n323_), .B(men_men_n462_), .C(men_men_n181_), .Y(men_men_n1054_));
  NOi31      u1026(.An(men_men_n1053_), .B(men_men_n1054_), .C(men_men_n222_), .Y(men_men_n1055_));
  NA2        u1027(.A(men_men_n455_), .B(men_men_n914_), .Y(men_men_n1056_));
  NO3        u1028(.A(men_men_n456_), .B(men_men_n326_), .C(men_men_n75_), .Y(men_men_n1057_));
  AOI220     u1029(.A0(men_men_n1057_), .A1(men_men_n1056_), .B0(men_men_n501_), .B1(g), .Y(men_men_n1058_));
  INV        u1030(.A(men_men_n1058_), .Y(men_men_n1059_));
  OAI220     u1031(.A0(men_men_n1046_), .A1(men_men_n242_), .B0(men_men_n1014_), .B1(men_men_n632_), .Y(men_men_n1060_));
  NO2        u1032(.A(men_men_n693_), .B(men_men_n395_), .Y(men_men_n1061_));
  NA2        u1033(.A(men_men_n974_), .B(men_men_n965_), .Y(men_men_n1062_));
  NO3        u1034(.A(men_men_n567_), .B(men_men_n153_), .C(men_men_n221_), .Y(men_men_n1063_));
  OAI210     u1035(.A0(men_men_n1063_), .A1(men_men_n547_), .B0(men_men_n396_), .Y(men_men_n1064_));
  OAI220     u1036(.A0(men_men_n971_), .A1(men_men_n979_), .B0(men_men_n568_), .B1(men_men_n445_), .Y(men_men_n1065_));
  NA4        u1037(.A(men_men_n1065_), .B(men_men_n1064_), .C(men_men_n1062_), .D(men_men_n651_), .Y(men_men_n1066_));
  OAI210     u1038(.A0(men_men_n974_), .A1(men_men_n966_), .B0(men_men_n1053_), .Y(men_men_n1067_));
  NA3        u1039(.A(men_men_n1010_), .B(men_men_n506_), .C(men_men_n46_), .Y(men_men_n1068_));
  AOI210     u1040(.A0(men_men_n398_), .A1(men_men_n396_), .B0(men_men_n346_), .Y(men_men_n1069_));
  NA4        u1041(.A(men_men_n1069_), .B(men_men_n1068_), .C(men_men_n1067_), .D(men_men_n285_), .Y(men_men_n1070_));
  OR4        u1042(.A(men_men_n1070_), .B(men_men_n1066_), .C(men_men_n1061_), .D(men_men_n1060_), .Y(men_men_n1071_));
  NO4        u1043(.A(men_men_n1071_), .B(men_men_n1059_), .C(men_men_n1055_), .D(men_men_n1052_), .Y(men_men_n1072_));
  NA4        u1044(.A(men_men_n1072_), .B(men_men_n1045_), .C(men_men_n1004_), .D(men_men_n990_), .Y(men13));
  NA2        u1045(.A(men_men_n46_), .B(men_men_n87_), .Y(men_men_n1074_));
  AN2        u1046(.A(c), .B(b), .Y(men_men_n1075_));
  NA3        u1047(.A(men_men_n260_), .B(men_men_n1075_), .C(m), .Y(men_men_n1076_));
  NA2        u1048(.A(men_men_n517_), .B(f), .Y(men_men_n1077_));
  NO4        u1049(.A(men_men_n1077_), .B(men_men_n1076_), .C(men_men_n1074_), .D(men_men_n610_), .Y(men_men_n1078_));
  NA2        u1050(.A(men_men_n276_), .B(men_men_n1075_), .Y(men_men_n1079_));
  NO4        u1051(.A(men_men_n1079_), .B(men_men_n1077_), .C(men_men_n1006_), .D(a), .Y(men_men_n1080_));
  NAi32      u1052(.An(d), .Bn(c), .C(e), .Y(men_men_n1081_));
  NA2        u1053(.A(men_men_n143_), .B(men_men_n45_), .Y(men_men_n1082_));
  NO4        u1054(.A(men_men_n1082_), .B(men_men_n1081_), .C(men_men_n617_), .D(men_men_n322_), .Y(men_men_n1083_));
  NA2        u1055(.A(men_men_n700_), .B(men_men_n233_), .Y(men_men_n1084_));
  NA2        u1056(.A(men_men_n429_), .B(men_men_n221_), .Y(men_men_n1085_));
  AN2        u1057(.A(d), .B(c), .Y(men_men_n1086_));
  NA2        u1058(.A(men_men_n1086_), .B(men_men_n117_), .Y(men_men_n1087_));
  NO4        u1059(.A(men_men_n1087_), .B(men_men_n1085_), .C(men_men_n182_), .D(men_men_n173_), .Y(men_men_n1088_));
  NA2        u1060(.A(men_men_n517_), .B(c), .Y(men_men_n1089_));
  NO4        u1061(.A(men_men_n1082_), .B(men_men_n613_), .C(men_men_n1089_), .D(men_men_n322_), .Y(men_men_n1090_));
  AO210      u1062(.A0(men_men_n1088_), .A1(men_men_n1084_), .B0(men_men_n1090_), .Y(men_men_n1091_));
  OR4        u1063(.A(men_men_n1091_), .B(men_men_n1083_), .C(men_men_n1080_), .D(men_men_n1078_), .Y(men_men_n1092_));
  NAi32      u1064(.An(f), .Bn(e), .C(c), .Y(men_men_n1093_));
  NO2        u1065(.A(men_men_n1093_), .B(men_men_n150_), .Y(men_men_n1094_));
  NA2        u1066(.A(men_men_n1094_), .B(g), .Y(men_men_n1095_));
  OR3        u1067(.A(men_men_n233_), .B(men_men_n182_), .C(men_men_n173_), .Y(men_men_n1096_));
  NO2        u1068(.A(men_men_n1096_), .B(men_men_n1095_), .Y(men_men_n1097_));
  NO2        u1069(.A(men_men_n1089_), .B(men_men_n322_), .Y(men_men_n1098_));
  NO2        u1070(.A(j), .B(men_men_n45_), .Y(men_men_n1099_));
  NA2        u1071(.A(men_men_n661_), .B(men_men_n1099_), .Y(men_men_n1100_));
  NOi21      u1072(.An(men_men_n1098_), .B(men_men_n1100_), .Y(men_men_n1101_));
  NO2        u1073(.A(men_men_n800_), .B(men_men_n113_), .Y(men_men_n1102_));
  NOi41      u1074(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1103_));
  NA2        u1075(.A(men_men_n1103_), .B(men_men_n1102_), .Y(men_men_n1104_));
  NO2        u1076(.A(men_men_n1104_), .B(men_men_n1095_), .Y(men_men_n1105_));
  OR3        u1077(.A(e), .B(d), .C(c), .Y(men_men_n1106_));
  NA3        u1078(.A(k), .B(j), .C(i), .Y(men_men_n1107_));
  NO3        u1079(.A(men_men_n1107_), .B(men_men_n322_), .C(men_men_n91_), .Y(men_men_n1108_));
  NOi21      u1080(.An(men_men_n1108_), .B(men_men_n1106_), .Y(men_men_n1109_));
  OR4        u1081(.A(men_men_n1109_), .B(men_men_n1105_), .C(men_men_n1101_), .D(men_men_n1097_), .Y(men_men_n1110_));
  NA3        u1082(.A(men_men_n485_), .B(men_men_n349_), .C(men_men_n56_), .Y(men_men_n1111_));
  NO2        u1083(.A(men_men_n1111_), .B(men_men_n1100_), .Y(men_men_n1112_));
  NO4        u1084(.A(men_men_n1111_), .B(men_men_n613_), .C(men_men_n469_), .D(men_men_n45_), .Y(men_men_n1113_));
  NO2        u1085(.A(f), .B(c), .Y(men_men_n1114_));
  NOi21      u1086(.An(men_men_n1114_), .B(men_men_n461_), .Y(men_men_n1115_));
  NA2        u1087(.A(men_men_n1115_), .B(men_men_n59_), .Y(men_men_n1116_));
  OR2        u1088(.A(k), .B(i), .Y(men_men_n1117_));
  NO3        u1089(.A(men_men_n1117_), .B(men_men_n253_), .C(l), .Y(men_men_n1118_));
  NOi31      u1090(.An(men_men_n1118_), .B(men_men_n1116_), .C(j), .Y(men_men_n1119_));
  OR3        u1091(.A(men_men_n1119_), .B(men_men_n1113_), .C(men_men_n1112_), .Y(men_men_n1120_));
  OR3        u1092(.A(men_men_n1120_), .B(men_men_n1110_), .C(men_men_n1092_), .Y(men02));
  OR2        u1093(.A(l), .B(k), .Y(men_men_n1122_));
  OR3        u1094(.A(h), .B(g), .C(f), .Y(men_men_n1123_));
  OR3        u1095(.A(n), .B(m), .C(i), .Y(men_men_n1124_));
  NO4        u1096(.A(men_men_n1124_), .B(men_men_n1123_), .C(men_men_n1122_), .D(men_men_n1106_), .Y(men_men_n1125_));
  NOi31      u1097(.An(e), .B(d), .C(c), .Y(men_men_n1126_));
  AOI210     u1098(.A0(men_men_n1108_), .A1(men_men_n1126_), .B0(men_men_n1083_), .Y(men_men_n1127_));
  AN3        u1099(.A(g), .B(f), .C(c), .Y(men_men_n1128_));
  NA3        u1100(.A(men_men_n1128_), .B(men_men_n485_), .C(h), .Y(men_men_n1129_));
  OR2        u1101(.A(men_men_n1107_), .B(men_men_n322_), .Y(men_men_n1130_));
  OR2        u1102(.A(men_men_n1130_), .B(men_men_n1129_), .Y(men_men_n1131_));
  NO3        u1103(.A(men_men_n1111_), .B(men_men_n1082_), .C(men_men_n613_), .Y(men_men_n1132_));
  NO2        u1104(.A(men_men_n1132_), .B(men_men_n1097_), .Y(men_men_n1133_));
  NA3        u1105(.A(l), .B(k), .C(j), .Y(men_men_n1134_));
  NA2        u1106(.A(i), .B(h), .Y(men_men_n1135_));
  NO3        u1107(.A(men_men_n1135_), .B(men_men_n1134_), .C(men_men_n134_), .Y(men_men_n1136_));
  NO3        u1108(.A(men_men_n145_), .B(men_men_n297_), .C(men_men_n222_), .Y(men_men_n1137_));
  AOI210     u1109(.A0(men_men_n1137_), .A1(men_men_n1136_), .B0(men_men_n1101_), .Y(men_men_n1138_));
  NA3        u1110(.A(c), .B(b), .C(a), .Y(men_men_n1139_));
  NO3        u1111(.A(men_men_n1139_), .B(men_men_n939_), .C(men_men_n221_), .Y(men_men_n1140_));
  NO4        u1112(.A(men_men_n1107_), .B(men_men_n315_), .C(men_men_n49_), .D(men_men_n113_), .Y(men_men_n1141_));
  AOI210     u1113(.A0(men_men_n1141_), .A1(men_men_n1140_), .B0(men_men_n1112_), .Y(men_men_n1142_));
  AN4        u1114(.A(men_men_n1142_), .B(men_men_n1138_), .C(men_men_n1133_), .D(men_men_n1131_), .Y(men_men_n1143_));
  NO2        u1115(.A(men_men_n1087_), .B(men_men_n1085_), .Y(men_men_n1144_));
  NA2        u1116(.A(men_men_n1104_), .B(men_men_n1096_), .Y(men_men_n1145_));
  AOI210     u1117(.A0(men_men_n1145_), .A1(men_men_n1144_), .B0(men_men_n1078_), .Y(men_men_n1146_));
  NAi41      u1118(.An(men_men_n1125_), .B(men_men_n1146_), .C(men_men_n1143_), .D(men_men_n1127_), .Y(men03));
  NO2        u1119(.A(men_men_n549_), .B(men_men_n626_), .Y(men_men_n1148_));
  NA4        u1120(.A(men_men_n88_), .B(men_men_n87_), .C(g), .D(men_men_n221_), .Y(men_men_n1149_));
  NA4        u1121(.A(men_men_n601_), .B(m), .C(men_men_n113_), .D(men_men_n221_), .Y(men_men_n1150_));
  NA3        u1122(.A(men_men_n1150_), .B(men_men_n386_), .C(men_men_n1149_), .Y(men_men_n1151_));
  NO3        u1123(.A(men_men_n1151_), .B(men_men_n1148_), .C(men_men_n1039_), .Y(men_men_n1152_));
  NOi41      u1124(.An(men_men_n842_), .B(men_men_n888_), .C(men_men_n877_), .D(men_men_n749_), .Y(men_men_n1153_));
  OAI220     u1125(.A0(men_men_n1153_), .A1(men_men_n724_), .B0(men_men_n1152_), .B1(men_men_n614_), .Y(men_men_n1154_));
  NA4        u1126(.A(i), .B(men_men_n1126_), .C(men_men_n358_), .D(men_men_n349_), .Y(men_men_n1155_));
  OAI210     u1127(.A0(men_men_n854_), .A1(men_men_n439_), .B0(men_men_n1155_), .Y(men_men_n1156_));
  NOi31      u1128(.An(m), .B(n), .C(f), .Y(men_men_n1157_));
  NA2        u1129(.A(men_men_n1157_), .B(men_men_n51_), .Y(men_men_n1158_));
  AN2        u1130(.A(e), .B(c), .Y(men_men_n1159_));
  NO2        u1131(.A(men_men_n922_), .B(men_men_n444_), .Y(men_men_n1160_));
  NA2        u1132(.A(men_men_n529_), .B(l), .Y(men_men_n1161_));
  NOi31      u1133(.An(men_men_n899_), .B(men_men_n1076_), .C(men_men_n1161_), .Y(men_men_n1162_));
  NO4        u1134(.A(men_men_n1162_), .B(men_men_n1160_), .C(men_men_n1156_), .D(men_men_n1038_), .Y(men_men_n1163_));
  NO2        u1135(.A(men_men_n297_), .B(a), .Y(men_men_n1164_));
  INV        u1136(.A(men_men_n1083_), .Y(men_men_n1165_));
  NO2        u1137(.A(men_men_n1135_), .B(men_men_n504_), .Y(men_men_n1166_));
  NO2        u1138(.A(men_men_n87_), .B(g), .Y(men_men_n1167_));
  AOI210     u1139(.A0(men_men_n1167_), .A1(men_men_n1166_), .B0(men_men_n1118_), .Y(men_men_n1168_));
  OR2        u1140(.A(men_men_n1168_), .B(men_men_n1116_), .Y(men_men_n1169_));
  NA3        u1141(.A(men_men_n1169_), .B(men_men_n1165_), .C(men_men_n1163_), .Y(men_men_n1170_));
  NO4        u1142(.A(men_men_n1170_), .B(men_men_n1154_), .C(men_men_n856_), .D(men_men_n590_), .Y(men_men_n1171_));
  NA2        u1143(.A(c), .B(b), .Y(men_men_n1172_));
  NO2        u1144(.A(men_men_n736_), .B(men_men_n1172_), .Y(men_men_n1173_));
  OAI210     u1145(.A0(men_men_n897_), .A1(men_men_n871_), .B0(men_men_n432_), .Y(men_men_n1174_));
  OAI210     u1146(.A0(men_men_n1174_), .A1(men_men_n898_), .B0(men_men_n1173_), .Y(men_men_n1175_));
  NA3        u1147(.A(men_men_n445_), .B(men_men_n583_), .C(f), .Y(men_men_n1176_));
  OAI210     u1148(.A0(men_men_n572_), .A1(men_men_n39_), .B0(men_men_n1164_), .Y(men_men_n1177_));
  NA2        u1149(.A(men_men_n1177_), .B(men_men_n1176_), .Y(men_men_n1178_));
  OAI210     u1150(.A0(k), .A1(men_men_n301_), .B0(g), .Y(men_men_n1179_));
  NAi21      u1151(.An(f), .B(d), .Y(men_men_n1180_));
  NO2        u1152(.A(men_men_n1180_), .B(men_men_n1139_), .Y(men_men_n1181_));
  INV        u1153(.A(men_men_n1181_), .Y(men_men_n1182_));
  AOI210     u1154(.A0(men_men_n1179_), .A1(men_men_n307_), .B0(men_men_n1182_), .Y(men_men_n1183_));
  AOI210     u1155(.A0(men_men_n1183_), .A1(men_men_n114_), .B0(men_men_n1178_), .Y(men_men_n1184_));
  NA2        u1156(.A(men_men_n487_), .B(men_men_n486_), .Y(men_men_n1185_));
  NO2        u1157(.A(men_men_n188_), .B(men_men_n246_), .Y(men_men_n1186_));
  NA2        u1158(.A(men_men_n1186_), .B(m), .Y(men_men_n1187_));
  NA3        u1159(.A(men_men_n955_), .B(men_men_n1161_), .C(men_men_n490_), .Y(men_men_n1188_));
  OAI210     u1160(.A0(men_men_n1188_), .A1(men_men_n327_), .B0(men_men_n488_), .Y(men_men_n1189_));
  AOI210     u1161(.A0(men_men_n1189_), .A1(men_men_n1185_), .B0(men_men_n1187_), .Y(men_men_n1190_));
  NA2        u1162(.A(men_men_n585_), .B(men_men_n428_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n163_), .B(men_men_n33_), .Y(men_men_n1192_));
  AOI210     u1164(.A0(men_men_n1002_), .A1(men_men_n1192_), .B0(men_men_n222_), .Y(men_men_n1193_));
  OAI210     u1165(.A0(men_men_n1193_), .A1(men_men_n465_), .B0(men_men_n1181_), .Y(men_men_n1194_));
  NO2        u1166(.A(men_men_n389_), .B(men_men_n388_), .Y(men_men_n1195_));
  AOI210     u1167(.A0(men_men_n1186_), .A1(men_men_n447_), .B0(men_men_n998_), .Y(men_men_n1196_));
  NAi41      u1168(.An(men_men_n1195_), .B(men_men_n1196_), .C(men_men_n1194_), .D(men_men_n1191_), .Y(men_men_n1197_));
  NO2        u1169(.A(men_men_n1197_), .B(men_men_n1190_), .Y(men_men_n1198_));
  NA4        u1170(.A(men_men_n1198_), .B(men_men_n1184_), .C(men_men_n1175_), .D(men_men_n1171_), .Y(men00));
  AOI210     u1171(.A0(men_men_n314_), .A1(men_men_n222_), .B0(men_men_n289_), .Y(men_men_n1200_));
  NO2        u1172(.A(men_men_n1200_), .B(men_men_n604_), .Y(men_men_n1201_));
  AOI210     u1173(.A0(men_men_n936_), .A1(men_men_n981_), .B0(men_men_n1156_), .Y(men_men_n1202_));
  NO3        u1174(.A(men_men_n1132_), .B(men_men_n998_), .C(men_men_n746_), .Y(men_men_n1203_));
  NA3        u1175(.A(men_men_n1203_), .B(men_men_n1202_), .C(men_men_n1040_), .Y(men_men_n1204_));
  NA2        u1176(.A(men_men_n531_), .B(f), .Y(men_men_n1205_));
  OAI210     u1177(.A0(men_men_n1047_), .A1(men_men_n40_), .B0(men_men_n678_), .Y(men_men_n1206_));
  NA3        u1178(.A(men_men_n1206_), .B(men_men_n268_), .C(n), .Y(men_men_n1207_));
  AOI210     u1179(.A0(men_men_n1207_), .A1(men_men_n1205_), .B0(men_men_n1087_), .Y(men_men_n1208_));
  NO4        u1180(.A(men_men_n1208_), .B(men_men_n1204_), .C(men_men_n1201_), .D(men_men_n1110_), .Y(men_men_n1209_));
  NA3        u1181(.A(men_men_n172_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1210_));
  NA3        u1182(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1211_));
  NOi31      u1183(.An(n), .B(m), .C(i), .Y(men_men_n1212_));
  NA3        u1184(.A(men_men_n1212_), .B(men_men_n681_), .C(men_men_n51_), .Y(men_men_n1213_));
  OAI210     u1185(.A0(men_men_n1211_), .A1(men_men_n1210_), .B0(men_men_n1213_), .Y(men_men_n1214_));
  INV        u1186(.A(men_men_n603_), .Y(men_men_n1215_));
  NO4        u1187(.A(men_men_n1215_), .B(men_men_n1214_), .C(men_men_n1195_), .D(men_men_n957_), .Y(men_men_n1216_));
  NO4        u1188(.A(men_men_n507_), .B(men_men_n373_), .C(men_men_n1172_), .D(men_men_n59_), .Y(men_men_n1217_));
  NA3        u1189(.A(men_men_n401_), .B(men_men_n229_), .C(g), .Y(men_men_n1218_));
  OA220      u1190(.A0(men_men_n1218_), .A1(men_men_n1211_), .B0(men_men_n402_), .B1(men_men_n137_), .Y(men_men_n1219_));
  NO2        u1191(.A(h), .B(g), .Y(men_men_n1220_));
  OAI220     u1192(.A0(men_men_n549_), .A1(men_men_n626_), .B0(men_men_n92_), .B1(men_men_n91_), .Y(men_men_n1221_));
  AOI220     u1193(.A0(men_men_n1221_), .A1(men_men_n558_), .B0(men_men_n986_), .B1(men_men_n602_), .Y(men_men_n1222_));
  AOI220     u1194(.A0(men_men_n334_), .A1(men_men_n257_), .B0(men_men_n183_), .B1(men_men_n152_), .Y(men_men_n1223_));
  NA3        u1195(.A(men_men_n1223_), .B(men_men_n1222_), .C(men_men_n1219_), .Y(men_men_n1224_));
  NO3        u1196(.A(men_men_n1224_), .B(men_men_n1217_), .C(men_men_n278_), .Y(men_men_n1225_));
  INV        u1197(.A(men_men_n339_), .Y(men_men_n1226_));
  AOI210     u1198(.A0(men_men_n257_), .A1(men_men_n363_), .B0(men_men_n605_), .Y(men_men_n1227_));
  NA3        u1199(.A(men_men_n1227_), .B(men_men_n1226_), .C(men_men_n158_), .Y(men_men_n1228_));
  NA3        u1200(.A(men_men_n185_), .B(men_men_n113_), .C(g), .Y(men_men_n1229_));
  NA3        u1201(.A(men_men_n485_), .B(men_men_n40_), .C(f), .Y(men_men_n1230_));
  NOi31      u1202(.An(men_men_n907_), .B(men_men_n1230_), .C(men_men_n1229_), .Y(men_men_n1231_));
  NAi31      u1203(.An(men_men_n192_), .B(men_men_n894_), .C(men_men_n485_), .Y(men_men_n1232_));
  NAi21      u1204(.An(men_men_n1231_), .B(men_men_n1232_), .Y(men_men_n1233_));
  NO2        u1205(.A(men_men_n288_), .B(men_men_n75_), .Y(men_men_n1234_));
  NO3        u1206(.A(men_men_n444_), .B(men_men_n867_), .C(n), .Y(men_men_n1235_));
  AOI210     u1207(.A0(men_men_n1235_), .A1(men_men_n1234_), .B0(men_men_n1125_), .Y(men_men_n1236_));
  NAi31      u1208(.An(men_men_n1090_), .B(men_men_n1236_), .C(men_men_n74_), .Y(men_men_n1237_));
  NO4        u1209(.A(men_men_n1237_), .B(men_men_n1233_), .C(men_men_n1228_), .D(men_men_n540_), .Y(men_men_n1238_));
  AN3        u1210(.A(men_men_n1238_), .B(men_men_n1225_), .C(men_men_n1216_), .Y(men_men_n1239_));
  NA2        u1211(.A(men_men_n558_), .B(men_men_n102_), .Y(men_men_n1240_));
  NA3        u1212(.A(men_men_n586_), .B(men_men_n1240_), .C(men_men_n251_), .Y(men_men_n1241_));
  NA2        u1213(.A(men_men_n1151_), .B(men_men_n558_), .Y(men_men_n1242_));
  NA4        u1214(.A(men_men_n681_), .B(men_men_n213_), .C(men_men_n229_), .D(men_men_n166_), .Y(men_men_n1243_));
  NA3        u1215(.A(men_men_n1243_), .B(men_men_n1242_), .C(men_men_n311_), .Y(men_men_n1244_));
  OAI210     u1216(.A0(men_men_n484_), .A1(men_men_n121_), .B0(men_men_n900_), .Y(men_men_n1245_));
  AOI220     u1217(.A0(men_men_n1245_), .A1(men_men_n1188_), .B0(men_men_n585_), .B1(men_men_n428_), .Y(men_men_n1246_));
  OR4        u1218(.A(men_men_n1087_), .B(men_men_n284_), .C(men_men_n231_), .D(e), .Y(men_men_n1247_));
  NO2        u1219(.A(men_men_n225_), .B(men_men_n222_), .Y(men_men_n1248_));
  NA2        u1220(.A(n), .B(e), .Y(men_men_n1249_));
  NO2        u1221(.A(men_men_n1249_), .B(men_men_n150_), .Y(men_men_n1250_));
  AOI220     u1222(.A0(men_men_n1250_), .A1(men_men_n286_), .B0(men_men_n881_), .B1(men_men_n1248_), .Y(men_men_n1251_));
  OAI210     u1223(.A0(men_men_n374_), .A1(men_men_n328_), .B0(men_men_n467_), .Y(men_men_n1252_));
  NA4        u1224(.A(men_men_n1252_), .B(men_men_n1251_), .C(men_men_n1247_), .D(men_men_n1246_), .Y(men_men_n1253_));
  AOI210     u1225(.A0(men_men_n1250_), .A1(men_men_n885_), .B0(men_men_n855_), .Y(men_men_n1254_));
  AOI220     u1226(.A0(men_men_n994_), .A1(men_men_n602_), .B0(men_men_n681_), .B1(men_men_n254_), .Y(men_men_n1255_));
  NO2        u1227(.A(men_men_n68_), .B(h), .Y(men_men_n1256_));
  NO3        u1228(.A(men_men_n1087_), .B(men_men_n1085_), .C(men_men_n762_), .Y(men_men_n1257_));
  NO2        u1229(.A(men_men_n1122_), .B(men_men_n134_), .Y(men_men_n1258_));
  AN2        u1230(.A(men_men_n1258_), .B(men_men_n1137_), .Y(men_men_n1259_));
  OAI210     u1231(.A0(men_men_n1259_), .A1(men_men_n1257_), .B0(men_men_n1256_), .Y(men_men_n1260_));
  NA4        u1232(.A(men_men_n1260_), .B(men_men_n1255_), .C(men_men_n1254_), .D(men_men_n902_), .Y(men_men_n1261_));
  NO4        u1233(.A(men_men_n1261_), .B(men_men_n1253_), .C(men_men_n1244_), .D(men_men_n1241_), .Y(men_men_n1262_));
  NA2        u1234(.A(men_men_n872_), .B(men_men_n795_), .Y(men_men_n1263_));
  NA4        u1235(.A(men_men_n1263_), .B(men_men_n1262_), .C(men_men_n1239_), .D(men_men_n1209_), .Y(men01));
  AN2        u1236(.A(men_men_n1064_), .B(men_men_n1062_), .Y(men_men_n1265_));
  NO4        u1237(.A(men_men_n839_), .B(men_men_n831_), .C(men_men_n498_), .D(men_men_n295_), .Y(men_men_n1266_));
  NO2        u1238(.A(men_men_n619_), .B(men_men_n304_), .Y(men_men_n1267_));
  OAI210     u1239(.A0(men_men_n1267_), .A1(men_men_n412_), .B0(i), .Y(men_men_n1268_));
  NA3        u1240(.A(men_men_n1268_), .B(men_men_n1266_), .C(men_men_n1265_), .Y(men_men_n1269_));
  NA2        u1241(.A(men_men_n615_), .B(men_men_n90_), .Y(men_men_n1270_));
  NA2        u1242(.A(men_men_n578_), .B(men_men_n283_), .Y(men_men_n1271_));
  NA2        u1243(.A(men_men_n1001_), .B(men_men_n1271_), .Y(men_men_n1272_));
  NA4        u1244(.A(men_men_n1272_), .B(men_men_n1270_), .C(men_men_n951_), .D(men_men_n348_), .Y(men_men_n1273_));
  NA2        u1245(.A(men_men_n741_), .B(men_men_n97_), .Y(men_men_n1274_));
  OAI220     u1246(.A0(men_men_n1274_), .A1(i), .B0(men_men_n370_), .B1(men_men_n299_), .Y(men_men_n1275_));
  OAI210     u1247(.A0(men_men_n818_), .A1(men_men_n632_), .B0(men_men_n1243_), .Y(men_men_n1276_));
  AOI210     u1248(.A0(men_men_n1275_), .A1(men_men_n668_), .B0(men_men_n1276_), .Y(men_men_n1277_));
  NA2        u1249(.A(men_men_n119_), .B(l), .Y(men_men_n1278_));
  OA220      u1250(.A0(men_men_n1278_), .A1(men_men_n612_), .B0(men_men_n694_), .B1(men_men_n386_), .Y(men_men_n1279_));
  NA3        u1251(.A(men_men_n1279_), .B(men_men_n1277_), .C(men_men_n935_), .Y(men_men_n1280_));
  NO3        u1252(.A(men_men_n819_), .B(men_men_n708_), .C(men_men_n534_), .Y(men_men_n1281_));
  NA4        u1253(.A(men_men_n741_), .B(men_men_n97_), .C(men_men_n45_), .D(men_men_n221_), .Y(men_men_n1282_));
  OA220      u1254(.A0(men_men_n1282_), .A1(men_men_n702_), .B0(men_men_n202_), .B1(men_men_n200_), .Y(men_men_n1283_));
  NA3        u1255(.A(men_men_n1283_), .B(men_men_n1281_), .C(men_men_n140_), .Y(men_men_n1284_));
  NO4        u1256(.A(men_men_n1284_), .B(men_men_n1280_), .C(men_men_n1273_), .D(men_men_n1269_), .Y(men_men_n1285_));
  NA2        u1257(.A(men_men_n1218_), .B(men_men_n214_), .Y(men_men_n1286_));
  OAI210     u1258(.A0(men_men_n1286_), .A1(men_men_n317_), .B0(men_men_n553_), .Y(men_men_n1287_));
  NA2        u1259(.A(men_men_n561_), .B(men_men_n414_), .Y(men_men_n1288_));
  NA2        u1260(.A(men_men_n76_), .B(i), .Y(men_men_n1289_));
  AOI210     u1261(.A0(men_men_n618_), .A1(men_men_n612_), .B0(men_men_n1289_), .Y(men_men_n1290_));
  NOi21      u1262(.An(men_men_n587_), .B(men_men_n609_), .Y(men_men_n1291_));
  AOI210     u1263(.A0(men_men_n1291_), .A1(men_men_n1288_), .B0(men_men_n1290_), .Y(men_men_n1292_));
  AOI210     u1264(.A0(men_men_n211_), .A1(men_men_n89_), .B0(men_men_n221_), .Y(men_men_n1293_));
  OAI210     u1265(.A0(men_men_n845_), .A1(men_men_n445_), .B0(men_men_n1293_), .Y(men_men_n1294_));
  NA2        u1266(.A(men_men_n210_), .B(men_men_n34_), .Y(men_men_n1295_));
  OR2        u1267(.A(men_men_n1295_), .B(men_men_n347_), .Y(men_men_n1296_));
  NA4        u1268(.A(men_men_n1296_), .B(men_men_n1294_), .C(men_men_n1292_), .D(men_men_n1287_), .Y(men_men_n1297_));
  AOI210     u1269(.A0(men_men_n624_), .A1(men_men_n119_), .B0(men_men_n630_), .Y(men_men_n1298_));
  OAI210     u1270(.A0(men_men_n1278_), .A1(men_men_n621_), .B0(men_men_n1298_), .Y(men_men_n1299_));
  NA2        u1271(.A(men_men_n294_), .B(men_men_n202_), .Y(men_men_n1300_));
  OAI210     u1272(.A0(men_men_n1300_), .A1(men_men_n403_), .B0(men_men_n699_), .Y(men_men_n1301_));
  NO3        u1273(.A(men_men_n854_), .B(men_men_n211_), .C(men_men_n426_), .Y(men_men_n1302_));
  NO2        u1274(.A(men_men_n1302_), .B(men_men_n998_), .Y(men_men_n1303_));
  NA3        u1275(.A(men_men_n1303_), .B(men_men_n1301_), .C(men_men_n821_), .Y(men_men_n1304_));
  NO3        u1276(.A(men_men_n1304_), .B(men_men_n1299_), .C(men_men_n1297_), .Y(men_men_n1305_));
  NA3        u1277(.A(men_men_n633_), .B(men_men_n29_), .C(f), .Y(men_men_n1306_));
  NO2        u1278(.A(men_men_n1306_), .B(men_men_n211_), .Y(men_men_n1307_));
  AOI210     u1279(.A0(men_men_n527_), .A1(men_men_n58_), .B0(men_men_n1307_), .Y(men_men_n1308_));
  OR3        u1280(.A(men_men_n1274_), .B(men_men_n634_), .C(i), .Y(men_men_n1309_));
  NA3        u1281(.A(men_men_n776_), .B(men_men_n76_), .C(i), .Y(men_men_n1310_));
  AOI210     u1282(.A0(men_men_n1310_), .A1(men_men_n1282_), .B0(men_men_n1017_), .Y(men_men_n1311_));
  NO2        u1283(.A(men_men_n214_), .B(men_men_n112_), .Y(men_men_n1312_));
  NO3        u1284(.A(men_men_n1312_), .B(men_men_n1311_), .C(men_men_n1214_), .Y(men_men_n1313_));
  NA4        u1285(.A(men_men_n1313_), .B(men_men_n1309_), .C(men_men_n1308_), .D(men_men_n794_), .Y(men_men_n1314_));
  NO2        u1286(.A(men_men_n1006_), .B(men_men_n241_), .Y(men_men_n1315_));
  NO2        u1287(.A(men_men_n1007_), .B(men_men_n580_), .Y(men_men_n1316_));
  OAI210     u1288(.A0(men_men_n1316_), .A1(men_men_n1315_), .B0(men_men_n356_), .Y(men_men_n1317_));
  NA2        u1289(.A(men_men_n597_), .B(men_men_n595_), .Y(men_men_n1318_));
  NO3        u1290(.A(men_men_n81_), .B(men_men_n315_), .C(men_men_n45_), .Y(men_men_n1319_));
  NA2        u1291(.A(men_men_n1319_), .B(men_men_n577_), .Y(men_men_n1320_));
  NA3        u1292(.A(men_men_n1320_), .B(men_men_n1318_), .C(men_men_n704_), .Y(men_men_n1321_));
  OR2        u1293(.A(men_men_n1218_), .B(men_men_n1211_), .Y(men_men_n1322_));
  NO2        u1294(.A(men_men_n386_), .B(men_men_n73_), .Y(men_men_n1323_));
  AOI210     u1295(.A0(men_men_n767_), .A1(men_men_n648_), .B0(men_men_n1323_), .Y(men_men_n1324_));
  NA3        u1296(.A(men_men_n1324_), .B(men_men_n1322_), .C(men_men_n404_), .Y(men_men_n1325_));
  NOi41      u1297(.An(men_men_n1317_), .B(men_men_n1325_), .C(men_men_n1321_), .D(men_men_n1314_), .Y(men_men_n1326_));
  NO2        u1298(.A(men_men_n133_), .B(men_men_n45_), .Y(men_men_n1327_));
  NO2        u1299(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1328_));
  AO220      u1300(.A0(men_men_n1328_), .A1(men_men_n654_), .B0(men_men_n1327_), .B1(men_men_n739_), .Y(men_men_n1329_));
  NA2        u1301(.A(men_men_n1329_), .B(men_men_n356_), .Y(men_men_n1330_));
  INV        u1302(.A(men_men_n137_), .Y(men_men_n1331_));
  NO3        u1303(.A(men_men_n1135_), .B(men_men_n182_), .C(men_men_n87_), .Y(men_men_n1332_));
  AOI220     u1304(.A0(men_men_n1332_), .A1(men_men_n1331_), .B0(men_men_n1319_), .B1(men_men_n1008_), .Y(men_men_n1333_));
  NA2        u1305(.A(men_men_n1333_), .B(men_men_n1330_), .Y(men_men_n1334_));
  NO2        u1306(.A(men_men_n645_), .B(men_men_n644_), .Y(men_men_n1335_));
  NO4        u1307(.A(men_men_n1135_), .B(men_men_n1335_), .C(men_men_n180_), .D(men_men_n87_), .Y(men_men_n1336_));
  NO3        u1308(.A(men_men_n1336_), .B(men_men_n1334_), .C(men_men_n672_), .Y(men_men_n1337_));
  NA4        u1309(.A(men_men_n1337_), .B(men_men_n1326_), .C(men_men_n1305_), .D(men_men_n1285_), .Y(men06));
  NO2        u1310(.A(men_men_n427_), .B(men_men_n584_), .Y(men_men_n1339_));
  NO2        u1311(.A(men_men_n769_), .B(i), .Y(men_men_n1340_));
  OAI210     u1312(.A0(men_men_n1340_), .A1(men_men_n279_), .B0(men_men_n1339_), .Y(men_men_n1341_));
  NO2        u1313(.A(men_men_n233_), .B(men_men_n104_), .Y(men_men_n1342_));
  OAI210     u1314(.A0(men_men_n1342_), .A1(men_men_n1332_), .B0(men_men_n400_), .Y(men_men_n1343_));
  NO3        u1315(.A(men_men_n628_), .B(men_men_n843_), .C(men_men_n631_), .Y(men_men_n1344_));
  OR2        u1316(.A(men_men_n1344_), .B(men_men_n922_), .Y(men_men_n1345_));
  NA4        u1317(.A(men_men_n1345_), .B(men_men_n1343_), .C(men_men_n1341_), .D(men_men_n1317_), .Y(men_men_n1346_));
  NO3        u1318(.A(men_men_n1346_), .B(men_men_n1321_), .C(men_men_n267_), .Y(men_men_n1347_));
  NO2        u1319(.A(men_men_n315_), .B(men_men_n45_), .Y(men_men_n1348_));
  AOI210     u1320(.A0(men_men_n1348_), .A1(men_men_n1009_), .B0(men_men_n1315_), .Y(men_men_n1349_));
  AOI210     u1321(.A0(men_men_n1348_), .A1(men_men_n581_), .B0(men_men_n1329_), .Y(men_men_n1350_));
  AOI210     u1322(.A0(men_men_n1350_), .A1(men_men_n1349_), .B0(men_men_n353_), .Y(men_men_n1351_));
  NO2        u1323(.A(men_men_n537_), .B(men_men_n177_), .Y(men_men_n1352_));
  NOi21      u1324(.An(men_men_n139_), .B(men_men_n45_), .Y(men_men_n1353_));
  NO2        u1325(.A(men_men_n638_), .B(men_men_n1158_), .Y(men_men_n1354_));
  NO2        u1326(.A(men_men_n480_), .B(men_men_n258_), .Y(men_men_n1355_));
  NO4        u1327(.A(men_men_n1355_), .B(men_men_n1354_), .C(men_men_n1353_), .D(men_men_n1352_), .Y(men_men_n1356_));
  OR2        u1328(.A(men_men_n629_), .B(men_men_n627_), .Y(men_men_n1357_));
  NO2        u1329(.A(men_men_n385_), .B(men_men_n138_), .Y(men_men_n1358_));
  AOI210     u1330(.A0(men_men_n1358_), .A1(men_men_n615_), .B0(men_men_n1357_), .Y(men_men_n1359_));
  NA2        u1331(.A(men_men_n1359_), .B(men_men_n1356_), .Y(men_men_n1360_));
  NO2        u1332(.A(men_men_n785_), .B(men_men_n384_), .Y(men_men_n1361_));
  NO3        u1333(.A(men_men_n709_), .B(men_men_n796_), .C(men_men_n668_), .Y(men_men_n1362_));
  NOi21      u1334(.An(men_men_n1361_), .B(men_men_n1362_), .Y(men_men_n1363_));
  AN2        u1335(.A(men_men_n994_), .B(men_men_n677_), .Y(men_men_n1364_));
  NO4        u1336(.A(men_men_n1364_), .B(men_men_n1363_), .C(men_men_n1360_), .D(men_men_n1351_), .Y(men_men_n1365_));
  NO2        u1337(.A(men_men_n838_), .B(men_men_n290_), .Y(men_men_n1366_));
  OAI220     u1338(.A0(men_men_n769_), .A1(men_men_n47_), .B0(men_men_n233_), .B1(men_men_n647_), .Y(men_men_n1367_));
  OAI210     u1339(.A0(men_men_n290_), .A1(c), .B0(men_men_n675_), .Y(men_men_n1368_));
  AOI220     u1340(.A0(men_men_n1368_), .A1(men_men_n1367_), .B0(men_men_n1366_), .B1(men_men_n279_), .Y(men_men_n1369_));
  NO3        u1341(.A(men_men_n253_), .B(men_men_n104_), .C(men_men_n297_), .Y(men_men_n1370_));
  OAI220     u1342(.A0(men_men_n733_), .A1(men_men_n258_), .B0(men_men_n533_), .B1(men_men_n537_), .Y(men_men_n1371_));
  OAI210     u1343(.A0(l), .A1(i), .B0(k), .Y(men_men_n1372_));
  NO3        u1344(.A(men_men_n1372_), .B(men_men_n626_), .C(j), .Y(men_men_n1373_));
  NOi21      u1345(.An(men_men_n1373_), .B(men_men_n702_), .Y(men_men_n1374_));
  NO4        u1346(.A(men_men_n1374_), .B(men_men_n1371_), .C(men_men_n1370_), .D(men_men_n1160_), .Y(men_men_n1375_));
  NA4        u1347(.A(men_men_n829_), .B(men_men_n828_), .C(men_men_n455_), .D(men_men_n914_), .Y(men_men_n1376_));
  NAi31      u1348(.An(men_men_n785_), .B(men_men_n1376_), .C(men_men_n210_), .Y(men_men_n1377_));
  NA4        u1349(.A(men_men_n1377_), .B(men_men_n1375_), .C(men_men_n1369_), .D(men_men_n1255_), .Y(men_men_n1378_));
  NOi31      u1350(.An(men_men_n1344_), .B(men_men_n483_), .C(men_men_n413_), .Y(men_men_n1379_));
  OR3        u1351(.A(men_men_n1379_), .B(men_men_n818_), .C(men_men_n564_), .Y(men_men_n1380_));
  OR3        u1352(.A(men_men_n388_), .B(men_men_n233_), .C(men_men_n647_), .Y(men_men_n1381_));
  AOI210     u1353(.A0(men_men_n597_), .A1(men_men_n467_), .B0(men_men_n390_), .Y(men_men_n1382_));
  NA2        u1354(.A(men_men_n1373_), .B(men_men_n825_), .Y(men_men_n1383_));
  NA4        u1355(.A(men_men_n1383_), .B(men_men_n1382_), .C(men_men_n1381_), .D(men_men_n1380_), .Y(men_men_n1384_));
  AOI220     u1356(.A0(men_men_n1361_), .A1(men_men_n795_), .B0(men_men_n1358_), .B1(men_men_n247_), .Y(men_men_n1385_));
  AN2        u1357(.A(men_men_n966_), .B(men_men_n965_), .Y(men_men_n1386_));
  NO4        u1358(.A(men_men_n1386_), .B(men_men_n912_), .C(men_men_n523_), .D(men_men_n501_), .Y(men_men_n1387_));
  NA2        u1359(.A(men_men_n1387_), .B(men_men_n1385_), .Y(men_men_n1388_));
  NAi21      u1360(.An(j), .B(i), .Y(men_men_n1389_));
  NO4        u1361(.A(men_men_n1335_), .B(men_men_n1389_), .C(men_men_n461_), .D(men_men_n244_), .Y(men_men_n1390_));
  NO4        u1362(.A(men_men_n1390_), .B(men_men_n1388_), .C(men_men_n1384_), .D(men_men_n1378_), .Y(men_men_n1391_));
  NA4        u1363(.A(men_men_n1391_), .B(men_men_n1365_), .C(men_men_n1347_), .D(men_men_n1337_), .Y(men07));
  NOi21      u1364(.An(j), .B(k), .Y(men_men_n1393_));
  NA4        u1365(.A(men_men_n185_), .B(men_men_n109_), .C(men_men_n1393_), .D(f), .Y(men_men_n1394_));
  NAi32      u1366(.An(m), .Bn(b), .C(n), .Y(men_men_n1395_));
  NO3        u1367(.A(men_men_n1395_), .B(g), .C(f), .Y(men_men_n1396_));
  OAI210     u1368(.A0(men_men_n338_), .A1(men_men_n503_), .B0(men_men_n1396_), .Y(men_men_n1397_));
  NAi21      u1369(.An(f), .B(c), .Y(men_men_n1398_));
  OR2        u1370(.A(e), .B(d), .Y(men_men_n1399_));
  NOi31      u1371(.An(n), .B(m), .C(b), .Y(men_men_n1400_));
  NO3        u1372(.A(men_men_n134_), .B(men_men_n469_), .C(h), .Y(men_men_n1401_));
  NA2        u1373(.A(men_men_n1397_), .B(men_men_n1394_), .Y(men_men_n1402_));
  NOi41      u1374(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1403_));
  NA3        u1375(.A(men_men_n1403_), .B(men_men_n904_), .C(men_men_n429_), .Y(men_men_n1404_));
  NO2        u1376(.A(men_men_n1404_), .B(men_men_n56_), .Y(men_men_n1405_));
  NA2        u1377(.A(men_men_n1137_), .B(men_men_n229_), .Y(men_men_n1406_));
  NO2        u1378(.A(men_men_n1406_), .B(men_men_n61_), .Y(men_men_n1407_));
  NO2        u1379(.A(k), .B(i), .Y(men_men_n1408_));
  NA3        u1380(.A(men_men_n1408_), .B(men_men_n934_), .C(men_men_n185_), .Y(men_men_n1409_));
  NA2        u1381(.A(men_men_n87_), .B(men_men_n45_), .Y(men_men_n1410_));
  NO2        u1382(.A(men_men_n1093_), .B(men_men_n461_), .Y(men_men_n1411_));
  NA3        u1383(.A(men_men_n1411_), .B(men_men_n1410_), .C(men_men_n222_), .Y(men_men_n1412_));
  NO2        u1384(.A(men_men_n1107_), .B(men_men_n322_), .Y(men_men_n1413_));
  NA2        u1385(.A(men_men_n1256_), .B(men_men_n305_), .Y(men_men_n1414_));
  NA3        u1386(.A(men_men_n1414_), .B(men_men_n1412_), .C(men_men_n1409_), .Y(men_men_n1415_));
  NO4        u1387(.A(men_men_n1415_), .B(men_men_n1407_), .C(men_men_n1405_), .D(men_men_n1402_), .Y(men_men_n1416_));
  NO3        u1388(.A(e), .B(d), .C(c), .Y(men_men_n1417_));
  AOI210     u1389(.A0(men_men_n1114_), .A1(men_men_n222_), .B0(men_men_n1417_), .Y(men_men_n1418_));
  OAI210     u1390(.A0(men_men_n134_), .A1(men_men_n222_), .B0(men_men_n635_), .Y(men_men_n1419_));
  NA2        u1391(.A(men_men_n1419_), .B(men_men_n1417_), .Y(men_men_n1420_));
  NO2        u1392(.A(men_men_n1420_), .B(men_men_n1418_), .Y(men_men_n1421_));
  OR2        u1393(.A(h), .B(f), .Y(men_men_n1422_));
  NO3        u1394(.A(n), .B(m), .C(i), .Y(men_men_n1423_));
  OAI210     u1395(.A0(men_men_n1159_), .A1(men_men_n161_), .B0(men_men_n1423_), .Y(men_men_n1424_));
  NO2        u1396(.A(i), .B(g), .Y(men_men_n1425_));
  OR3        u1397(.A(men_men_n1425_), .B(men_men_n1395_), .C(men_men_n72_), .Y(men_men_n1426_));
  OAI220     u1398(.A0(men_men_n1426_), .A1(men_men_n503_), .B0(men_men_n1424_), .B1(men_men_n1422_), .Y(men_men_n1427_));
  NA3        u1399(.A(men_men_n730_), .B(men_men_n716_), .C(men_men_n113_), .Y(men_men_n1428_));
  NA3        u1400(.A(men_men_n1400_), .B(men_men_n1102_), .C(men_men_n706_), .Y(men_men_n1429_));
  AOI210     u1401(.A0(men_men_n1429_), .A1(men_men_n1428_), .B0(men_men_n45_), .Y(men_men_n1430_));
  NA2        u1402(.A(men_men_n1423_), .B(men_men_n674_), .Y(men_men_n1431_));
  NO2        u1403(.A(l), .B(k), .Y(men_men_n1432_));
  NO3        u1404(.A(men_men_n461_), .B(d), .C(c), .Y(men_men_n1433_));
  NO3        u1405(.A(men_men_n1430_), .B(men_men_n1427_), .C(men_men_n1421_), .Y(men_men_n1434_));
  NO2        u1406(.A(men_men_n151_), .B(h), .Y(men_men_n1435_));
  NO2        u1407(.A(men_men_n1117_), .B(l), .Y(men_men_n1436_));
  NO2        u1408(.A(g), .B(c), .Y(men_men_n1437_));
  NA3        u1409(.A(men_men_n1437_), .B(men_men_n145_), .C(men_men_n193_), .Y(men_men_n1438_));
  NO2        u1410(.A(men_men_n1438_), .B(men_men_n1436_), .Y(men_men_n1439_));
  NA2        u1411(.A(men_men_n1439_), .B(men_men_n185_), .Y(men_men_n1440_));
  NO2        u1412(.A(men_men_n471_), .B(a), .Y(men_men_n1441_));
  NA3        u1413(.A(men_men_n1441_), .B(k), .C(men_men_n114_), .Y(men_men_n1442_));
  NO2        u1414(.A(i), .B(h), .Y(men_men_n1443_));
  NA2        u1415(.A(men_men_n1443_), .B(men_men_n229_), .Y(men_men_n1444_));
  AOI210     u1416(.A0(men_men_n1180_), .A1(h), .B0(men_men_n433_), .Y(men_men_n1445_));
  NA2        u1417(.A(men_men_n141_), .B(men_men_n229_), .Y(men_men_n1446_));
  AOI210     u1418(.A0(men_men_n268_), .A1(men_men_n117_), .B0(men_men_n553_), .Y(men_men_n1447_));
  OAI220     u1419(.A0(men_men_n1447_), .A1(men_men_n1444_), .B0(men_men_n1446_), .B1(men_men_n1445_), .Y(men_men_n1448_));
  NO2        u1420(.A(men_men_n792_), .B(men_men_n194_), .Y(men_men_n1449_));
  NOi31      u1421(.An(m), .B(n), .C(b), .Y(men_men_n1450_));
  NOi31      u1422(.An(f), .B(d), .C(c), .Y(men_men_n1451_));
  NA2        u1423(.A(men_men_n1451_), .B(men_men_n1450_), .Y(men_men_n1452_));
  INV        u1424(.A(men_men_n1452_), .Y(men_men_n1453_));
  NO3        u1425(.A(men_men_n1453_), .B(men_men_n1449_), .C(men_men_n1448_), .Y(men_men_n1454_));
  NA2        u1426(.A(men_men_n1128_), .B(men_men_n485_), .Y(men_men_n1455_));
  NO4        u1427(.A(men_men_n1455_), .B(men_men_n1102_), .C(men_men_n461_), .D(men_men_n45_), .Y(men_men_n1456_));
  OAI210     u1428(.A0(men_men_n188_), .A1(men_men_n548_), .B0(men_men_n1103_), .Y(men_men_n1457_));
  NO3        u1429(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1458_));
  INV        u1430(.A(men_men_n1457_), .Y(men_men_n1459_));
  NO2        u1431(.A(men_men_n1459_), .B(men_men_n1456_), .Y(men_men_n1460_));
  AN4        u1432(.A(men_men_n1460_), .B(men_men_n1454_), .C(men_men_n1442_), .D(men_men_n1440_), .Y(men_men_n1461_));
  NA2        u1433(.A(men_men_n1400_), .B(men_men_n397_), .Y(men_men_n1462_));
  NO2        u1434(.A(men_men_n1462_), .B(men_men_n1084_), .Y(men_men_n1463_));
  NA2        u1435(.A(men_men_n1433_), .B(men_men_n223_), .Y(men_men_n1464_));
  NO2        u1436(.A(men_men_n194_), .B(b), .Y(men_men_n1465_));
  AOI220     u1437(.A0(men_men_n1212_), .A1(men_men_n1465_), .B0(men_men_n1136_), .B1(men_men_n1455_), .Y(men_men_n1466_));
  NO2        u1438(.A(i), .B(men_men_n221_), .Y(men_men_n1467_));
  NA4        u1439(.A(men_men_n1186_), .B(men_men_n1467_), .C(men_men_n105_), .D(m), .Y(men_men_n1468_));
  NAi41      u1440(.An(men_men_n1463_), .B(men_men_n1468_), .C(men_men_n1466_), .D(men_men_n1464_), .Y(men_men_n1469_));
  NO4        u1441(.A(men_men_n134_), .B(g), .C(f), .D(e), .Y(men_men_n1470_));
  NA3        u1442(.A(men_men_n1408_), .B(men_men_n306_), .C(h), .Y(men_men_n1471_));
  NA2        u1443(.A(men_men_n201_), .B(men_men_n99_), .Y(men_men_n1472_));
  NA2        u1444(.A(men_men_n30_), .B(h), .Y(men_men_n1473_));
  NO2        u1445(.A(men_men_n1473_), .B(men_men_n1124_), .Y(men_men_n1474_));
  NOi41      u1446(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1475_));
  NA2        u1447(.A(men_men_n1475_), .B(men_men_n114_), .Y(men_men_n1476_));
  NA2        u1448(.A(men_men_n1403_), .B(men_men_n1432_), .Y(men_men_n1477_));
  NA2        u1449(.A(men_men_n1477_), .B(men_men_n1476_), .Y(men_men_n1478_));
  OR3        u1450(.A(men_men_n564_), .B(men_men_n563_), .C(men_men_n113_), .Y(men_men_n1479_));
  NA2        u1451(.A(men_men_n1157_), .B(men_men_n426_), .Y(men_men_n1480_));
  OAI220     u1452(.A0(men_men_n1480_), .A1(men_men_n454_), .B0(men_men_n1479_), .B1(men_men_n315_), .Y(men_men_n1481_));
  AO210      u1453(.A0(men_men_n1481_), .A1(men_men_n117_), .B0(men_men_n1478_), .Y(men_men_n1482_));
  NO3        u1454(.A(men_men_n1482_), .B(men_men_n1474_), .C(men_men_n1469_), .Y(men_men_n1483_));
  NA4        u1455(.A(men_men_n1483_), .B(men_men_n1461_), .C(men_men_n1434_), .D(men_men_n1416_), .Y(men_men_n1484_));
  NO2        u1456(.A(men_men_n1172_), .B(men_men_n111_), .Y(men_men_n1485_));
  NA2        u1457(.A(men_men_n397_), .B(men_men_n56_), .Y(men_men_n1486_));
  AOI210     u1458(.A0(men_men_n1486_), .A1(men_men_n1093_), .B0(men_men_n1431_), .Y(men_men_n1487_));
  NA2        u1459(.A(men_men_n223_), .B(men_men_n185_), .Y(men_men_n1488_));
  AOI210     u1460(.A0(men_men_n1488_), .A1(men_men_n1229_), .B0(men_men_n1486_), .Y(men_men_n1489_));
  NO2        u1461(.A(men_men_n1129_), .B(men_men_n1124_), .Y(men_men_n1490_));
  NO3        u1462(.A(men_men_n1490_), .B(men_men_n1489_), .C(men_men_n1487_), .Y(men_men_n1491_));
  NO2        u1463(.A(men_men_n409_), .B(j), .Y(men_men_n1492_));
  NA3        u1464(.A(men_men_n1458_), .B(men_men_n1399_), .C(men_men_n1157_), .Y(men_men_n1493_));
  NAi41      u1465(.An(men_men_n1443_), .B(men_men_n1115_), .C(men_men_n173_), .D(men_men_n154_), .Y(men_men_n1494_));
  NA2        u1466(.A(men_men_n1494_), .B(men_men_n1493_), .Y(men_men_n1495_));
  NA3        u1467(.A(g), .B(men_men_n1492_), .C(men_men_n163_), .Y(men_men_n1496_));
  INV        u1468(.A(men_men_n1496_), .Y(men_men_n1497_));
  NO3        u1469(.A(men_men_n785_), .B(men_men_n180_), .C(men_men_n429_), .Y(men_men_n1498_));
  NO3        u1470(.A(men_men_n1498_), .B(men_men_n1497_), .C(men_men_n1495_), .Y(men_men_n1499_));
  NO3        u1471(.A(men_men_n1124_), .B(men_men_n609_), .C(g), .Y(men_men_n1500_));
  NOi21      u1472(.An(men_men_n1488_), .B(men_men_n1500_), .Y(men_men_n1501_));
  AOI210     u1473(.A0(men_men_n1501_), .A1(men_men_n1472_), .B0(men_men_n1093_), .Y(men_men_n1502_));
  OR2        u1474(.A(n), .B(i), .Y(men_men_n1503_));
  OAI210     u1475(.A0(men_men_n1503_), .A1(men_men_n1114_), .B0(men_men_n49_), .Y(men_men_n1504_));
  AOI220     u1476(.A0(men_men_n1504_), .A1(men_men_n1220_), .B0(men_men_n859_), .B1(men_men_n201_), .Y(men_men_n1505_));
  INV        u1477(.A(men_men_n1505_), .Y(men_men_n1506_));
  OAI220     u1478(.A0(men_men_n700_), .A1(g), .B0(men_men_n233_), .B1(c), .Y(men_men_n1507_));
  AOI210     u1479(.A0(men_men_n1465_), .A1(men_men_n41_), .B0(men_men_n1507_), .Y(men_men_n1508_));
  NO2        u1480(.A(men_men_n233_), .B(k), .Y(men_men_n1509_));
  NO2        u1481(.A(men_men_n1508_), .B(men_men_n182_), .Y(men_men_n1510_));
  NO3        u1482(.A(men_men_n1510_), .B(men_men_n1506_), .C(men_men_n1502_), .Y(men_men_n1511_));
  NO2        u1483(.A(men_men_n49_), .B(men_men_n609_), .Y(men_men_n1512_));
  NO3        u1484(.A(men_men_n1139_), .B(men_men_n1399_), .C(men_men_n49_), .Y(men_men_n1513_));
  NA2        u1485(.A(men_men_n1140_), .B(men_men_n1512_), .Y(men_men_n1514_));
  NO2        u1486(.A(men_men_n1124_), .B(h), .Y(men_men_n1515_));
  NA3        u1487(.A(men_men_n1515_), .B(d), .C(men_men_n1085_), .Y(men_men_n1516_));
  OAI220     u1488(.A0(men_men_n1516_), .A1(c), .B0(men_men_n1514_), .B1(j), .Y(men_men_n1517_));
  NA3        u1489(.A(men_men_n1485_), .B(men_men_n485_), .C(f), .Y(men_men_n1518_));
  NA2        u1490(.A(men_men_n185_), .B(men_men_n113_), .Y(men_men_n1519_));
  NO2        u1491(.A(men_men_n1393_), .B(men_men_n42_), .Y(men_men_n1520_));
  AOI210     u1492(.A0(men_men_n114_), .A1(men_men_n40_), .B0(men_men_n1520_), .Y(men_men_n1521_));
  NO2        u1493(.A(men_men_n1521_), .B(men_men_n1518_), .Y(men_men_n1522_));
  AOI210     u1494(.A0(men_men_n548_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1523_));
  NA2        u1495(.A(men_men_n1523_), .B(men_men_n1441_), .Y(men_men_n1524_));
  NO2        u1496(.A(men_men_n1389_), .B(men_men_n180_), .Y(men_men_n1525_));
  NOi21      u1497(.An(d), .B(f), .Y(men_men_n1526_));
  NO3        u1498(.A(men_men_n1451_), .B(men_men_n1526_), .C(men_men_n40_), .Y(men_men_n1527_));
  NA2        u1499(.A(men_men_n1527_), .B(men_men_n1525_), .Y(men_men_n1528_));
  NO2        u1500(.A(men_men_n1399_), .B(f), .Y(men_men_n1529_));
  NA2        u1501(.A(men_men_n1441_), .B(men_men_n1520_), .Y(men_men_n1530_));
  NO2        u1502(.A(men_men_n315_), .B(c), .Y(men_men_n1531_));
  NA2        u1503(.A(men_men_n1531_), .B(men_men_n565_), .Y(men_men_n1532_));
  NA4        u1504(.A(men_men_n1532_), .B(men_men_n1530_), .C(men_men_n1528_), .D(men_men_n1524_), .Y(men_men_n1533_));
  NO3        u1505(.A(men_men_n1533_), .B(men_men_n1522_), .C(men_men_n1517_), .Y(men_men_n1534_));
  NA4        u1506(.A(men_men_n1534_), .B(men_men_n1511_), .C(men_men_n1499_), .D(men_men_n1491_), .Y(men_men_n1535_));
  NO3        u1507(.A(men_men_n1128_), .B(men_men_n1114_), .C(men_men_n40_), .Y(men_men_n1536_));
  OAI220     u1508(.A0(men_men_n485_), .A1(men_men_n315_), .B0(men_men_n133_), .B1(men_men_n59_), .Y(men_men_n1537_));
  OAI210     u1509(.A0(men_men_n1537_), .A1(men_men_n1536_), .B0(men_men_n1413_), .Y(men_men_n1538_));
  OAI210     u1510(.A0(men_men_n1470_), .A1(men_men_n1400_), .B0(men_men_n919_), .Y(men_men_n1539_));
  OAI220     u1511(.A0(men_men_n1081_), .A1(men_men_n134_), .B0(men_men_n700_), .B1(men_men_n180_), .Y(men_men_n1540_));
  NA2        u1512(.A(men_men_n1540_), .B(men_men_n653_), .Y(men_men_n1541_));
  NA3        u1513(.A(men_men_n1541_), .B(men_men_n1539_), .C(men_men_n1538_), .Y(men_men_n1542_));
  NA2        u1514(.A(men_men_n1437_), .B(men_men_n1526_), .Y(men_men_n1543_));
  NO2        u1515(.A(men_men_n1543_), .B(m), .Y(men_men_n1544_));
  NA3        u1516(.A(men_men_n1137_), .B(men_men_n109_), .C(men_men_n229_), .Y(men_men_n1545_));
  OAI220     u1517(.A0(men_men_n155_), .A1(men_men_n187_), .B0(men_men_n469_), .B1(g), .Y(men_men_n1546_));
  OAI210     u1518(.A0(men_men_n1546_), .A1(men_men_n111_), .B0(men_men_n1450_), .Y(men_men_n1547_));
  NA2        u1519(.A(men_men_n1547_), .B(men_men_n1545_), .Y(men_men_n1548_));
  NO3        u1520(.A(men_men_n1548_), .B(men_men_n1544_), .C(men_men_n1542_), .Y(men_men_n1549_));
  NO2        u1521(.A(men_men_n1398_), .B(e), .Y(men_men_n1550_));
  NA2        u1522(.A(men_men_n1550_), .B(men_men_n424_), .Y(men_men_n1551_));
  OAI210     u1523(.A0(men_men_n1529_), .A1(men_men_n1167_), .B0(men_men_n664_), .Y(men_men_n1552_));
  OR3        u1524(.A(men_men_n1509_), .B(men_men_n1256_), .C(men_men_n134_), .Y(men_men_n1553_));
  OAI220     u1525(.A0(men_men_n1553_), .A1(men_men_n1551_), .B0(men_men_n1552_), .B1(men_men_n463_), .Y(men_men_n1554_));
  NO3        u1526(.A(men_men_n1479_), .B(men_men_n370_), .C(a), .Y(men_men_n1555_));
  NO2        u1527(.A(men_men_n1555_), .B(men_men_n1554_), .Y(men_men_n1556_));
  NO2        u1528(.A(men_men_n187_), .B(c), .Y(men_men_n1557_));
  OAI210     u1529(.A0(men_men_n1557_), .A1(men_men_n1550_), .B0(men_men_n185_), .Y(men_men_n1558_));
  AOI220     u1530(.A0(men_men_n1558_), .A1(men_men_n1116_), .B0(men_men_n555_), .B1(men_men_n384_), .Y(men_men_n1559_));
  NA2        u1531(.A(men_men_n563_), .B(g), .Y(men_men_n1560_));
  AOI210     u1532(.A0(men_men_n1560_), .A1(men_men_n1433_), .B0(men_men_n1513_), .Y(men_men_n1561_));
  NO2        u1533(.A(men_men_n1561_), .B(men_men_n221_), .Y(men_men_n1562_));
  AOI210     u1534(.A0(men_men_n939_), .A1(men_men_n435_), .B0(men_men_n106_), .Y(men_men_n1563_));
  OR2        u1535(.A(men_men_n1563_), .B(men_men_n563_), .Y(men_men_n1564_));
  NO2        u1536(.A(men_men_n1564_), .B(men_men_n180_), .Y(men_men_n1565_));
  NA2        u1537(.A(men_men_n1401_), .B(men_men_n188_), .Y(men_men_n1566_));
  NO2        u1538(.A(men_men_n49_), .B(l), .Y(men_men_n1567_));
  INV        u1539(.A(men_men_n503_), .Y(men_men_n1568_));
  OAI210     u1540(.A0(men_men_n1568_), .A1(men_men_n1140_), .B0(men_men_n1567_), .Y(men_men_n1569_));
  NO2        u1541(.A(m), .B(i), .Y(men_men_n1570_));
  BUFFER     u1542(.A(men_men_n1570_), .Y(men_men_n1571_));
  NA2        u1543(.A(men_men_n1571_), .B(men_men_n1435_), .Y(men_men_n1572_));
  NA3        u1544(.A(men_men_n1572_), .B(men_men_n1569_), .C(men_men_n1566_), .Y(men_men_n1573_));
  NO4        u1545(.A(men_men_n1573_), .B(men_men_n1565_), .C(men_men_n1562_), .D(men_men_n1559_), .Y(men_men_n1574_));
  NA3        u1546(.A(men_men_n1574_), .B(men_men_n1556_), .C(men_men_n1549_), .Y(men_men_n1575_));
  NA3        u1547(.A(men_men_n1000_), .B(men_men_n141_), .C(men_men_n46_), .Y(men_men_n1576_));
  AOI210     u1548(.A0(men_men_n152_), .A1(c), .B0(men_men_n1576_), .Y(men_men_n1577_));
  INV        u1549(.A(men_men_n191_), .Y(men_men_n1578_));
  NA2        u1550(.A(men_men_n1578_), .B(men_men_n1515_), .Y(men_men_n1579_));
  AO210      u1551(.A0(men_men_n135_), .A1(l), .B0(men_men_n1462_), .Y(men_men_n1580_));
  NO2        u1552(.A(men_men_n72_), .B(c), .Y(men_men_n1581_));
  NO4        u1553(.A(men_men_n1422_), .B(men_men_n192_), .C(men_men_n469_), .D(men_men_n45_), .Y(men_men_n1582_));
  AOI210     u1554(.A0(men_men_n1525_), .A1(men_men_n1581_), .B0(men_men_n1582_), .Y(men_men_n1583_));
  NA3        u1555(.A(men_men_n1583_), .B(men_men_n1580_), .C(men_men_n1579_), .Y(men_men_n1584_));
  NO2        u1556(.A(men_men_n1584_), .B(men_men_n1577_), .Y(men_men_n1585_));
  NO4        u1557(.A(men_men_n233_), .B(men_men_n192_), .C(men_men_n268_), .D(k), .Y(men_men_n1586_));
  AOI210     u1558(.A0(men_men_n161_), .A1(men_men_n56_), .B0(men_men_n1550_), .Y(men_men_n1587_));
  NO2        u1559(.A(men_men_n1587_), .B(men_men_n1519_), .Y(men_men_n1588_));
  NO2        u1560(.A(men_men_n1576_), .B(men_men_n111_), .Y(men_men_n1589_));
  NO3        u1561(.A(men_men_n1589_), .B(men_men_n1588_), .C(men_men_n1586_), .Y(men_men_n1590_));
  NO2        u1562(.A(men_men_n1518_), .B(men_men_n69_), .Y(men_men_n1591_));
  NA2        u1563(.A(men_men_n59_), .B(a), .Y(men_men_n1592_));
  NO2        u1564(.A(men_men_n1480_), .B(men_men_n1592_), .Y(men_men_n1593_));
  NO2        u1565(.A(men_men_n1593_), .B(men_men_n1591_), .Y(men_men_n1594_));
  NA3        u1566(.A(men_men_n1594_), .B(men_men_n1590_), .C(men_men_n1585_), .Y(men_men_n1595_));
  OR4        u1567(.A(men_men_n1595_), .B(men_men_n1575_), .C(men_men_n1535_), .D(men_men_n1484_), .Y(men04));
  NOi31      u1568(.An(men_men_n1470_), .B(men_men_n1471_), .C(men_men_n1087_), .Y(men_men_n1597_));
  NA2        u1569(.A(men_men_n1529_), .B(men_men_n859_), .Y(men_men_n1598_));
  NO4        u1570(.A(men_men_n1598_), .B(men_men_n1076_), .C(men_men_n504_), .D(j), .Y(men_men_n1599_));
  OR3        u1571(.A(men_men_n1599_), .B(men_men_n1597_), .C(men_men_n1105_), .Y(men_men_n1600_));
  NO3        u1572(.A(men_men_n1410_), .B(men_men_n91_), .C(k), .Y(men_men_n1601_));
  AOI210     u1573(.A0(men_men_n1601_), .A1(men_men_n1098_), .B0(men_men_n1231_), .Y(men_men_n1602_));
  NA2        u1574(.A(men_men_n1602_), .B(men_men_n1260_), .Y(men_men_n1603_));
  NO4        u1575(.A(men_men_n1603_), .B(men_men_n1600_), .C(men_men_n1113_), .D(men_men_n1092_), .Y(men_men_n1604_));
  NA4        u1576(.A(men_men_n1604_), .B(men_men_n1169_), .C(men_men_n1155_), .D(men_men_n1143_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule