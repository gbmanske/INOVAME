// Benchmark "top" written by ABC on Thu Jun 20 14:00:09 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n138_, new_new_n139_,
    new_new_n140_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1024_, new_new_n1025_, new_new_n1026_, new_new_n1027_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(mai1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n51_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  INV        g0062(.A(i_6_), .Y(new_new_n85_));
  OR4        g0063(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n86_));
  INV        g0064(.A(new_new_n86_), .Y(new_new_n87_));
  NO2        g0065(.A(i_2_), .B(i_7_), .Y(new_new_n88_));
  NAi21      g0066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g0067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g0068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n63_), .Y(new_new_n91_));
  NA2        g0069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  NO3        g0070(.A(new_new_n92_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n93_));
  NO2        g0071(.A(new_new_n93_), .B(new_new_n91_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n1027_), .B0(new_new_n80_), .Y(new_new_n95_));
  AN3        g0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g0074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NO2        g0075(.A(i_5_), .B(i_8_), .Y(new_new_n98_));
  NOi21      g0076(.An(new_new_n98_), .B(new_new_n97_), .Y(new_new_n99_));
  AOI220     g0077(.A0(new_new_n99_), .A1(new_new_n62_), .B0(new_new_n96_), .B1(new_new_n32_), .Y(new_new_n100_));
  INV        g0078(.A(i_7_), .Y(new_new_n101_));
  NA2        g0079(.A(new_new_n47_), .B(new_new_n101_), .Y(new_new_n102_));
  NO2        g0080(.A(i_0_), .B(i_5_), .Y(new_new_n103_));
  NO2        g0081(.A(new_new_n103_), .B(new_new_n85_), .Y(new_new_n104_));
  NA2        g0082(.A(i_12_), .B(i_3_), .Y(new_new_n105_));
  INV        g0083(.A(new_new_n105_), .Y(new_new_n106_));
  NA3        g0084(.A(new_new_n106_), .B(new_new_n104_), .C(new_new_n102_), .Y(new_new_n107_));
  NAi21      g0085(.An(i_7_), .B(i_11_), .Y(new_new_n108_));
  NO3        g0086(.A(new_new_n108_), .B(new_new_n89_), .C(new_new_n54_), .Y(new_new_n109_));
  AN2        g0087(.A(i_2_), .B(i_10_), .Y(new_new_n110_));
  NO2        g0088(.A(new_new_n110_), .B(i_7_), .Y(new_new_n111_));
  OR2        g0089(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n112_));
  NO2        g0090(.A(i_8_), .B(new_new_n101_), .Y(new_new_n113_));
  NO3        g0091(.A(new_new_n113_), .B(new_new_n112_), .C(new_new_n111_), .Y(new_new_n114_));
  NA2        g0092(.A(i_12_), .B(i_7_), .Y(new_new_n115_));
  NO2        g0093(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n116_));
  NA2        g0094(.A(new_new_n116_), .B(i_0_), .Y(new_new_n117_));
  NA2        g0095(.A(i_11_), .B(i_12_), .Y(new_new_n118_));
  OAI210     g0096(.A0(new_new_n117_), .A1(new_new_n115_), .B0(new_new_n118_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n119_), .B(new_new_n114_), .Y(new_new_n120_));
  NAi41      g0098(.An(new_new_n109_), .B(new_new_n120_), .C(new_new_n107_), .D(new_new_n100_), .Y(new_new_n121_));
  NOi21      g0099(.An(i_1_), .B(i_5_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(i_11_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n124_));
  NA2        g0102(.A(i_7_), .B(new_new_n25_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n125_), .B(new_new_n124_), .Y(new_new_n126_));
  NO2        g0104(.A(new_new_n126_), .B(new_new_n47_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n128_));
  NAi21      g0106(.An(i_3_), .B(i_8_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n129_), .B(new_new_n62_), .Y(new_new_n130_));
  NOi31      g0108(.An(new_new_n130_), .B(new_new_n128_), .C(new_new_n127_), .Y(new_new_n131_));
  NO2        g0109(.A(i_1_), .B(new_new_n85_), .Y(new_new_n132_));
  NO2        g0110(.A(i_6_), .B(i_5_), .Y(new_new_n133_));
  NA2        g0111(.A(new_new_n133_), .B(i_3_), .Y(new_new_n134_));
  OAI220     g0112(.A0(new_new_n134_), .A1(new_new_n108_), .B0(new_new_n131_), .B1(new_new_n123_), .Y(new_new_n135_));
  NO3        g0113(.A(new_new_n135_), .B(new_new_n121_), .C(new_new_n95_), .Y(new_new_n136_));
  NA3        g0114(.A(new_new_n136_), .B(new_new_n79_), .C(new_new_n56_), .Y(mai2));
  NO2        g0115(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n138_));
  NA2        g0116(.A(i_6_), .B(new_new_n25_), .Y(new_new_n139_));
  NA2        g0117(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n140_));
  NA4        g0118(.A(new_new_n140_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(mai0));
  AN2        g0119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(i_6_), .Y(new_new_n143_));
  NO2        g0121(.A(i_12_), .B(i_13_), .Y(new_new_n144_));
  NAi21      g0122(.An(i_5_), .B(i_11_), .Y(new_new_n145_));
  NOi21      g0123(.An(new_new_n144_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g0124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NA2        g0125(.A(i_2_), .B(i_3_), .Y(new_new_n148_));
  NO2        g0126(.A(new_new_n148_), .B(i_4_), .Y(new_new_n149_));
  NA2        g0127(.A(new_new_n149_), .B(new_new_n146_), .Y(new_new_n150_));
  AN2        g0128(.A(new_new_n144_), .B(new_new_n83_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(new_new_n27_), .Y(new_new_n152_));
  NA2        g0130(.A(i_1_), .B(i_5_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n73_), .B(new_new_n47_), .Y(new_new_n154_));
  NA2        g0132(.A(new_new_n154_), .B(new_new_n36_), .Y(new_new_n155_));
  NO3        g0133(.A(new_new_n155_), .B(new_new_n153_), .C(new_new_n152_), .Y(new_new_n156_));
  OR2        g0134(.A(i_0_), .B(i_1_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n158_));
  NAi32      g0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NAi21      g0137(.An(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  NOi21      g0138(.An(i_4_), .B(i_10_), .Y(new_new_n161_));
  NA2        g0139(.A(new_new_n161_), .B(new_new_n40_), .Y(new_new_n162_));
  NO2        g0140(.A(i_3_), .B(i_5_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  OAI210     g0143(.A0(new_new_n165_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n166_));
  NO2        g0144(.A(new_new_n166_), .B(new_new_n156_), .Y(new_new_n167_));
  AOI210     g0145(.A0(new_new_n167_), .A1(new_new_n150_), .B0(new_new_n143_), .Y(new_new_n168_));
  NA2        g0146(.A(new_new_n73_), .B(i_1_), .Y(new_new_n169_));
  NA2        g0147(.A(i_3_), .B(new_new_n49_), .Y(new_new_n170_));
  NOi21      g0148(.An(i_4_), .B(i_9_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_11_), .B(i_13_), .Y(new_new_n172_));
  NA2        g0150(.A(new_new_n172_), .B(new_new_n171_), .Y(new_new_n173_));
  OR2        g0151(.A(new_new_n173_), .B(new_new_n170_), .Y(new_new_n174_));
  NO2        g0152(.A(i_4_), .B(i_5_), .Y(new_new_n175_));
  NAi21      g0153(.An(i_12_), .B(i_11_), .Y(new_new_n176_));
  NO2        g0154(.A(new_new_n176_), .B(i_13_), .Y(new_new_n177_));
  NA3        g0155(.A(new_new_n177_), .B(new_new_n175_), .C(new_new_n83_), .Y(new_new_n178_));
  AOI210     g0156(.A0(new_new_n178_), .A1(new_new_n174_), .B0(new_new_n169_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n180_));
  NA2        g0158(.A(new_new_n180_), .B(new_new_n47_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n36_), .B(i_5_), .Y(new_new_n182_));
  NAi31      g0160(.An(new_new_n182_), .B(new_new_n151_), .C(i_11_), .Y(new_new_n183_));
  NA2        g0161(.A(i_3_), .B(i_5_), .Y(new_new_n184_));
  OR2        g0162(.A(new_new_n184_), .B(new_new_n173_), .Y(new_new_n185_));
  AOI210     g0163(.A0(new_new_n185_), .A1(new_new_n183_), .B0(new_new_n181_), .Y(new_new_n186_));
  NO2        g0164(.A(new_new_n73_), .B(i_5_), .Y(new_new_n187_));
  NO2        g0165(.A(i_13_), .B(i_10_), .Y(new_new_n188_));
  NA3        g0166(.A(new_new_n188_), .B(new_new_n187_), .C(new_new_n45_), .Y(new_new_n189_));
  NO2        g0167(.A(i_2_), .B(i_1_), .Y(new_new_n190_));
  NA2        g0168(.A(new_new_n190_), .B(i_3_), .Y(new_new_n191_));
  NAi21      g0169(.An(i_4_), .B(i_12_), .Y(new_new_n192_));
  NO4        g0170(.A(new_new_n192_), .B(new_new_n191_), .C(new_new_n189_), .D(new_new_n25_), .Y(new_new_n193_));
  NO3        g0171(.A(new_new_n193_), .B(new_new_n186_), .C(new_new_n179_), .Y(new_new_n194_));
  INV        g0172(.A(i_8_), .Y(new_new_n195_));
  NA2        g0173(.A(i_8_), .B(i_6_), .Y(new_new_n196_));
  NO3        g0174(.A(i_3_), .B(new_new_n85_), .C(new_new_n49_), .Y(new_new_n197_));
  NA2        g0175(.A(new_new_n197_), .B(new_new_n113_), .Y(new_new_n198_));
  NO3        g0176(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n199_));
  NA3        g0177(.A(new_new_n199_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n200_));
  NO3        g0178(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n201_));
  OAI210     g0179(.A0(new_new_n96_), .A1(i_12_), .B0(new_new_n201_), .Y(new_new_n202_));
  AOI210     g0180(.A0(new_new_n202_), .A1(new_new_n200_), .B0(new_new_n198_), .Y(new_new_n203_));
  NO2        g0181(.A(i_3_), .B(i_8_), .Y(new_new_n204_));
  NO3        g0182(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n205_));
  NA3        g0183(.A(new_new_n205_), .B(new_new_n204_), .C(new_new_n40_), .Y(new_new_n206_));
  NO2        g0184(.A(i_13_), .B(i_9_), .Y(new_new_n207_));
  NA2        g0185(.A(new_new_n207_), .B(i_6_), .Y(new_new_n208_));
  NAi21      g0186(.An(i_12_), .B(i_3_), .Y(new_new_n209_));
  NO2        g0187(.A(new_new_n45_), .B(i_5_), .Y(new_new_n210_));
  NO3        g0188(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n211_));
  NA3        g0189(.A(new_new_n211_), .B(new_new_n210_), .C(i_10_), .Y(new_new_n212_));
  OAI220     g0190(.A0(new_new_n212_), .A1(new_new_n208_), .B0(new_new_n58_), .B1(new_new_n206_), .Y(new_new_n213_));
  AOI210     g0191(.A0(new_new_n213_), .A1(i_7_), .B0(new_new_n203_), .Y(new_new_n214_));
  OAI220     g0192(.A0(new_new_n214_), .A1(i_4_), .B0(new_new_n196_), .B1(new_new_n194_), .Y(new_new_n215_));
  NAi21      g0193(.An(i_12_), .B(i_7_), .Y(new_new_n216_));
  NA3        g0194(.A(i_13_), .B(new_new_n195_), .C(i_10_), .Y(new_new_n217_));
  NO2        g0195(.A(new_new_n217_), .B(new_new_n216_), .Y(new_new_n218_));
  NA2        g0196(.A(i_0_), .B(i_5_), .Y(new_new_n219_));
  OAI220     g0197(.A0(new_new_n85_), .A1(new_new_n191_), .B0(new_new_n181_), .B1(new_new_n134_), .Y(new_new_n220_));
  NAi31      g0198(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n221_));
  NO2        g0199(.A(new_new_n36_), .B(i_13_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n224_));
  NA3        g0202(.A(new_new_n224_), .B(new_new_n223_), .C(new_new_n222_), .Y(new_new_n225_));
  INV        g0203(.A(i_13_), .Y(new_new_n226_));
  NO2        g0204(.A(i_12_), .B(new_new_n226_), .Y(new_new_n227_));
  NA3        g0205(.A(new_new_n227_), .B(new_new_n199_), .C(new_new_n197_), .Y(new_new_n228_));
  OAI210     g0206(.A0(new_new_n225_), .A1(new_new_n221_), .B0(new_new_n228_), .Y(new_new_n229_));
  AOI220     g0207(.A0(new_new_n229_), .A1(new_new_n142_), .B0(new_new_n220_), .B1(new_new_n218_), .Y(new_new_n230_));
  NO2        g0208(.A(i_12_), .B(new_new_n37_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n184_), .B(i_4_), .Y(new_new_n232_));
  NA2        g0210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  OR2        g0211(.A(i_8_), .B(i_7_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n234_), .B(new_new_n85_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n54_), .B(i_1_), .Y(new_new_n236_));
  NA2        g0214(.A(new_new_n236_), .B(new_new_n235_), .Y(new_new_n237_));
  INV        g0215(.A(i_12_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n45_), .B(new_new_n238_), .Y(new_new_n239_));
  NO3        g0217(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n240_));
  NA2        g0218(.A(i_2_), .B(i_1_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n237_), .B(new_new_n233_), .Y(new_new_n242_));
  NO3        g0220(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n243_));
  NAi21      g0221(.An(i_4_), .B(i_3_), .Y(new_new_n244_));
  INV        g0222(.A(new_new_n75_), .Y(new_new_n245_));
  NO2        g0223(.A(i_0_), .B(i_6_), .Y(new_new_n246_));
  NOi41      g0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n247_));
  NA2        g0225(.A(new_new_n247_), .B(new_new_n246_), .Y(new_new_n248_));
  NO2        g0226(.A(new_new_n241_), .B(new_new_n184_), .Y(new_new_n249_));
  NAi21      g0227(.An(new_new_n248_), .B(new_new_n249_), .Y(new_new_n250_));
  INV        g0228(.A(new_new_n250_), .Y(new_new_n251_));
  AOI210     g0229(.A0(new_new_n251_), .A1(new_new_n40_), .B0(new_new_n242_), .Y(new_new_n252_));
  NO2        g0230(.A(i_11_), .B(new_new_n226_), .Y(new_new_n253_));
  NOi21      g0231(.An(i_1_), .B(i_6_), .Y(new_new_n254_));
  NAi21      g0232(.An(i_3_), .B(i_7_), .Y(new_new_n255_));
  NO2        g0233(.A(i_12_), .B(i_3_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n73_), .B(i_5_), .Y(new_new_n257_));
  NAi21      g0235(.An(i_7_), .B(i_10_), .Y(new_new_n258_));
  NA3        g0236(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n259_));
  INV        g0237(.A(new_new_n143_), .Y(new_new_n260_));
  NA2        g0238(.A(new_new_n238_), .B(i_13_), .Y(new_new_n261_));
  NO2        g0239(.A(new_new_n261_), .B(new_new_n75_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n262_), .B(new_new_n260_), .Y(new_new_n263_));
  NO2        g0241(.A(new_new_n234_), .B(new_new_n37_), .Y(new_new_n264_));
  NA2        g0242(.A(i_12_), .B(i_6_), .Y(new_new_n265_));
  OR2        g0243(.A(i_13_), .B(i_9_), .Y(new_new_n266_));
  NO3        g0244(.A(new_new_n266_), .B(new_new_n265_), .C(new_new_n49_), .Y(new_new_n267_));
  NO2        g0245(.A(new_new_n244_), .B(i_2_), .Y(new_new_n268_));
  NA3        g0246(.A(new_new_n268_), .B(new_new_n267_), .C(new_new_n45_), .Y(new_new_n269_));
  NA2        g0247(.A(new_new_n253_), .B(i_9_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n257_), .B(new_new_n64_), .Y(new_new_n271_));
  OAI210     g0249(.A0(new_new_n271_), .A1(new_new_n270_), .B0(new_new_n269_), .Y(new_new_n272_));
  NA2        g0250(.A(new_new_n154_), .B(new_new_n63_), .Y(new_new_n273_));
  NO3        g0251(.A(i_11_), .B(new_new_n226_), .C(new_new_n25_), .Y(new_new_n274_));
  NO2        g0252(.A(new_new_n255_), .B(i_8_), .Y(new_new_n275_));
  NO2        g0253(.A(i_6_), .B(new_new_n49_), .Y(new_new_n276_));
  NA3        g0254(.A(new_new_n276_), .B(new_new_n275_), .C(new_new_n274_), .Y(new_new_n277_));
  NO3        g0255(.A(new_new_n26_), .B(new_new_n85_), .C(i_5_), .Y(new_new_n278_));
  NA3        g0256(.A(new_new_n278_), .B(new_new_n264_), .C(new_new_n227_), .Y(new_new_n279_));
  AOI210     g0257(.A0(new_new_n279_), .A1(new_new_n277_), .B0(new_new_n273_), .Y(new_new_n280_));
  AOI210     g0258(.A0(new_new_n272_), .A1(new_new_n264_), .B0(new_new_n280_), .Y(new_new_n281_));
  NA4        g0259(.A(new_new_n281_), .B(new_new_n263_), .C(new_new_n252_), .D(new_new_n230_), .Y(new_new_n282_));
  NO3        g0260(.A(i_12_), .B(new_new_n226_), .C(new_new_n37_), .Y(new_new_n283_));
  INV        g0261(.A(new_new_n283_), .Y(new_new_n284_));
  NA2        g0262(.A(i_8_), .B(new_new_n101_), .Y(new_new_n285_));
  NO3        g0263(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n286_));
  AOI220     g0264(.A0(new_new_n286_), .A1(new_new_n197_), .B0(new_new_n163_), .B1(new_new_n236_), .Y(new_new_n287_));
  NO2        g0265(.A(new_new_n287_), .B(new_new_n285_), .Y(new_new_n288_));
  NO2        g0266(.A(new_new_n241_), .B(i_0_), .Y(new_new_n289_));
  AOI220     g0267(.A0(new_new_n289_), .A1(i_8_), .B0(i_1_), .B1(new_new_n142_), .Y(new_new_n290_));
  NA2        g0268(.A(new_new_n276_), .B(new_new_n26_), .Y(new_new_n291_));
  NO2        g0269(.A(new_new_n291_), .B(new_new_n290_), .Y(new_new_n292_));
  NA2        g0270(.A(i_0_), .B(i_1_), .Y(new_new_n293_));
  NO2        g0271(.A(new_new_n293_), .B(i_2_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n59_), .B(i_6_), .Y(new_new_n295_));
  NA3        g0273(.A(new_new_n295_), .B(new_new_n294_), .C(new_new_n163_), .Y(new_new_n296_));
  OAI210     g0274(.A0(new_new_n165_), .A1(new_new_n143_), .B0(new_new_n296_), .Y(new_new_n297_));
  NO3        g0275(.A(new_new_n297_), .B(new_new_n292_), .C(new_new_n288_), .Y(new_new_n298_));
  NO2        g0276(.A(i_3_), .B(i_10_), .Y(new_new_n299_));
  NA3        g0277(.A(new_new_n299_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n300_));
  NO2        g0278(.A(i_2_), .B(new_new_n101_), .Y(new_new_n301_));
  NA2        g0279(.A(i_1_), .B(new_new_n36_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n302_), .B(i_8_), .Y(new_new_n303_));
  NA2        g0281(.A(new_new_n303_), .B(new_new_n301_), .Y(new_new_n304_));
  AN2        g0282(.A(i_3_), .B(i_10_), .Y(new_new_n305_));
  NA4        g0283(.A(new_new_n305_), .B(new_new_n199_), .C(new_new_n177_), .D(new_new_n175_), .Y(new_new_n306_));
  NO2        g0284(.A(i_5_), .B(new_new_n37_), .Y(new_new_n307_));
  NO2        g0285(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n308_));
  OR2        g0286(.A(new_new_n304_), .B(new_new_n300_), .Y(new_new_n309_));
  OAI220     g0287(.A0(new_new_n309_), .A1(i_6_), .B0(new_new_n298_), .B1(new_new_n284_), .Y(new_new_n310_));
  NO4        g0288(.A(new_new_n310_), .B(new_new_n282_), .C(new_new_n215_), .D(new_new_n168_), .Y(new_new_n311_));
  NO3        g0289(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n312_));
  NO2        g0290(.A(new_new_n59_), .B(new_new_n85_), .Y(new_new_n313_));
  NO3        g0291(.A(i_6_), .B(new_new_n195_), .C(i_7_), .Y(new_new_n314_));
  NA2        g0292(.A(new_new_n314_), .B(new_new_n199_), .Y(new_new_n315_));
  INV        g0293(.A(new_new_n315_), .Y(new_new_n316_));
  NO2        g0294(.A(i_2_), .B(i_3_), .Y(new_new_n317_));
  OR2        g0295(.A(i_0_), .B(i_5_), .Y(new_new_n318_));
  NA3        g0296(.A(new_new_n235_), .B(new_new_n317_), .C(i_1_), .Y(new_new_n319_));
  NA3        g0297(.A(new_new_n289_), .B(new_new_n163_), .C(new_new_n113_), .Y(new_new_n320_));
  NAi21      g0298(.An(i_8_), .B(i_7_), .Y(new_new_n321_));
  NO2        g0299(.A(new_new_n321_), .B(i_6_), .Y(new_new_n322_));
  NO2        g0300(.A(new_new_n157_), .B(new_new_n47_), .Y(new_new_n323_));
  NA3        g0301(.A(new_new_n323_), .B(new_new_n322_), .C(new_new_n163_), .Y(new_new_n324_));
  NA3        g0302(.A(new_new_n324_), .B(new_new_n320_), .C(new_new_n319_), .Y(new_new_n325_));
  OAI210     g0303(.A0(new_new_n325_), .A1(new_new_n316_), .B0(i_4_), .Y(new_new_n326_));
  NO2        g0304(.A(i_12_), .B(i_10_), .Y(new_new_n327_));
  NOi21      g0305(.An(i_5_), .B(i_0_), .Y(new_new_n328_));
  NO3        g0306(.A(new_new_n302_), .B(new_new_n328_), .C(new_new_n129_), .Y(new_new_n329_));
  NA4        g0307(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n85_), .D(i_8_), .Y(new_new_n330_));
  NA2        g0308(.A(new_new_n329_), .B(new_new_n327_), .Y(new_new_n331_));
  NO2        g0309(.A(i_6_), .B(i_8_), .Y(new_new_n332_));
  NOi21      g0310(.An(i_0_), .B(i_2_), .Y(new_new_n333_));
  AN2        g0311(.A(new_new_n333_), .B(new_new_n332_), .Y(new_new_n334_));
  NO2        g0312(.A(i_1_), .B(i_7_), .Y(new_new_n335_));
  AO220      g0313(.A0(new_new_n335_), .A1(new_new_n334_), .B0(new_new_n322_), .B1(new_new_n236_), .Y(new_new_n336_));
  NA2        g0314(.A(new_new_n336_), .B(new_new_n42_), .Y(new_new_n337_));
  NA3        g0315(.A(new_new_n337_), .B(new_new_n331_), .C(new_new_n326_), .Y(new_new_n338_));
  NO3        g0316(.A(new_new_n234_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n339_));
  NO3        g0317(.A(new_new_n321_), .B(i_2_), .C(i_1_), .Y(new_new_n340_));
  OAI210     g0318(.A0(new_new_n340_), .A1(new_new_n339_), .B0(i_6_), .Y(new_new_n341_));
  NA2        g0319(.A(new_new_n254_), .B(new_new_n301_), .Y(new_new_n342_));
  NA2        g0320(.A(new_new_n342_), .B(new_new_n341_), .Y(new_new_n343_));
  NA2        g0321(.A(new_new_n343_), .B(i_3_), .Y(new_new_n344_));
  INV        g0322(.A(new_new_n84_), .Y(new_new_n345_));
  NO2        g0323(.A(new_new_n293_), .B(new_new_n81_), .Y(new_new_n346_));
  NA2        g0324(.A(new_new_n346_), .B(new_new_n133_), .Y(new_new_n347_));
  NO2        g0325(.A(new_new_n92_), .B(new_new_n195_), .Y(new_new_n348_));
  NA2        g0326(.A(new_new_n348_), .B(new_new_n63_), .Y(new_new_n349_));
  AOI210     g0327(.A0(new_new_n349_), .A1(new_new_n347_), .B0(new_new_n345_), .Y(new_new_n350_));
  NO2        g0328(.A(new_new_n195_), .B(i_9_), .Y(new_new_n351_));
  NA2        g0329(.A(new_new_n351_), .B(i_6_), .Y(new_new_n352_));
  NO2        g0330(.A(new_new_n350_), .B(new_new_n292_), .Y(new_new_n353_));
  AOI210     g0331(.A0(new_new_n353_), .A1(new_new_n344_), .B0(new_new_n162_), .Y(new_new_n354_));
  AOI210     g0332(.A0(new_new_n338_), .A1(new_new_n312_), .B0(new_new_n354_), .Y(new_new_n355_));
  NOi32      g0333(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n356_));
  INV        g0334(.A(new_new_n356_), .Y(new_new_n357_));
  NAi21      g0335(.An(i_0_), .B(i_6_), .Y(new_new_n358_));
  NAi21      g0336(.An(i_1_), .B(i_5_), .Y(new_new_n359_));
  NA2        g0337(.A(new_new_n359_), .B(new_new_n358_), .Y(new_new_n360_));
  NA2        g0338(.A(new_new_n360_), .B(new_new_n25_), .Y(new_new_n361_));
  OAI210     g0339(.A0(new_new_n361_), .A1(new_new_n159_), .B0(new_new_n248_), .Y(new_new_n362_));
  NAi41      g0340(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n363_));
  OAI220     g0341(.A0(new_new_n363_), .A1(new_new_n359_), .B0(new_new_n221_), .B1(new_new_n159_), .Y(new_new_n364_));
  AOI210     g0342(.A0(new_new_n363_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n365_));
  NOi32      g0343(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n366_));
  NAi21      g0344(.An(i_6_), .B(i_1_), .Y(new_new_n367_));
  NA3        g0345(.A(new_new_n367_), .B(new_new_n366_), .C(new_new_n47_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n368_), .B(i_0_), .Y(new_new_n369_));
  OR3        g0347(.A(new_new_n369_), .B(new_new_n365_), .C(new_new_n364_), .Y(new_new_n370_));
  NO2        g0348(.A(i_1_), .B(new_new_n101_), .Y(new_new_n371_));
  NAi21      g0349(.An(i_3_), .B(i_4_), .Y(new_new_n372_));
  NA2        g0350(.A(i_2_), .B(i_7_), .Y(new_new_n373_));
  NO2        g0351(.A(new_new_n372_), .B(i_10_), .Y(new_new_n374_));
  AOI210     g0352(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n375_));
  OAI210     g0353(.A0(new_new_n375_), .A1(new_new_n190_), .B0(new_new_n374_), .Y(new_new_n376_));
  AOI220     g0354(.A0(new_new_n374_), .A1(new_new_n335_), .B0(new_new_n240_), .B1(new_new_n190_), .Y(new_new_n377_));
  AOI210     g0355(.A0(new_new_n377_), .A1(new_new_n376_), .B0(i_5_), .Y(new_new_n378_));
  NO3        g0356(.A(new_new_n378_), .B(new_new_n370_), .C(new_new_n362_), .Y(new_new_n379_));
  NO2        g0357(.A(new_new_n379_), .B(new_new_n357_), .Y(new_new_n380_));
  NO2        g0358(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n381_));
  AN2        g0359(.A(i_12_), .B(i_5_), .Y(new_new_n382_));
  NA2        g0360(.A(i_3_), .B(new_new_n382_), .Y(new_new_n383_));
  NO2        g0361(.A(i_11_), .B(i_6_), .Y(new_new_n384_));
  NA3        g0362(.A(new_new_n384_), .B(new_new_n323_), .C(new_new_n226_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n385_), .B(new_new_n383_), .Y(new_new_n386_));
  NO2        g0364(.A(new_new_n244_), .B(i_5_), .Y(new_new_n387_));
  NO2        g0365(.A(i_5_), .B(i_10_), .Y(new_new_n388_));
  AOI220     g0366(.A0(new_new_n388_), .A1(new_new_n268_), .B0(new_new_n387_), .B1(new_new_n199_), .Y(new_new_n389_));
  NA2        g0367(.A(new_new_n144_), .B(new_new_n46_), .Y(new_new_n390_));
  NO2        g0368(.A(new_new_n390_), .B(new_new_n389_), .Y(new_new_n391_));
  OAI210     g0369(.A0(new_new_n391_), .A1(new_new_n386_), .B0(new_new_n381_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n393_));
  NA2        g0371(.A(new_new_n386_), .B(new_new_n393_), .Y(new_new_n394_));
  NO3        g0372(.A(new_new_n85_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n299_), .B(new_new_n90_), .Y(new_new_n396_));
  NO2        g0374(.A(i_11_), .B(i_12_), .Y(new_new_n397_));
  NA2        g0375(.A(new_new_n397_), .B(new_new_n36_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n396_), .B(new_new_n398_), .Y(new_new_n399_));
  NA2        g0377(.A(new_new_n388_), .B(new_new_n238_), .Y(new_new_n400_));
  NA2        g0378(.A(new_new_n42_), .B(i_11_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n401_), .B(new_new_n221_), .Y(new_new_n402_));
  NAi21      g0380(.An(i_13_), .B(i_0_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n403_), .B(new_new_n241_), .Y(new_new_n404_));
  OAI210     g0382(.A0(new_new_n402_), .A1(new_new_n399_), .B0(new_new_n404_), .Y(new_new_n405_));
  NA3        g0383(.A(new_new_n405_), .B(new_new_n394_), .C(new_new_n392_), .Y(new_new_n406_));
  NA2        g0384(.A(new_new_n45_), .B(new_new_n226_), .Y(new_new_n407_));
  NO2        g0385(.A(i_0_), .B(i_11_), .Y(new_new_n408_));
  AN2        g0386(.A(i_1_), .B(i_6_), .Y(new_new_n409_));
  NOi21      g0387(.An(i_2_), .B(i_12_), .Y(new_new_n410_));
  NA2        g0388(.A(new_new_n410_), .B(new_new_n409_), .Y(new_new_n411_));
  INV        g0389(.A(new_new_n411_), .Y(new_new_n412_));
  NA2        g0390(.A(new_new_n142_), .B(i_9_), .Y(new_new_n413_));
  NO2        g0391(.A(new_new_n413_), .B(i_4_), .Y(new_new_n414_));
  NA2        g0392(.A(new_new_n412_), .B(new_new_n414_), .Y(new_new_n415_));
  NAi21      g0393(.An(i_9_), .B(i_4_), .Y(new_new_n416_));
  OR2        g0394(.A(i_13_), .B(i_10_), .Y(new_new_n417_));
  NO3        g0395(.A(new_new_n417_), .B(new_new_n118_), .C(new_new_n416_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n173_), .B(new_new_n124_), .Y(new_new_n419_));
  OR2        g0397(.A(new_new_n217_), .B(new_new_n216_), .Y(new_new_n420_));
  NO2        g0398(.A(new_new_n101_), .B(new_new_n25_), .Y(new_new_n421_));
  NA2        g0399(.A(new_new_n276_), .B(new_new_n211_), .Y(new_new_n422_));
  NO2        g0400(.A(new_new_n422_), .B(new_new_n420_), .Y(new_new_n423_));
  INV        g0401(.A(new_new_n423_), .Y(new_new_n424_));
  AOI210     g0402(.A0(new_new_n424_), .A1(new_new_n415_), .B0(new_new_n26_), .Y(new_new_n425_));
  NA2        g0403(.A(new_new_n320_), .B(new_new_n319_), .Y(new_new_n426_));
  AOI220     g0404(.A0(new_new_n295_), .A1(new_new_n286_), .B0(new_new_n289_), .B1(new_new_n313_), .Y(new_new_n427_));
  NO2        g0405(.A(new_new_n427_), .B(new_new_n170_), .Y(new_new_n428_));
  NO2        g0406(.A(new_new_n184_), .B(new_new_n85_), .Y(new_new_n429_));
  AOI220     g0407(.A0(new_new_n429_), .A1(new_new_n294_), .B0(new_new_n278_), .B1(new_new_n211_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n430_), .B(new_new_n285_), .Y(new_new_n431_));
  NO3        g0409(.A(new_new_n431_), .B(new_new_n428_), .C(new_new_n426_), .Y(new_new_n432_));
  NA2        g0410(.A(new_new_n197_), .B(new_new_n96_), .Y(new_new_n433_));
  NA3        g0411(.A(new_new_n323_), .B(new_new_n163_), .C(new_new_n85_), .Y(new_new_n434_));
  AOI210     g0412(.A0(new_new_n434_), .A1(new_new_n433_), .B0(new_new_n321_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n295_), .B(new_new_n236_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n436_), .B(new_new_n184_), .Y(new_new_n437_));
  NO2        g0415(.A(i_3_), .B(new_new_n49_), .Y(new_new_n438_));
  NA3        g0416(.A(new_new_n335_), .B(new_new_n334_), .C(new_new_n438_), .Y(new_new_n439_));
  INV        g0417(.A(new_new_n314_), .Y(new_new_n440_));
  OAI210     g0418(.A0(new_new_n440_), .A1(new_new_n191_), .B0(new_new_n439_), .Y(new_new_n441_));
  NO3        g0419(.A(new_new_n441_), .B(new_new_n437_), .C(new_new_n435_), .Y(new_new_n442_));
  AOI210     g0420(.A0(new_new_n442_), .A1(new_new_n432_), .B0(new_new_n270_), .Y(new_new_n443_));
  NO4        g0421(.A(new_new_n443_), .B(new_new_n425_), .C(new_new_n406_), .D(new_new_n380_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n73_), .B(i_13_), .Y(new_new_n445_));
  NO2        g0423(.A(i_10_), .B(i_9_), .Y(new_new_n446_));
  NAi21      g0424(.An(i_12_), .B(i_8_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n447_), .B(i_3_), .Y(new_new_n448_));
  NO2        g0426(.A(new_new_n47_), .B(i_4_), .Y(new_new_n449_));
  NA2        g0427(.A(new_new_n449_), .B(new_new_n104_), .Y(new_new_n450_));
  NO2        g0428(.A(new_new_n450_), .B(new_new_n206_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n308_), .B(i_0_), .Y(new_new_n452_));
  NO3        g0430(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n453_));
  NA2        g0431(.A(new_new_n265_), .B(new_new_n97_), .Y(new_new_n454_));
  NA2        g0432(.A(new_new_n454_), .B(new_new_n453_), .Y(new_new_n455_));
  NA2        g0433(.A(i_8_), .B(i_9_), .Y(new_new_n456_));
  NO2        g0434(.A(new_new_n455_), .B(new_new_n452_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n253_), .B(new_new_n307_), .Y(new_new_n458_));
  NO3        g0436(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n459_));
  INV        g0437(.A(new_new_n459_), .Y(new_new_n460_));
  NA3        g0438(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n461_));
  NA4        g0439(.A(new_new_n145_), .B(new_new_n116_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n462_));
  OAI220     g0440(.A0(new_new_n462_), .A1(new_new_n461_), .B0(new_new_n460_), .B1(new_new_n458_), .Y(new_new_n463_));
  NO3        g0441(.A(new_new_n463_), .B(new_new_n457_), .C(new_new_n451_), .Y(new_new_n464_));
  OR2        g0442(.A(new_new_n293_), .B(new_new_n208_), .Y(new_new_n465_));
  OA210      g0443(.A0(new_new_n352_), .A1(new_new_n101_), .B0(new_new_n296_), .Y(new_new_n466_));
  OA220      g0444(.A0(new_new_n466_), .A1(new_new_n162_), .B0(new_new_n465_), .B1(new_new_n233_), .Y(new_new_n467_));
  NA2        g0445(.A(new_new_n96_), .B(i_13_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n429_), .B(new_new_n381_), .Y(new_new_n469_));
  NO2        g0447(.A(i_2_), .B(i_13_), .Y(new_new_n470_));
  NA3        g0448(.A(new_new_n470_), .B(new_new_n161_), .C(new_new_n99_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n469_), .B(new_new_n468_), .Y(new_new_n472_));
  NO3        g0450(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n473_));
  NO2        g0451(.A(i_6_), .B(i_7_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n474_), .B(new_new_n473_), .Y(new_new_n475_));
  NO2        g0453(.A(i_11_), .B(i_1_), .Y(new_new_n476_));
  OR2        g0454(.A(i_11_), .B(i_8_), .Y(new_new_n477_));
  NOi21      g0455(.An(i_2_), .B(i_7_), .Y(new_new_n478_));
  NAi31      g0456(.An(new_new_n477_), .B(new_new_n478_), .C(i_0_), .Y(new_new_n479_));
  NO2        g0457(.A(new_new_n417_), .B(i_6_), .Y(new_new_n480_));
  NA2        g0458(.A(new_new_n480_), .B(i_1_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n481_), .B(new_new_n479_), .Y(new_new_n482_));
  NO2        g0460(.A(i_3_), .B(new_new_n195_), .Y(new_new_n483_));
  NO2        g0461(.A(i_6_), .B(i_10_), .Y(new_new_n484_));
  NA4        g0462(.A(new_new_n484_), .B(new_new_n312_), .C(new_new_n483_), .D(new_new_n238_), .Y(new_new_n485_));
  NO2        g0463(.A(new_new_n485_), .B(new_new_n155_), .Y(new_new_n486_));
  NA2        g0464(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n487_));
  NO2        g0465(.A(new_new_n157_), .B(i_3_), .Y(new_new_n488_));
  NAi31      g0466(.An(new_new_n487_), .B(new_new_n488_), .C(new_new_n227_), .Y(new_new_n489_));
  NA3        g0467(.A(new_new_n393_), .B(new_new_n180_), .C(new_new_n149_), .Y(new_new_n490_));
  NA2        g0468(.A(new_new_n490_), .B(new_new_n489_), .Y(new_new_n491_));
  NO4        g0469(.A(new_new_n491_), .B(new_new_n486_), .C(new_new_n482_), .D(new_new_n472_), .Y(new_new_n492_));
  NA2        g0470(.A(new_new_n453_), .B(new_new_n382_), .Y(new_new_n493_));
  NAi21      g0471(.An(new_new_n217_), .B(new_new_n397_), .Y(new_new_n494_));
  NA2        g0472(.A(new_new_n335_), .B(new_new_n219_), .Y(new_new_n495_));
  NA3        g0473(.A(i_6_), .B(i_3_), .C(new_new_n142_), .Y(new_new_n496_));
  OR3        g0474(.A(new_new_n302_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n497_));
  OAI220     g0475(.A0(new_new_n497_), .A1(new_new_n496_), .B0(new_new_n495_), .B1(new_new_n494_), .Y(new_new_n498_));
  NA3        g0476(.A(new_new_n305_), .B(new_new_n224_), .C(new_new_n73_), .Y(new_new_n499_));
  NO2        g0477(.A(new_new_n499_), .B(new_new_n475_), .Y(new_new_n500_));
  NO2        g0478(.A(new_new_n500_), .B(new_new_n498_), .Y(new_new_n501_));
  NA4        g0479(.A(new_new_n501_), .B(new_new_n492_), .C(new_new_n467_), .D(new_new_n464_), .Y(new_new_n502_));
  NA3        g0480(.A(new_new_n305_), .B(new_new_n177_), .C(new_new_n175_), .Y(new_new_n503_));
  INV        g0481(.A(new_new_n503_), .Y(new_new_n504_));
  BUFFER     g0482(.A(new_new_n286_), .Y(new_new_n505_));
  NA2        g0483(.A(new_new_n505_), .B(new_new_n504_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n123_), .B(new_new_n112_), .Y(new_new_n507_));
  AO220      g0485(.A0(new_new_n507_), .A1(new_new_n453_), .B0(new_new_n418_), .B1(i_6_), .Y(new_new_n508_));
  NA2        g0486(.A(new_new_n312_), .B(new_new_n164_), .Y(new_new_n509_));
  OAI210     g0487(.A0(new_new_n509_), .A1(new_new_n233_), .B0(new_new_n306_), .Y(new_new_n510_));
  AOI220     g0488(.A0(new_new_n510_), .A1(new_new_n322_), .B0(new_new_n508_), .B1(new_new_n308_), .Y(new_new_n511_));
  NA2        g0489(.A(new_new_n356_), .B(new_new_n73_), .Y(new_new_n512_));
  NO2        g0490(.A(new_new_n36_), .B(i_8_), .Y(new_new_n513_));
  AOI210     g0491(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n418_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n257_), .B(new_new_n64_), .Y(new_new_n515_));
  OAI210     g0493(.A0(i_8_), .A1(new_new_n515_), .B0(new_new_n134_), .Y(new_new_n516_));
  NO2        g0494(.A(i_7_), .B(new_new_n200_), .Y(new_new_n517_));
  OR2        g0495(.A(new_new_n184_), .B(i_4_), .Y(new_new_n518_));
  NO2        g0496(.A(new_new_n518_), .B(new_new_n85_), .Y(new_new_n519_));
  AOI220     g0497(.A0(new_new_n519_), .A1(new_new_n517_), .B0(new_new_n516_), .B1(new_new_n419_), .Y(new_new_n520_));
  NA4        g0498(.A(new_new_n520_), .B(new_new_n514_), .C(new_new_n511_), .D(new_new_n506_), .Y(new_new_n521_));
  NA2        g0499(.A(new_new_n387_), .B(new_new_n294_), .Y(new_new_n522_));
  OAI210     g0500(.A0(new_new_n383_), .A1(new_new_n169_), .B0(new_new_n522_), .Y(new_new_n523_));
  NA2        g0501(.A(new_new_n1026_), .B(new_new_n226_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n484_), .B(new_new_n27_), .Y(new_new_n525_));
  NO2        g0503(.A(new_new_n525_), .B(new_new_n524_), .Y(new_new_n526_));
  NOi31      g0504(.An(new_new_n314_), .B(new_new_n417_), .C(new_new_n38_), .Y(new_new_n527_));
  OAI210     g0505(.A0(new_new_n527_), .A1(new_new_n526_), .B0(new_new_n523_), .Y(new_new_n528_));
  NO2        g0506(.A(i_8_), .B(i_7_), .Y(new_new_n529_));
  OAI210     g0507(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n530_));
  NA2        g0508(.A(new_new_n530_), .B(new_new_n224_), .Y(new_new_n531_));
  OAI220     g0509(.A0(new_new_n47_), .A1(new_new_n518_), .B0(new_new_n531_), .B1(new_new_n244_), .Y(new_new_n532_));
  NA2        g0510(.A(new_new_n45_), .B(i_10_), .Y(new_new_n533_));
  NO2        g0511(.A(new_new_n533_), .B(i_6_), .Y(new_new_n534_));
  NA3        g0512(.A(new_new_n534_), .B(new_new_n532_), .C(new_new_n529_), .Y(new_new_n535_));
  AOI220     g0513(.A0(new_new_n429_), .A1(new_new_n323_), .B0(new_new_n249_), .B1(new_new_n246_), .Y(new_new_n536_));
  OAI220     g0514(.A0(new_new_n536_), .A1(new_new_n261_), .B0(new_new_n468_), .B1(new_new_n134_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n537_), .B(new_new_n264_), .Y(new_new_n538_));
  NOi31      g0516(.An(new_new_n289_), .B(new_new_n300_), .C(new_new_n182_), .Y(new_new_n539_));
  NA3        g0517(.A(new_new_n305_), .B(new_new_n175_), .C(new_new_n96_), .Y(new_new_n540_));
  NO2        g0518(.A(new_new_n222_), .B(new_new_n45_), .Y(new_new_n541_));
  NO2        g0519(.A(new_new_n157_), .B(i_5_), .Y(new_new_n542_));
  NA3        g0520(.A(new_new_n542_), .B(new_new_n407_), .C(new_new_n317_), .Y(new_new_n543_));
  OAI210     g0521(.A0(new_new_n543_), .A1(new_new_n541_), .B0(new_new_n540_), .Y(new_new_n544_));
  OAI210     g0522(.A0(new_new_n544_), .A1(new_new_n539_), .B0(new_new_n459_), .Y(new_new_n545_));
  NA4        g0523(.A(new_new_n545_), .B(new_new_n538_), .C(new_new_n535_), .D(new_new_n528_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n283_), .B(new_new_n84_), .Y(new_new_n547_));
  NO2        g0525(.A(new_new_n347_), .B(new_new_n547_), .Y(new_new_n548_));
  NA2        g0526(.A(new_new_n295_), .B(new_new_n286_), .Y(new_new_n549_));
  NO2        g0527(.A(new_new_n549_), .B(new_new_n174_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n551_));
  NA2        g0529(.A(new_new_n446_), .B(new_new_n222_), .Y(new_new_n552_));
  NO2        g0530(.A(new_new_n551_), .B(new_new_n552_), .Y(new_new_n553_));
  NO3        g0531(.A(new_new_n553_), .B(new_new_n550_), .C(new_new_n548_), .Y(new_new_n554_));
  NO4        g0532(.A(new_new_n254_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n555_));
  NO3        g0533(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n556_));
  NO2        g0534(.A(new_new_n234_), .B(new_new_n36_), .Y(new_new_n557_));
  AN2        g0535(.A(new_new_n557_), .B(new_new_n556_), .Y(new_new_n558_));
  OA210      g0536(.A0(new_new_n558_), .A1(new_new_n555_), .B0(new_new_n356_), .Y(new_new_n559_));
  NO2        g0537(.A(new_new_n417_), .B(i_1_), .Y(new_new_n560_));
  NOi31      g0538(.An(new_new_n560_), .B(new_new_n454_), .C(new_new_n73_), .Y(new_new_n561_));
  AN4        g0539(.A(new_new_n561_), .B(new_new_n414_), .C(i_3_), .D(i_2_), .Y(new_new_n562_));
  NO2        g0540(.A(new_new_n427_), .B(new_new_n178_), .Y(new_new_n563_));
  NO3        g0541(.A(new_new_n563_), .B(new_new_n562_), .C(new_new_n559_), .Y(new_new_n564_));
  NOi21      g0542(.An(i_10_), .B(i_6_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n566_));
  AOI220     g0544(.A0(new_new_n283_), .A1(new_new_n566_), .B0(new_new_n274_), .B1(new_new_n565_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n567_), .B(new_new_n452_), .Y(new_new_n568_));
  NO2        g0546(.A(new_new_n115_), .B(new_new_n23_), .Y(new_new_n569_));
  NA2        g0547(.A(new_new_n314_), .B(new_new_n164_), .Y(new_new_n570_));
  AOI220     g0548(.A0(new_new_n570_), .A1(new_new_n436_), .B0(new_new_n185_), .B1(new_new_n183_), .Y(new_new_n571_));
  NOi21      g0549(.An(new_new_n146_), .B(new_new_n330_), .Y(new_new_n572_));
  NO3        g0550(.A(new_new_n572_), .B(new_new_n571_), .C(new_new_n568_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n512_), .B(new_new_n377_), .Y(new_new_n574_));
  INV        g0552(.A(new_new_n317_), .Y(new_new_n575_));
  NO2        g0553(.A(i_12_), .B(new_new_n85_), .Y(new_new_n576_));
  NA3        g0554(.A(new_new_n576_), .B(new_new_n274_), .C(i_5_), .Y(new_new_n577_));
  NA3        g0555(.A(new_new_n384_), .B(new_new_n283_), .C(new_new_n219_), .Y(new_new_n578_));
  AOI210     g0556(.A0(new_new_n578_), .A1(new_new_n577_), .B0(new_new_n575_), .Y(new_new_n579_));
  NO3        g0557(.A(i_4_), .B(new_new_n341_), .C(new_new_n300_), .Y(new_new_n580_));
  NO3        g0558(.A(new_new_n580_), .B(new_new_n579_), .C(new_new_n574_), .Y(new_new_n581_));
  NA4        g0559(.A(new_new_n581_), .B(new_new_n573_), .C(new_new_n564_), .D(new_new_n554_), .Y(new_new_n582_));
  NO4        g0560(.A(new_new_n582_), .B(new_new_n546_), .C(new_new_n521_), .D(new_new_n502_), .Y(new_new_n583_));
  NA4        g0561(.A(new_new_n583_), .B(new_new_n444_), .C(new_new_n355_), .D(new_new_n311_), .Y(mai7));
  NO2        g0562(.A(new_new_n92_), .B(new_new_n55_), .Y(new_new_n585_));
  NO2        g0563(.A(new_new_n108_), .B(new_new_n89_), .Y(new_new_n586_));
  NA2        g0564(.A(i_3_), .B(new_new_n586_), .Y(new_new_n587_));
  NA2        g0565(.A(i_11_), .B(new_new_n195_), .Y(new_new_n588_));
  INV        g0566(.A(new_new_n587_), .Y(new_new_n589_));
  NA3        g0567(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n590_));
  NO2        g0568(.A(new_new_n238_), .B(i_4_), .Y(new_new_n591_));
  NA2        g0569(.A(new_new_n591_), .B(i_8_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n105_), .B(new_new_n590_), .Y(new_new_n593_));
  NA2        g0571(.A(i_2_), .B(new_new_n85_), .Y(new_new_n594_));
  OAI210     g0572(.A0(new_new_n88_), .A1(new_new_n204_), .B0(new_new_n205_), .Y(new_new_n595_));
  NO2        g0573(.A(i_7_), .B(new_new_n37_), .Y(new_new_n596_));
  NA2        g0574(.A(i_4_), .B(i_8_), .Y(new_new_n597_));
  AOI210     g0575(.A0(new_new_n597_), .A1(new_new_n305_), .B0(new_new_n596_), .Y(new_new_n598_));
  OAI220     g0576(.A0(new_new_n598_), .A1(new_new_n594_), .B0(new_new_n595_), .B1(i_13_), .Y(new_new_n599_));
  NO4        g0577(.A(new_new_n599_), .B(new_new_n593_), .C(new_new_n589_), .D(new_new_n585_), .Y(new_new_n600_));
  AOI210     g0578(.A0(new_new_n129_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n601_));
  AOI210     g0579(.A0(new_new_n601_), .A1(new_new_n238_), .B0(new_new_n161_), .Y(new_new_n602_));
  OR2        g0580(.A(i_6_), .B(i_10_), .Y(new_new_n603_));
  NO2        g0581(.A(new_new_n603_), .B(new_new_n23_), .Y(new_new_n604_));
  OR3        g0582(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n605_));
  NO3        g0583(.A(new_new_n605_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n606_));
  INV        g0584(.A(new_new_n201_), .Y(new_new_n607_));
  NO2        g0585(.A(new_new_n606_), .B(new_new_n604_), .Y(new_new_n608_));
  OA220      g0586(.A0(new_new_n608_), .A1(new_new_n575_), .B0(new_new_n602_), .B1(new_new_n266_), .Y(new_new_n609_));
  AOI210     g0587(.A0(new_new_n609_), .A1(new_new_n600_), .B0(new_new_n63_), .Y(new_new_n610_));
  NOi21      g0588(.An(i_11_), .B(i_7_), .Y(new_new_n611_));
  AO210      g0589(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n612_));
  NO2        g0590(.A(new_new_n612_), .B(new_new_n611_), .Y(new_new_n613_));
  NA2        g0591(.A(new_new_n613_), .B(new_new_n207_), .Y(new_new_n614_));
  NA3        g0592(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n615_));
  NAi31      g0593(.An(new_new_n615_), .B(new_new_n216_), .C(i_11_), .Y(new_new_n616_));
  AOI210     g0594(.A0(new_new_n616_), .A1(new_new_n614_), .B0(new_new_n63_), .Y(new_new_n617_));
  NA2        g0595(.A(new_new_n87_), .B(new_new_n63_), .Y(new_new_n618_));
  AO210      g0596(.A0(new_new_n618_), .A1(new_new_n377_), .B0(new_new_n41_), .Y(new_new_n619_));
  NO3        g0597(.A(new_new_n258_), .B(new_new_n209_), .C(new_new_n588_), .Y(new_new_n620_));
  OAI210     g0598(.A0(new_new_n620_), .A1(new_new_n227_), .B0(new_new_n63_), .Y(new_new_n621_));
  NA2        g0599(.A(new_new_n410_), .B(new_new_n31_), .Y(new_new_n622_));
  OR2        g0600(.A(new_new_n209_), .B(new_new_n108_), .Y(new_new_n623_));
  NA2        g0601(.A(new_new_n623_), .B(new_new_n622_), .Y(new_new_n624_));
  NO2        g0602(.A(new_new_n63_), .B(i_9_), .Y(new_new_n625_));
  NO2        g0603(.A(new_new_n625_), .B(i_4_), .Y(new_new_n626_));
  NA2        g0604(.A(new_new_n626_), .B(new_new_n624_), .Y(new_new_n627_));
  NO2        g0605(.A(i_1_), .B(i_12_), .Y(new_new_n628_));
  NA3        g0606(.A(new_new_n628_), .B(new_new_n110_), .C(new_new_n24_), .Y(new_new_n629_));
  NA4        g0607(.A(new_new_n629_), .B(new_new_n627_), .C(new_new_n621_), .D(new_new_n619_), .Y(new_new_n630_));
  OAI210     g0608(.A0(new_new_n630_), .A1(new_new_n617_), .B0(i_6_), .Y(new_new_n631_));
  NO2        g0609(.A(i_6_), .B(i_11_), .Y(new_new_n632_));
  INV        g0610(.A(new_new_n455_), .Y(new_new_n633_));
  NO4        g0611(.A(new_new_n216_), .B(new_new_n129_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n634_));
  NA2        g0612(.A(new_new_n634_), .B(new_new_n625_), .Y(new_new_n635_));
  INV        g0613(.A(new_new_n635_), .Y(new_new_n636_));
  NA3        g0614(.A(new_new_n529_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n637_));
  NA2        g0615(.A(new_new_n138_), .B(i_9_), .Y(new_new_n638_));
  NA3        g0616(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n639_));
  NO2        g0617(.A(new_new_n47_), .B(i_1_), .Y(new_new_n640_));
  NA3        g0618(.A(new_new_n640_), .B(new_new_n265_), .C(new_new_n45_), .Y(new_new_n641_));
  OAI220     g0619(.A0(new_new_n641_), .A1(new_new_n639_), .B0(new_new_n638_), .B1(new_new_n1024_), .Y(new_new_n642_));
  NA3        g0620(.A(new_new_n625_), .B(new_new_n317_), .C(i_6_), .Y(new_new_n643_));
  NO2        g0621(.A(new_new_n643_), .B(new_new_n23_), .Y(new_new_n644_));
  AOI210     g0622(.A0(new_new_n476_), .A1(new_new_n421_), .B0(new_new_n243_), .Y(new_new_n645_));
  NO2        g0623(.A(new_new_n645_), .B(new_new_n594_), .Y(new_new_n646_));
  NAi21      g0624(.An(new_new_n637_), .B(new_new_n91_), .Y(new_new_n647_));
  NA2        g0625(.A(new_new_n640_), .B(new_new_n265_), .Y(new_new_n648_));
  NO2        g0626(.A(i_11_), .B(new_new_n37_), .Y(new_new_n649_));
  NA2        g0627(.A(new_new_n649_), .B(new_new_n24_), .Y(new_new_n650_));
  OAI210     g0628(.A0(new_new_n650_), .A1(new_new_n648_), .B0(new_new_n647_), .Y(new_new_n651_));
  OR4        g0629(.A(new_new_n651_), .B(new_new_n646_), .C(new_new_n644_), .D(new_new_n642_), .Y(new_new_n652_));
  NO3        g0630(.A(new_new_n652_), .B(new_new_n636_), .C(new_new_n633_), .Y(new_new_n653_));
  NO2        g0631(.A(new_new_n238_), .B(new_new_n101_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n654_), .B(new_new_n611_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n655_), .B(i_1_), .Y(new_new_n656_));
  NO2        g0634(.A(new_new_n656_), .B(new_new_n605_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n657_), .B(new_new_n47_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n234_), .B(new_new_n45_), .Y(new_new_n659_));
  NO3        g0637(.A(new_new_n659_), .B(new_new_n308_), .C(new_new_n239_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n118_), .B(new_new_n37_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n661_), .B(i_6_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n85_), .B(i_9_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n663_), .B(new_new_n63_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n664_), .B(new_new_n628_), .Y(new_new_n665_));
  NO4        g0643(.A(new_new_n665_), .B(new_new_n662_), .C(new_new_n660_), .D(i_4_), .Y(new_new_n666_));
  NA2        g0644(.A(i_1_), .B(i_3_), .Y(new_new_n667_));
  INV        g0645(.A(new_new_n666_), .Y(new_new_n668_));
  NA4        g0646(.A(new_new_n668_), .B(new_new_n658_), .C(new_new_n653_), .D(new_new_n631_), .Y(new_new_n669_));
  NO3        g0647(.A(new_new_n477_), .B(i_3_), .C(i_7_), .Y(new_new_n670_));
  NOi21      g0648(.An(new_new_n670_), .B(i_10_), .Y(new_new_n671_));
  OA210      g0649(.A0(new_new_n671_), .A1(new_new_n247_), .B0(new_new_n85_), .Y(new_new_n672_));
  NA3        g0650(.A(new_new_n484_), .B(new_new_n513_), .C(new_new_n47_), .Y(new_new_n673_));
  NO3        g0651(.A(new_new_n478_), .B(new_new_n597_), .C(new_new_n85_), .Y(new_new_n674_));
  NA2        g0652(.A(new_new_n674_), .B(new_new_n25_), .Y(new_new_n675_));
  NA3        g0653(.A(new_new_n161_), .B(new_new_n84_), .C(new_new_n85_), .Y(new_new_n676_));
  NA3        g0654(.A(new_new_n676_), .B(new_new_n675_), .C(new_new_n673_), .Y(new_new_n677_));
  OAI210     g0655(.A0(new_new_n677_), .A1(new_new_n672_), .B0(i_1_), .Y(new_new_n678_));
  AOI210     g0656(.A0(new_new_n265_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n679_));
  NO2        g0657(.A(new_new_n372_), .B(i_2_), .Y(new_new_n680_));
  NA2        g0658(.A(new_new_n680_), .B(new_new_n679_), .Y(new_new_n681_));
  OAI210     g0659(.A0(new_new_n643_), .A1(new_new_n447_), .B0(new_new_n681_), .Y(new_new_n682_));
  INV        g0660(.A(new_new_n682_), .Y(new_new_n683_));
  AOI210     g0661(.A0(new_new_n683_), .A1(new_new_n678_), .B0(i_13_), .Y(new_new_n684_));
  OR2        g0662(.A(i_11_), .B(i_7_), .Y(new_new_n685_));
  NA3        g0663(.A(new_new_n685_), .B(new_new_n106_), .C(new_new_n138_), .Y(new_new_n686_));
  AOI220     g0664(.A0(new_new_n470_), .A1(new_new_n161_), .B0(new_new_n449_), .B1(new_new_n138_), .Y(new_new_n687_));
  OAI210     g0665(.A0(new_new_n687_), .A1(new_new_n45_), .B0(new_new_n686_), .Y(new_new_n688_));
  AOI210     g0666(.A0(new_new_n639_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n689_));
  INV        g0667(.A(new_new_n689_), .Y(new_new_n690_));
  NA2        g0668(.A(new_new_n247_), .B(new_new_n132_), .Y(new_new_n691_));
  OAI220     g0669(.A0(new_new_n691_), .A1(new_new_n41_), .B0(new_new_n690_), .B1(new_new_n92_), .Y(new_new_n692_));
  AOI210     g0670(.A0(new_new_n688_), .A1(new_new_n332_), .B0(new_new_n692_), .Y(new_new_n693_));
  INV        g0671(.A(new_new_n115_), .Y(new_new_n694_));
  AOI220     g0672(.A0(new_new_n694_), .A1(new_new_n72_), .B0(new_new_n384_), .B1(new_new_n640_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n695_), .B(new_new_n244_), .Y(new_new_n696_));
  AOI210     g0674(.A0(new_new_n447_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n697_));
  NA2        g0675(.A(new_new_n128_), .B(i_13_), .Y(new_new_n698_));
  NO2        g0676(.A(new_new_n639_), .B(new_new_n115_), .Y(new_new_n699_));
  INV        g0677(.A(new_new_n699_), .Y(new_new_n700_));
  OAI220     g0678(.A0(new_new_n700_), .A1(new_new_n71_), .B0(new_new_n698_), .B1(new_new_n679_), .Y(new_new_n701_));
  NO3        g0679(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n101_), .Y(new_new_n702_));
  NA2        g0680(.A(new_new_n26_), .B(new_new_n195_), .Y(new_new_n703_));
  INV        g0681(.A(new_new_n703_), .Y(new_new_n704_));
  NO3        g0682(.A(new_new_n478_), .B(new_new_n238_), .C(new_new_n85_), .Y(new_new_n705_));
  AOI210     g0683(.A0(new_new_n705_), .A1(new_new_n704_), .B0(new_new_n702_), .Y(new_new_n706_));
  NA2        g0684(.A(new_new_n91_), .B(new_new_n102_), .Y(new_new_n707_));
  OAI220     g0685(.A0(new_new_n707_), .A1(new_new_n592_), .B0(new_new_n706_), .B1(new_new_n607_), .Y(new_new_n708_));
  NO3        g0686(.A(new_new_n708_), .B(new_new_n701_), .C(new_new_n696_), .Y(new_new_n709_));
  OR2        g0687(.A(i_11_), .B(i_6_), .Y(new_new_n710_));
  NA3        g0688(.A(new_new_n591_), .B(new_new_n703_), .C(i_7_), .Y(new_new_n711_));
  AOI210     g0689(.A0(new_new_n711_), .A1(new_new_n700_), .B0(new_new_n710_), .Y(new_new_n712_));
  NA3        g0690(.A(new_new_n410_), .B(new_new_n596_), .C(new_new_n97_), .Y(new_new_n713_));
  NA2        g0691(.A(new_new_n632_), .B(i_13_), .Y(new_new_n714_));
  NA2        g0692(.A(new_new_n102_), .B(new_new_n703_), .Y(new_new_n715_));
  NAi21      g0693(.An(i_11_), .B(i_12_), .Y(new_new_n716_));
  NOi41      g0694(.An(new_new_n111_), .B(new_new_n716_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n717_));
  NO3        g0695(.A(new_new_n478_), .B(new_new_n576_), .C(new_new_n597_), .Y(new_new_n718_));
  AOI220     g0696(.A0(new_new_n718_), .A1(new_new_n312_), .B0(new_new_n717_), .B1(new_new_n715_), .Y(new_new_n719_));
  NA3        g0697(.A(new_new_n719_), .B(new_new_n714_), .C(new_new_n713_), .Y(new_new_n720_));
  OAI210     g0698(.A0(new_new_n720_), .A1(new_new_n712_), .B0(new_new_n63_), .Y(new_new_n721_));
  NO2        g0699(.A(i_2_), .B(i_12_), .Y(new_new_n722_));
  NA2        g0700(.A(new_new_n371_), .B(new_new_n722_), .Y(new_new_n723_));
  NO3        g0701(.A(i_9_), .B(i_3_), .C(new_new_n591_), .Y(new_new_n724_));
  NA2        g0702(.A(new_new_n724_), .B(new_new_n371_), .Y(new_new_n725_));
  NO2        g0703(.A(new_new_n129_), .B(i_2_), .Y(new_new_n726_));
  NA2        g0704(.A(new_new_n726_), .B(new_new_n628_), .Y(new_new_n727_));
  NA3        g0705(.A(new_new_n727_), .B(new_new_n725_), .C(new_new_n723_), .Y(new_new_n728_));
  NA3        g0706(.A(new_new_n728_), .B(new_new_n46_), .C(new_new_n226_), .Y(new_new_n729_));
  NA4        g0707(.A(new_new_n729_), .B(new_new_n721_), .C(new_new_n709_), .D(new_new_n693_), .Y(new_new_n730_));
  OR4        g0708(.A(new_new_n730_), .B(new_new_n684_), .C(new_new_n669_), .D(new_new_n610_), .Y(mai5));
  AOI210     g0709(.A0(new_new_n655_), .A1(new_new_n268_), .B0(new_new_n419_), .Y(new_new_n732_));
  AN2        g0710(.A(new_new_n24_), .B(i_10_), .Y(new_new_n733_));
  NA3        g0711(.A(new_new_n733_), .B(new_new_n722_), .C(new_new_n108_), .Y(new_new_n734_));
  NO2        g0712(.A(new_new_n592_), .B(i_11_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n88_), .B(new_new_n735_), .Y(new_new_n736_));
  NA3        g0714(.A(new_new_n736_), .B(new_new_n734_), .C(new_new_n732_), .Y(new_new_n737_));
  NO3        g0715(.A(i_11_), .B(new_new_n238_), .C(i_13_), .Y(new_new_n738_));
  NO2        g0716(.A(new_new_n125_), .B(new_new_n23_), .Y(new_new_n739_));
  NA2        g0717(.A(i_12_), .B(i_8_), .Y(new_new_n740_));
  OAI210     g0718(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n740_), .Y(new_new_n741_));
  INV        g0719(.A(new_new_n446_), .Y(new_new_n742_));
  AOI220     g0720(.A0(new_new_n317_), .A1(new_new_n569_), .B0(new_new_n741_), .B1(new_new_n739_), .Y(new_new_n743_));
  INV        g0721(.A(new_new_n743_), .Y(new_new_n744_));
  NO2        g0722(.A(new_new_n744_), .B(new_new_n737_), .Y(new_new_n745_));
  INV        g0723(.A(new_new_n172_), .Y(new_new_n746_));
  INV        g0724(.A(new_new_n247_), .Y(new_new_n747_));
  OAI210     g0725(.A0(new_new_n680_), .A1(new_new_n448_), .B0(new_new_n111_), .Y(new_new_n748_));
  AOI210     g0726(.A0(new_new_n748_), .A1(new_new_n747_), .B0(new_new_n746_), .Y(new_new_n749_));
  NO2        g0727(.A(new_new_n456_), .B(new_new_n26_), .Y(new_new_n750_));
  NO2        g0728(.A(new_new_n750_), .B(new_new_n421_), .Y(new_new_n751_));
  NA2        g0729(.A(new_new_n751_), .B(i_2_), .Y(new_new_n752_));
  INV        g0730(.A(new_new_n752_), .Y(new_new_n753_));
  AOI210     g0731(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n417_), .Y(new_new_n754_));
  AOI210     g0732(.A0(new_new_n754_), .A1(new_new_n753_), .B0(new_new_n749_), .Y(new_new_n755_));
  NO2        g0733(.A(new_new_n192_), .B(new_new_n126_), .Y(new_new_n756_));
  OAI210     g0734(.A0(new_new_n756_), .A1(new_new_n739_), .B0(i_2_), .Y(new_new_n757_));
  INV        g0735(.A(new_new_n173_), .Y(new_new_n758_));
  NO3        g0736(.A(new_new_n612_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n759_));
  AOI210     g0737(.A0(new_new_n758_), .A1(new_new_n88_), .B0(new_new_n759_), .Y(new_new_n760_));
  AOI210     g0738(.A0(new_new_n760_), .A1(new_new_n757_), .B0(new_new_n195_), .Y(new_new_n761_));
  OA210      g0739(.A0(new_new_n613_), .A1(new_new_n127_), .B0(i_13_), .Y(new_new_n762_));
  NA2        g0740(.A(new_new_n201_), .B(new_new_n204_), .Y(new_new_n763_));
  NA2        g0741(.A(new_new_n151_), .B(new_new_n588_), .Y(new_new_n764_));
  AOI210     g0742(.A0(new_new_n764_), .A1(new_new_n763_), .B0(new_new_n373_), .Y(new_new_n765_));
  AOI210     g0743(.A0(new_new_n209_), .A1(new_new_n148_), .B0(new_new_n513_), .Y(new_new_n766_));
  NA2        g0744(.A(new_new_n766_), .B(new_new_n421_), .Y(new_new_n767_));
  NO2        g0745(.A(new_new_n102_), .B(new_new_n45_), .Y(new_new_n768_));
  INV        g0746(.A(new_new_n301_), .Y(new_new_n769_));
  NA4        g0747(.A(new_new_n769_), .B(new_new_n305_), .C(new_new_n125_), .D(new_new_n43_), .Y(new_new_n770_));
  OAI210     g0748(.A0(new_new_n770_), .A1(new_new_n768_), .B0(new_new_n767_), .Y(new_new_n771_));
  NO4        g0749(.A(new_new_n771_), .B(new_new_n765_), .C(new_new_n762_), .D(new_new_n761_), .Y(new_new_n772_));
  NA2        g0750(.A(new_new_n569_), .B(new_new_n28_), .Y(new_new_n773_));
  NA2        g0751(.A(new_new_n738_), .B(new_new_n275_), .Y(new_new_n774_));
  NA2        g0752(.A(new_new_n774_), .B(new_new_n773_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n62_), .B(i_12_), .Y(new_new_n776_));
  NO2        g0754(.A(new_new_n776_), .B(new_new_n127_), .Y(new_new_n777_));
  NO2        g0755(.A(new_new_n777_), .B(new_new_n588_), .Y(new_new_n778_));
  AOI220     g0756(.A0(new_new_n778_), .A1(new_new_n36_), .B0(new_new_n775_), .B1(new_new_n47_), .Y(new_new_n779_));
  NA4        g0757(.A(new_new_n779_), .B(new_new_n772_), .C(new_new_n755_), .D(new_new_n745_), .Y(mai6));
  NO3        g0758(.A(i_9_), .B(new_new_n307_), .C(i_1_), .Y(new_new_n781_));
  NO2        g0759(.A(new_new_n187_), .B(new_new_n139_), .Y(new_new_n782_));
  OAI210     g0760(.A0(new_new_n782_), .A1(new_new_n781_), .B0(new_new_n726_), .Y(new_new_n783_));
  NA4        g0761(.A(new_new_n388_), .B(new_new_n483_), .C(new_new_n71_), .D(new_new_n101_), .Y(new_new_n784_));
  INV        g0762(.A(new_new_n784_), .Y(new_new_n785_));
  NO2        g0763(.A(i_11_), .B(i_9_), .Y(new_new_n786_));
  NO2        g0764(.A(new_new_n785_), .B(new_new_n328_), .Y(new_new_n787_));
  AO210      g0765(.A0(new_new_n787_), .A1(new_new_n783_), .B0(i_12_), .Y(new_new_n788_));
  NA2        g0766(.A(new_new_n374_), .B(new_new_n335_), .Y(new_new_n789_));
  NA2        g0767(.A(new_new_n576_), .B(new_new_n63_), .Y(new_new_n790_));
  NA2        g0768(.A(new_new_n671_), .B(new_new_n71_), .Y(new_new_n791_));
  BUFFER     g0769(.A(new_new_n618_), .Y(new_new_n792_));
  NA4        g0770(.A(new_new_n792_), .B(new_new_n791_), .C(new_new_n790_), .D(new_new_n789_), .Y(new_new_n793_));
  INV        g0771(.A(new_new_n198_), .Y(new_new_n794_));
  AOI220     g0772(.A0(new_new_n794_), .A1(new_new_n786_), .B0(new_new_n793_), .B1(new_new_n73_), .Y(new_new_n795_));
  INV        g0773(.A(new_new_n327_), .Y(new_new_n796_));
  NA2        g0774(.A(new_new_n75_), .B(new_new_n132_), .Y(new_new_n797_));
  INV        g0775(.A(new_new_n125_), .Y(new_new_n798_));
  NA2        g0776(.A(new_new_n798_), .B(new_new_n47_), .Y(new_new_n799_));
  AOI210     g0777(.A0(new_new_n799_), .A1(new_new_n797_), .B0(new_new_n796_), .Y(new_new_n800_));
  NO2        g0778(.A(new_new_n32_), .B(i_11_), .Y(new_new_n801_));
  NA3        g0779(.A(new_new_n801_), .B(new_new_n474_), .C(new_new_n388_), .Y(new_new_n802_));
  NAi32      g0780(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n803_));
  AOI210     g0781(.A0(new_new_n710_), .A1(new_new_n86_), .B0(new_new_n803_), .Y(new_new_n804_));
  OAI210     g0782(.A0(new_new_n670_), .A1(new_new_n557_), .B0(new_new_n556_), .Y(new_new_n805_));
  NAi31      g0783(.An(new_new_n804_), .B(new_new_n805_), .C(new_new_n802_), .Y(new_new_n806_));
  OR2        g0784(.A(new_new_n806_), .B(new_new_n800_), .Y(new_new_n807_));
  NO2        g0785(.A(new_new_n685_), .B(i_2_), .Y(new_new_n808_));
  NA2        g0786(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n809_));
  OAI210     g0787(.A0(new_new_n809_), .A1(new_new_n409_), .B0(new_new_n361_), .Y(new_new_n810_));
  NA2        g0788(.A(new_new_n810_), .B(new_new_n808_), .Y(new_new_n811_));
  AO210      g0789(.A0(new_new_n360_), .A1(new_new_n351_), .B0(new_new_n395_), .Y(new_new_n812_));
  NA3        g0790(.A(new_new_n812_), .B(new_new_n256_), .C(i_7_), .Y(new_new_n813_));
  OR2        g0791(.A(new_new_n613_), .B(new_new_n448_), .Y(new_new_n814_));
  NA3        g0792(.A(new_new_n814_), .B(new_new_n147_), .C(new_new_n69_), .Y(new_new_n815_));
  OR2        g0793(.A(new_new_n742_), .B(new_new_n36_), .Y(new_new_n816_));
  NA4        g0794(.A(new_new_n816_), .B(new_new_n815_), .C(new_new_n813_), .D(new_new_n811_), .Y(new_new_n817_));
  OAI210     g0795(.A0(i_6_), .A1(i_11_), .B0(new_new_n86_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n818_), .B(new_new_n556_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n395_), .B(new_new_n70_), .Y(new_new_n820_));
  NA3        g0798(.A(new_new_n820_), .B(new_new_n819_), .C(new_new_n595_), .Y(new_new_n821_));
  AO210      g0799(.A0(new_new_n513_), .A1(new_new_n47_), .B0(new_new_n87_), .Y(new_new_n822_));
  NA3        g0800(.A(new_new_n822_), .B(new_new_n484_), .C(new_new_n219_), .Y(new_new_n823_));
  AOI210     g0801(.A0(new_new_n448_), .A1(new_new_n446_), .B0(new_new_n555_), .Y(new_new_n824_));
  NA2        g0802(.A(new_new_n112_), .B(new_new_n408_), .Y(new_new_n825_));
  NA2        g0803(.A(new_new_n246_), .B(new_new_n47_), .Y(new_new_n826_));
  NA3        g0804(.A(new_new_n825_), .B(new_new_n824_), .C(new_new_n823_), .Y(new_new_n827_));
  NO4        g0805(.A(new_new_n827_), .B(new_new_n821_), .C(new_new_n817_), .D(new_new_n807_), .Y(new_new_n828_));
  NA4        g0806(.A(new_new_n828_), .B(new_new_n795_), .C(new_new_n788_), .D(new_new_n379_), .Y(mai3));
  NA2        g0807(.A(i_6_), .B(i_7_), .Y(new_new_n830_));
  NO2        g0808(.A(new_new_n830_), .B(i_0_), .Y(new_new_n831_));
  NO2        g0809(.A(i_11_), .B(new_new_n238_), .Y(new_new_n832_));
  OAI210     g0810(.A0(new_new_n831_), .A1(new_new_n289_), .B0(new_new_n832_), .Y(new_new_n833_));
  NO2        g0811(.A(new_new_n833_), .B(new_new_n195_), .Y(new_new_n834_));
  NO3        g0812(.A(new_new_n452_), .B(new_new_n89_), .C(new_new_n45_), .Y(new_new_n835_));
  OA210      g0813(.A0(new_new_n835_), .A1(new_new_n834_), .B0(new_new_n175_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n410_), .B(new_new_n46_), .Y(new_new_n837_));
  NO4        g0815(.A(new_new_n375_), .B(new_new_n382_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n838_));
  INV        g0816(.A(new_new_n838_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n697_), .B(new_new_n663_), .Y(new_new_n840_));
  NA2        g0818(.A(new_new_n333_), .B(new_new_n438_), .Y(new_new_n841_));
  OAI220     g0819(.A0(new_new_n841_), .A1(new_new_n840_), .B0(new_new_n839_), .B1(new_new_n63_), .Y(new_new_n842_));
  NOi21      g0820(.An(i_5_), .B(i_9_), .Y(new_new_n843_));
  NA2        g0821(.A(new_new_n843_), .B(new_new_n445_), .Y(new_new_n844_));
  AOI210     g0822(.A0(new_new_n265_), .A1(new_new_n476_), .B0(new_new_n674_), .Y(new_new_n845_));
  NO3        g0823(.A(new_new_n413_), .B(new_new_n265_), .C(new_new_n73_), .Y(new_new_n846_));
  NO2        g0824(.A(new_new_n176_), .B(new_new_n148_), .Y(new_new_n847_));
  AOI210     g0825(.A0(new_new_n847_), .A1(new_new_n246_), .B0(new_new_n846_), .Y(new_new_n848_));
  OAI220     g0826(.A0(new_new_n848_), .A1(new_new_n182_), .B0(new_new_n845_), .B1(new_new_n844_), .Y(new_new_n849_));
  NO3        g0827(.A(new_new_n849_), .B(new_new_n842_), .C(new_new_n836_), .Y(new_new_n850_));
  NA2        g0828(.A(new_new_n187_), .B(new_new_n24_), .Y(new_new_n851_));
  NO2        g0829(.A(new_new_n661_), .B(new_new_n586_), .Y(new_new_n852_));
  NO2        g0830(.A(new_new_n852_), .B(new_new_n851_), .Y(new_new_n853_));
  NA2        g0831(.A(new_new_n312_), .B(new_new_n130_), .Y(new_new_n854_));
  NAi21      g0832(.An(new_new_n162_), .B(new_new_n438_), .Y(new_new_n855_));
  OAI220     g0833(.A0(new_new_n855_), .A1(new_new_n826_), .B0(new_new_n854_), .B1(new_new_n400_), .Y(new_new_n856_));
  NO2        g0834(.A(new_new_n856_), .B(new_new_n853_), .Y(new_new_n857_));
  NO2        g0835(.A(new_new_n388_), .B(new_new_n293_), .Y(new_new_n858_));
  NA2        g0836(.A(new_new_n858_), .B(new_new_n699_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n566_), .B(i_0_), .Y(new_new_n860_));
  NO3        g0838(.A(new_new_n860_), .B(new_new_n383_), .C(new_new_n88_), .Y(new_new_n861_));
  INV        g0839(.A(new_new_n861_), .Y(new_new_n862_));
  AN2        g0840(.A(new_new_n96_), .B(new_new_n245_), .Y(new_new_n863_));
  NA2        g0841(.A(new_new_n738_), .B(new_new_n328_), .Y(new_new_n864_));
  INV        g0842(.A(new_new_n58_), .Y(new_new_n865_));
  OAI220     g0843(.A0(new_new_n865_), .A1(new_new_n864_), .B0(new_new_n650_), .B1(new_new_n531_), .Y(new_new_n866_));
  NA2        g0844(.A(i_0_), .B(i_10_), .Y(new_new_n867_));
  NA2        g0845(.A(new_new_n187_), .B(new_new_n84_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n560_), .B(i_4_), .Y(new_new_n869_));
  NA2        g0847(.A(new_new_n190_), .B(new_new_n204_), .Y(new_new_n870_));
  OAI220     g0848(.A0(new_new_n870_), .A1(new_new_n864_), .B0(new_new_n869_), .B1(new_new_n868_), .Y(new_new_n871_));
  NO3        g0849(.A(new_new_n871_), .B(new_new_n866_), .C(new_new_n863_), .Y(new_new_n872_));
  NA4        g0850(.A(new_new_n872_), .B(new_new_n862_), .C(new_new_n859_), .D(new_new_n857_), .Y(new_new_n873_));
  NA2        g0851(.A(i_11_), .B(i_9_), .Y(new_new_n874_));
  NO2        g0852(.A(new_new_n49_), .B(i_7_), .Y(new_new_n875_));
  NA2        g0853(.A(new_new_n393_), .B(new_new_n180_), .Y(new_new_n876_));
  NA2        g0854(.A(new_new_n876_), .B(new_new_n160_), .Y(new_new_n877_));
  NO2        g0855(.A(new_new_n874_), .B(new_new_n73_), .Y(new_new_n878_));
  NO2        g0856(.A(new_new_n176_), .B(i_0_), .Y(new_new_n879_));
  INV        g0857(.A(new_new_n879_), .Y(new_new_n880_));
  NA2        g0858(.A(new_new_n474_), .B(new_new_n232_), .Y(new_new_n881_));
  NO2        g0859(.A(new_new_n881_), .B(new_new_n880_), .Y(new_new_n882_));
  NO2        g0860(.A(new_new_n882_), .B(new_new_n877_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n649_), .B(new_new_n122_), .Y(new_new_n884_));
  NO2        g0862(.A(i_6_), .B(new_new_n884_), .Y(new_new_n885_));
  AOI210     g0863(.A0(new_new_n447_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n172_), .B(new_new_n103_), .Y(new_new_n887_));
  NOi32      g0865(.An(new_new_n886_), .Bn(new_new_n190_), .C(new_new_n887_), .Y(new_new_n888_));
  NA2        g0866(.A(new_new_n596_), .B(new_new_n328_), .Y(new_new_n889_));
  NO2        g0867(.A(new_new_n889_), .B(new_new_n837_), .Y(new_new_n890_));
  NO3        g0868(.A(new_new_n890_), .B(new_new_n888_), .C(new_new_n885_), .Y(new_new_n891_));
  NOi21      g0869(.An(i_7_), .B(i_5_), .Y(new_new_n892_));
  NOi31      g0870(.An(new_new_n892_), .B(i_0_), .C(new_new_n716_), .Y(new_new_n893_));
  NA3        g0871(.A(new_new_n893_), .B(i_3_), .C(i_6_), .Y(new_new_n894_));
  BUFFER     g0872(.A(new_new_n894_), .Y(new_new_n895_));
  NO3        g0873(.A(new_new_n403_), .B(new_new_n363_), .C(new_new_n359_), .Y(new_new_n896_));
  NO2        g0874(.A(new_new_n259_), .B(new_new_n318_), .Y(new_new_n897_));
  INV        g0875(.A(new_new_n716_), .Y(new_new_n898_));
  AOI210     g0876(.A0(new_new_n898_), .A1(new_new_n897_), .B0(new_new_n896_), .Y(new_new_n899_));
  NA4        g0877(.A(new_new_n899_), .B(new_new_n895_), .C(new_new_n891_), .D(new_new_n883_), .Y(new_new_n900_));
  NO2        g0878(.A(new_new_n851_), .B(new_new_n241_), .Y(new_new_n901_));
  AN2        g0879(.A(new_new_n332_), .B(new_new_n328_), .Y(new_new_n902_));
  AN2        g0880(.A(new_new_n902_), .B(new_new_n847_), .Y(new_new_n903_));
  OAI210     g0881(.A0(new_new_n903_), .A1(new_new_n901_), .B0(i_10_), .Y(new_new_n904_));
  OA210      g0882(.A0(new_new_n474_), .A1(new_new_n224_), .B0(new_new_n473_), .Y(new_new_n905_));
  NA3        g0883(.A(new_new_n473_), .B(new_new_n410_), .C(new_new_n46_), .Y(new_new_n906_));
  OAI210     g0884(.A0(new_new_n855_), .A1(i_6_), .B0(new_new_n906_), .Y(new_new_n907_));
  NA2        g0885(.A(new_new_n878_), .B(new_new_n305_), .Y(new_new_n908_));
  NA2        g0886(.A(new_new_n189_), .B(new_new_n908_), .Y(new_new_n909_));
  AOI220     g0887(.A0(new_new_n909_), .A1(new_new_n474_), .B0(new_new_n907_), .B1(new_new_n73_), .Y(new_new_n910_));
  NO2        g0888(.A(new_new_n75_), .B(new_new_n740_), .Y(new_new_n911_));
  AOI220     g0889(.A0(new_new_n911_), .A1(i_11_), .B0(new_new_n175_), .B1(new_new_n586_), .Y(new_new_n912_));
  NO2        g0890(.A(new_new_n912_), .B(new_new_n48_), .Y(new_new_n913_));
  NO3        g0891(.A(i_5_), .B(new_new_n358_), .C(new_new_n24_), .Y(new_new_n914_));
  INV        g0892(.A(new_new_n914_), .Y(new_new_n915_));
  NAi21      g0893(.An(i_9_), .B(i_5_), .Y(new_new_n916_));
  NO2        g0894(.A(new_new_n590_), .B(new_new_n105_), .Y(new_new_n917_));
  NA2        g0895(.A(new_new_n917_), .B(i_0_), .Y(new_new_n918_));
  OAI220     g0896(.A0(new_new_n918_), .A1(new_new_n85_), .B0(new_new_n915_), .B1(new_new_n173_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n919_), .B(new_new_n913_), .Y(new_new_n920_));
  NA3        g0898(.A(new_new_n920_), .B(new_new_n910_), .C(new_new_n904_), .Y(new_new_n921_));
  NO3        g0899(.A(new_new_n921_), .B(new_new_n900_), .C(new_new_n873_), .Y(new_new_n922_));
  NO2        g0900(.A(i_0_), .B(new_new_n716_), .Y(new_new_n923_));
  NA2        g0901(.A(new_new_n73_), .B(new_new_n45_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n790_), .B(new_new_n887_), .Y(new_new_n925_));
  INV        g0903(.A(new_new_n925_), .Y(new_new_n926_));
  NA2        g0904(.A(new_new_n726_), .B(new_new_n146_), .Y(new_new_n927_));
  INV        g0905(.A(new_new_n927_), .Y(new_new_n928_));
  NA3        g0906(.A(new_new_n928_), .B(new_new_n663_), .C(new_new_n73_), .Y(new_new_n929_));
  NO2        g0907(.A(new_new_n805_), .B(new_new_n403_), .Y(new_new_n930_));
  NA2        g0908(.A(new_new_n246_), .B(new_new_n231_), .Y(new_new_n931_));
  AOI210     g0909(.A0(new_new_n931_), .A1(new_new_n860_), .B0(new_new_n153_), .Y(new_new_n932_));
  NO2        g0910(.A(new_new_n932_), .B(new_new_n930_), .Y(new_new_n933_));
  NA3        g0911(.A(new_new_n933_), .B(new_new_n929_), .C(new_new_n926_), .Y(new_new_n934_));
  NA2        g0912(.A(new_new_n902_), .B(new_new_n373_), .Y(new_new_n935_));
  AOI210     g0913(.A0(new_new_n300_), .A1(new_new_n162_), .B0(new_new_n935_), .Y(new_new_n936_));
  NA3        g0914(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n875_), .B(new_new_n488_), .Y(new_new_n938_));
  AOI210     g0916(.A0(new_new_n937_), .A1(new_new_n162_), .B0(new_new_n938_), .Y(new_new_n939_));
  NO2        g0917(.A(new_new_n939_), .B(new_new_n936_), .Y(new_new_n940_));
  NO3        g0918(.A(new_new_n867_), .B(new_new_n843_), .C(new_new_n192_), .Y(new_new_n941_));
  AOI220     g0919(.A0(new_new_n941_), .A1(i_11_), .B0(new_new_n561_), .B1(new_new_n75_), .Y(new_new_n942_));
  NO3        g0920(.A(new_new_n210_), .B(new_new_n382_), .C(i_0_), .Y(new_new_n943_));
  OAI210     g0921(.A0(new_new_n943_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n944_));
  INV        g0922(.A(new_new_n219_), .Y(new_new_n945_));
  NO2        g0923(.A(new_new_n524_), .B(new_new_n139_), .Y(new_new_n946_));
  NA3        g0924(.A(new_new_n946_), .B(i_7_), .C(new_new_n945_), .Y(new_new_n947_));
  NA4        g0925(.A(new_new_n947_), .B(new_new_n944_), .C(new_new_n942_), .D(new_new_n940_), .Y(new_new_n948_));
  INV        g0926(.A(new_new_n92_), .Y(new_new_n949_));
  AOI210     g0927(.A0(new_new_n949_), .A1(new_new_n923_), .B0(new_new_n109_), .Y(new_new_n950_));
  AOI220     g0928(.A0(new_new_n892_), .A1(new_new_n488_), .B0(new_new_n831_), .B1(new_new_n163_), .Y(new_new_n951_));
  NA2        g0929(.A(new_new_n351_), .B(new_new_n177_), .Y(new_new_n952_));
  OA220      g0930(.A0(new_new_n952_), .A1(new_new_n951_), .B0(new_new_n950_), .B1(i_5_), .Y(new_new_n953_));
  AOI210     g0931(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n176_), .Y(new_new_n954_));
  NA2        g0932(.A(new_new_n954_), .B(new_new_n905_), .Y(new_new_n955_));
  NO3        g0933(.A(new_new_n837_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n956_));
  NA2        g0934(.A(new_new_n493_), .B(new_new_n471_), .Y(new_new_n957_));
  NO2        g0935(.A(new_new_n957_), .B(new_new_n956_), .Y(new_new_n958_));
  NA3        g0936(.A(new_new_n388_), .B(new_new_n172_), .C(new_new_n171_), .Y(new_new_n959_));
  NA3        g0937(.A(new_new_n875_), .B(new_new_n289_), .C(new_new_n231_), .Y(new_new_n960_));
  NA2        g0938(.A(new_new_n960_), .B(new_new_n959_), .Y(new_new_n961_));
  NA3        g0939(.A(new_new_n388_), .B(new_new_n334_), .C(new_new_n222_), .Y(new_new_n962_));
  INV        g0940(.A(new_new_n962_), .Y(new_new_n963_));
  NOi31      g0941(.An(new_new_n387_), .B(new_new_n924_), .C(new_new_n241_), .Y(new_new_n964_));
  NO3        g0942(.A(new_new_n874_), .B(new_new_n219_), .C(new_new_n192_), .Y(new_new_n965_));
  NO4        g0943(.A(new_new_n965_), .B(new_new_n964_), .C(new_new_n963_), .D(new_new_n961_), .Y(new_new_n966_));
  NA4        g0944(.A(new_new_n966_), .B(new_new_n958_), .C(new_new_n955_), .D(new_new_n953_), .Y(new_new_n967_));
  NA2        g0945(.A(new_new_n305_), .B(i_5_), .Y(new_new_n968_));
  NA2        g0946(.A(new_new_n968_), .B(new_new_n244_), .Y(new_new_n969_));
  NO4        g0947(.A(new_new_n241_), .B(new_new_n210_), .C(i_0_), .D(i_12_), .Y(new_new_n970_));
  AOI220     g0948(.A0(new_new_n970_), .A1(new_new_n969_), .B0(new_new_n785_), .B1(new_new_n177_), .Y(new_new_n971_));
  AN2        g0949(.A(new_new_n867_), .B(new_new_n153_), .Y(new_new_n972_));
  NO4        g0950(.A(new_new_n972_), .B(i_12_), .C(new_new_n637_), .D(new_new_n132_), .Y(new_new_n973_));
  NA2        g0951(.A(new_new_n973_), .B(new_new_n219_), .Y(new_new_n974_));
  NA3        g0952(.A(new_new_n98_), .B(new_new_n565_), .C(i_11_), .Y(new_new_n975_));
  NO2        g0953(.A(new_new_n975_), .B(new_new_n155_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n892_), .B(new_new_n470_), .Y(new_new_n977_));
  NA2        g0955(.A(new_new_n64_), .B(new_new_n101_), .Y(new_new_n978_));
  OAI220     g0956(.A0(new_new_n978_), .A1(new_new_n968_), .B0(new_new_n977_), .B1(new_new_n664_), .Y(new_new_n979_));
  AOI210     g0957(.A0(new_new_n979_), .A1(new_new_n879_), .B0(new_new_n976_), .Y(new_new_n980_));
  NA3        g0958(.A(new_new_n980_), .B(new_new_n974_), .C(new_new_n971_), .Y(new_new_n981_));
  NO4        g0959(.A(new_new_n981_), .B(new_new_n967_), .C(new_new_n948_), .D(new_new_n934_), .Y(new_new_n982_));
  OAI210     g0960(.A0(new_new_n808_), .A1(new_new_n801_), .B0(new_new_n37_), .Y(new_new_n983_));
  NA3        g0961(.A(new_new_n886_), .B(new_new_n371_), .C(i_5_), .Y(new_new_n984_));
  NA3        g0962(.A(new_new_n984_), .B(new_new_n983_), .C(new_new_n602_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n985_), .B(new_new_n207_), .Y(new_new_n986_));
  NA2        g0964(.A(new_new_n188_), .B(new_new_n190_), .Y(new_new_n987_));
  AO210      g0965(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n987_), .Y(new_new_n988_));
  OAI210     g0966(.A0(new_new_n606_), .A1(new_new_n604_), .B0(new_new_n317_), .Y(new_new_n989_));
  NA2        g0967(.A(new_new_n989_), .B(new_new_n988_), .Y(new_new_n990_));
  NO2        g0968(.A(new_new_n461_), .B(new_new_n265_), .Y(new_new_n991_));
  NO4        g0969(.A(new_new_n234_), .B(new_new_n145_), .C(new_new_n667_), .D(new_new_n37_), .Y(new_new_n992_));
  NO2        g0970(.A(new_new_n992_), .B(new_new_n991_), .Y(new_new_n993_));
  OAI210     g0971(.A0(new_new_n975_), .A1(new_new_n148_), .B0(new_new_n993_), .Y(new_new_n994_));
  AOI210     g0972(.A0(new_new_n990_), .A1(new_new_n49_), .B0(new_new_n994_), .Y(new_new_n995_));
  AOI210     g0973(.A0(new_new_n995_), .A1(new_new_n986_), .B0(new_new_n73_), .Y(new_new_n996_));
  NO2        g0974(.A(new_new_n558_), .B(new_new_n378_), .Y(new_new_n997_));
  NO2        g0975(.A(new_new_n997_), .B(new_new_n746_), .Y(new_new_n998_));
  INV        g0976(.A(new_new_n76_), .Y(new_new_n999_));
  AOI210     g0977(.A0(new_new_n954_), .A1(new_new_n875_), .B0(new_new_n893_), .Y(new_new_n1000_));
  AOI210     g0978(.A0(new_new_n1000_), .A1(new_new_n999_), .B0(new_new_n667_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n259_), .B(new_new_n57_), .Y(new_new_n1002_));
  NA2        g0980(.A(new_new_n1002_), .B(new_new_n76_), .Y(new_new_n1003_));
  NO2        g0981(.A(new_new_n1003_), .B(new_new_n238_), .Y(new_new_n1004_));
  NA3        g0982(.A(new_new_n96_), .B(new_new_n307_), .C(new_new_n31_), .Y(new_new_n1005_));
  INV        g0983(.A(new_new_n1005_), .Y(new_new_n1006_));
  NO3        g0984(.A(new_new_n1006_), .B(new_new_n1004_), .C(new_new_n1001_), .Y(new_new_n1007_));
  OAI210     g0985(.A0(new_new_n267_), .A1(new_new_n158_), .B0(new_new_n88_), .Y(new_new_n1008_));
  NA3        g0986(.A(new_new_n750_), .B(new_new_n289_), .C(new_new_n80_), .Y(new_new_n1009_));
  AOI210     g0987(.A0(new_new_n1009_), .A1(new_new_n1008_), .B0(i_11_), .Y(new_new_n1010_));
  OAI210     g0988(.A0(new_new_n1025_), .A1(new_new_n886_), .B0(new_new_n207_), .Y(new_new_n1011_));
  NA2        g0989(.A(new_new_n164_), .B(i_5_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n1011_), .A1(new_new_n763_), .B0(new_new_n1012_), .Y(new_new_n1013_));
  NO4        g0991(.A(new_new_n916_), .B(new_new_n477_), .C(new_new_n255_), .D(new_new_n254_), .Y(new_new_n1014_));
  NO2        g0992(.A(new_new_n1014_), .B(new_new_n555_), .Y(new_new_n1015_));
  INV        g0993(.A(new_new_n364_), .Y(new_new_n1016_));
  AOI210     g0994(.A0(new_new_n1016_), .A1(new_new_n1015_), .B0(new_new_n41_), .Y(new_new_n1017_));
  NO3        g0995(.A(new_new_n1017_), .B(new_new_n1013_), .C(new_new_n1010_), .Y(new_new_n1018_));
  OAI210     g0996(.A0(new_new_n1007_), .A1(i_4_), .B0(new_new_n1018_), .Y(new_new_n1019_));
  NO3        g0997(.A(new_new_n1019_), .B(new_new_n998_), .C(new_new_n996_), .Y(new_new_n1020_));
  NA4        g0998(.A(new_new_n1020_), .B(new_new_n982_), .C(new_new_n922_), .D(new_new_n850_), .Y(mai4));
  INV        g0999(.A(i_2_), .Y(new_new_n1024_));
  INV        g1000(.A(i_12_), .Y(new_new_n1025_));
  INV        g1001(.A(i_12_), .Y(new_new_n1026_));
  INV        g1002(.A(new_new_n82_), .Y(new_new_n1027_));
endmodule


