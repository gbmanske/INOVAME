// Benchmark "top" written by ABC on Thu Jun 20 14:59:19 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n134_, new_new_n135_,
    new_new_n136_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n678_,
    new_new_n679_, new_new_n680_, new_new_n681_, new_new_n682_,
    new_new_n683_, new_new_n684_, new_new_n685_, new_new_n686_,
    new_new_n687_, new_new_n688_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n720_, new_new_n721_, new_new_n722_, new_new_n723_,
    new_new_n724_, new_new_n725_, new_new_n726_, new_new_n727_,
    new_new_n728_, new_new_n729_, new_new_n730_, new_new_n731_,
    new_new_n732_, new_new_n733_, new_new_n734_, new_new_n735_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n963_,
    new_new_n964_, new_new_n965_, new_new_n966_, new_new_n967_,
    new_new_n968_, new_new_n969_, new_new_n970_, new_new_n971_,
    new_new_n972_, new_new_n973_, new_new_n974_, new_new_n975_,
    new_new_n976_, new_new_n977_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g021(.A(new_new_n35_), .Y(men1));
  INV        g022(.A(i_11_), .Y(new_new_n45_));
  NO2        g023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g024(.A(i_2_), .Y(new_new_n47_));
  NA2        g025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g026(.A(i_5_), .Y(new_new_n49_));
  NO2        g027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NO2        g035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  NAi21      g037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g038(.A(i_1_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n51_), .B(i_2_), .Y(new_new_n63_));
  AOI210     g041(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n64_));
  NA2        g042(.A(i_1_), .B(i_6_), .Y(new_new_n65_));
  NO2        g043(.A(new_new_n65_), .B(new_new_n25_), .Y(new_new_n66_));
  INV        g044(.A(i_0_), .Y(new_new_n67_));
  NAi21      g045(.An(i_5_), .B(i_10_), .Y(new_new_n68_));
  NA2        g046(.A(i_5_), .B(i_9_), .Y(new_new_n69_));
  AOI210     g047(.A0(new_new_n69_), .A1(new_new_n68_), .B0(new_new_n67_), .Y(new_new_n70_));
  NO2        g048(.A(new_new_n70_), .B(new_new_n66_), .Y(new_new_n71_));
  OAI210     g049(.A0(new_new_n64_), .A1(new_new_n63_), .B0(new_new_n71_), .Y(new_new_n72_));
  NA2        g050(.A(new_new_n72_), .B(i_0_), .Y(new_new_n73_));
  NA2        g051(.A(i_12_), .B(i_5_), .Y(new_new_n74_));
  NA2        g052(.A(i_2_), .B(i_8_), .Y(new_new_n75_));
  NO2        g053(.A(i_3_), .B(i_9_), .Y(new_new_n76_));
  NO2        g054(.A(i_3_), .B(i_7_), .Y(new_new_n77_));
  NO3        g055(.A(new_new_n77_), .B(new_new_n76_), .C(new_new_n61_), .Y(new_new_n78_));
  INV        g056(.A(i_6_), .Y(new_new_n79_));
  OR4        g057(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n80_));
  INV        g058(.A(new_new_n80_), .Y(new_new_n81_));
  NO2        g059(.A(i_2_), .B(i_7_), .Y(new_new_n82_));
  OAI210     g060(.A0(new_new_n78_), .A1(i_8_), .B0(i_2_), .Y(new_new_n83_));
  NAi21      g061(.An(i_6_), .B(i_10_), .Y(new_new_n84_));
  NA2        g062(.A(i_6_), .B(i_9_), .Y(new_new_n85_));
  AOI210     g063(.A0(new_new_n85_), .A1(new_new_n84_), .B0(new_new_n61_), .Y(new_new_n86_));
  NA2        g064(.A(i_2_), .B(i_6_), .Y(new_new_n87_));
  NO3        g065(.A(new_new_n87_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n88_));
  NO2        g066(.A(new_new_n88_), .B(new_new_n86_), .Y(new_new_n89_));
  AOI210     g067(.A0(new_new_n89_), .A1(new_new_n83_), .B0(new_new_n74_), .Y(new_new_n90_));
  AN3        g068(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n91_));
  NAi21      g069(.An(i_6_), .B(i_11_), .Y(new_new_n92_));
  NO2        g070(.A(i_5_), .B(i_8_), .Y(new_new_n93_));
  NOi21      g071(.An(new_new_n93_), .B(new_new_n92_), .Y(new_new_n94_));
  AOI220     g072(.A0(new_new_n94_), .A1(new_new_n60_), .B0(new_new_n91_), .B1(new_new_n32_), .Y(new_new_n95_));
  INV        g073(.A(i_7_), .Y(new_new_n96_));
  NA2        g074(.A(new_new_n47_), .B(new_new_n96_), .Y(new_new_n97_));
  NO2        g075(.A(i_0_), .B(i_5_), .Y(new_new_n98_));
  NO2        g076(.A(new_new_n98_), .B(new_new_n79_), .Y(new_new_n99_));
  NA2        g077(.A(i_12_), .B(i_3_), .Y(new_new_n100_));
  INV        g078(.A(new_new_n100_), .Y(new_new_n101_));
  NA3        g079(.A(new_new_n101_), .B(new_new_n99_), .C(new_new_n97_), .Y(new_new_n102_));
  NAi21      g080(.An(i_7_), .B(i_11_), .Y(new_new_n103_));
  NO3        g081(.A(new_new_n103_), .B(new_new_n84_), .C(new_new_n54_), .Y(new_new_n104_));
  AN2        g082(.A(i_2_), .B(i_10_), .Y(new_new_n105_));
  NO2        g083(.A(new_new_n105_), .B(i_7_), .Y(new_new_n106_));
  OR2        g084(.A(new_new_n74_), .B(new_new_n58_), .Y(new_new_n107_));
  NO2        g085(.A(i_8_), .B(new_new_n96_), .Y(new_new_n108_));
  NO3        g086(.A(new_new_n108_), .B(new_new_n107_), .C(new_new_n106_), .Y(new_new_n109_));
  NA2        g087(.A(i_12_), .B(i_7_), .Y(new_new_n110_));
  NO2        g088(.A(new_new_n61_), .B(new_new_n26_), .Y(new_new_n111_));
  NA2        g089(.A(new_new_n111_), .B(i_0_), .Y(new_new_n112_));
  NA2        g090(.A(i_11_), .B(i_12_), .Y(new_new_n113_));
  OAI210     g091(.A0(new_new_n112_), .A1(new_new_n110_), .B0(new_new_n113_), .Y(new_new_n114_));
  NO2        g092(.A(new_new_n114_), .B(new_new_n109_), .Y(new_new_n115_));
  NAi41      g093(.An(new_new_n104_), .B(new_new_n115_), .C(new_new_n102_), .D(new_new_n95_), .Y(new_new_n116_));
  NOi21      g094(.An(i_1_), .B(i_5_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(i_11_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n96_), .B(new_new_n37_), .Y(new_new_n119_));
  NA2        g097(.A(i_7_), .B(new_new_n25_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(new_new_n119_), .Y(new_new_n121_));
  NO2        g099(.A(new_new_n121_), .B(new_new_n47_), .Y(new_new_n122_));
  NA2        g100(.A(new_new_n85_), .B(new_new_n84_), .Y(new_new_n123_));
  NAi21      g101(.An(i_3_), .B(i_8_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(new_new_n60_), .Y(new_new_n125_));
  NOi31      g103(.An(new_new_n125_), .B(new_new_n123_), .C(new_new_n122_), .Y(new_new_n126_));
  NO2        g104(.A(i_1_), .B(new_new_n79_), .Y(new_new_n127_));
  NO2        g105(.A(i_6_), .B(i_5_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(i_3_), .Y(new_new_n129_));
  AO210      g107(.A0(new_new_n129_), .A1(new_new_n48_), .B0(new_new_n127_), .Y(new_new_n130_));
  OAI220     g108(.A0(new_new_n130_), .A1(new_new_n103_), .B0(new_new_n126_), .B1(new_new_n118_), .Y(new_new_n131_));
  NO3        g109(.A(new_new_n131_), .B(new_new_n116_), .C(new_new_n90_), .Y(new_new_n132_));
  NA3        g110(.A(new_new_n132_), .B(new_new_n73_), .C(new_new_n57_), .Y(men2));
  NO2        g111(.A(new_new_n61_), .B(new_new_n37_), .Y(new_new_n134_));
  NA2        g112(.A(i_6_), .B(new_new_n25_), .Y(new_new_n135_));
  NA2        g113(.A(new_new_n135_), .B(new_new_n134_), .Y(new_new_n136_));
  NA4        g114(.A(new_new_n136_), .B(new_new_n71_), .C(new_new_n63_), .D(new_new_n30_), .Y(men0));
  AN2        g115(.A(i_8_), .B(i_7_), .Y(new_new_n138_));
  NA2        g116(.A(new_new_n138_), .B(i_6_), .Y(new_new_n139_));
  NO2        g117(.A(i_12_), .B(i_13_), .Y(new_new_n140_));
  NAi21      g118(.An(i_5_), .B(i_11_), .Y(new_new_n141_));
  NOi21      g119(.An(new_new_n140_), .B(new_new_n141_), .Y(new_new_n142_));
  NO2        g120(.A(i_0_), .B(i_1_), .Y(new_new_n143_));
  NA2        g121(.A(i_2_), .B(i_3_), .Y(new_new_n144_));
  NO2        g122(.A(new_new_n144_), .B(i_4_), .Y(new_new_n145_));
  NA3        g123(.A(new_new_n145_), .B(new_new_n143_), .C(new_new_n142_), .Y(new_new_n146_));
  OR2        g124(.A(new_new_n146_), .B(new_new_n25_), .Y(new_new_n147_));
  AN2        g125(.A(new_new_n140_), .B(new_new_n76_), .Y(new_new_n148_));
  NO2        g126(.A(new_new_n148_), .B(new_new_n27_), .Y(new_new_n149_));
  NA2        g127(.A(i_1_), .B(i_5_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n67_), .B(new_new_n47_), .Y(new_new_n151_));
  NA2        g129(.A(new_new_n151_), .B(new_new_n36_), .Y(new_new_n152_));
  NO3        g130(.A(new_new_n152_), .B(new_new_n150_), .C(new_new_n149_), .Y(new_new_n153_));
  OR2        g131(.A(i_0_), .B(i_1_), .Y(new_new_n154_));
  NO3        g132(.A(new_new_n154_), .B(new_new_n74_), .C(i_13_), .Y(new_new_n155_));
  NAi32      g133(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n156_));
  NAi21      g134(.An(new_new_n156_), .B(new_new_n155_), .Y(new_new_n157_));
  NOi21      g135(.An(i_4_), .B(i_10_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n40_), .Y(new_new_n159_));
  NO2        g137(.A(i_3_), .B(i_5_), .Y(new_new_n160_));
  NO3        g138(.A(new_new_n67_), .B(i_2_), .C(i_1_), .Y(new_new_n161_));
  OAI210     g139(.A0(i_3_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n162_));
  NO2        g140(.A(new_new_n162_), .B(new_new_n153_), .Y(new_new_n163_));
  AOI210     g141(.A0(new_new_n163_), .A1(new_new_n147_), .B0(new_new_n139_), .Y(new_new_n164_));
  NA2        g142(.A(i_3_), .B(new_new_n49_), .Y(new_new_n165_));
  NOi21      g143(.An(i_4_), .B(i_9_), .Y(new_new_n166_));
  NOi21      g144(.An(i_11_), .B(i_13_), .Y(new_new_n167_));
  NA2        g145(.A(new_new_n167_), .B(new_new_n166_), .Y(new_new_n168_));
  OR2        g146(.A(new_new_n168_), .B(new_new_n165_), .Y(new_new_n169_));
  NO2        g147(.A(i_4_), .B(i_5_), .Y(new_new_n170_));
  NAi21      g148(.An(i_12_), .B(i_11_), .Y(new_new_n171_));
  NO2        g149(.A(new_new_n171_), .B(i_13_), .Y(new_new_n172_));
  NA3        g150(.A(new_new_n172_), .B(new_new_n170_), .C(new_new_n76_), .Y(new_new_n173_));
  AOI210     g151(.A0(new_new_n173_), .A1(new_new_n169_), .B0(i_0_), .Y(new_new_n174_));
  NO2        g152(.A(new_new_n67_), .B(new_new_n61_), .Y(new_new_n175_));
  NA2        g153(.A(new_new_n175_), .B(new_new_n47_), .Y(new_new_n176_));
  NA2        g154(.A(new_new_n36_), .B(i_5_), .Y(new_new_n177_));
  NAi31      g155(.An(new_new_n177_), .B(new_new_n148_), .C(i_11_), .Y(new_new_n178_));
  NA2        g156(.A(i_3_), .B(i_5_), .Y(new_new_n179_));
  OR2        g157(.A(new_new_n179_), .B(new_new_n168_), .Y(new_new_n180_));
  AOI210     g158(.A0(new_new_n180_), .A1(new_new_n178_), .B0(new_new_n176_), .Y(new_new_n181_));
  NO2        g159(.A(new_new_n67_), .B(i_5_), .Y(new_new_n182_));
  NO2        g160(.A(i_13_), .B(i_10_), .Y(new_new_n183_));
  NA3        g161(.A(new_new_n183_), .B(new_new_n182_), .C(new_new_n45_), .Y(new_new_n184_));
  NO2        g162(.A(i_2_), .B(i_1_), .Y(new_new_n185_));
  NA2        g163(.A(new_new_n185_), .B(i_3_), .Y(new_new_n186_));
  NAi21      g164(.An(i_4_), .B(i_12_), .Y(new_new_n187_));
  NO3        g165(.A(new_new_n187_), .B(new_new_n186_), .C(new_new_n25_), .Y(new_new_n188_));
  NO3        g166(.A(new_new_n188_), .B(new_new_n181_), .C(new_new_n174_), .Y(new_new_n189_));
  INV        g167(.A(i_8_), .Y(new_new_n190_));
  NO2        g168(.A(new_new_n190_), .B(i_7_), .Y(new_new_n191_));
  NA2        g169(.A(new_new_n191_), .B(i_6_), .Y(new_new_n192_));
  NO3        g170(.A(i_3_), .B(new_new_n79_), .C(new_new_n49_), .Y(new_new_n193_));
  NA2        g171(.A(new_new_n193_), .B(new_new_n108_), .Y(new_new_n194_));
  NO3        g172(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n195_));
  NA3        g173(.A(new_new_n195_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n196_));
  NO3        g174(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n197_));
  OAI210     g175(.A0(new_new_n91_), .A1(i_12_), .B0(new_new_n197_), .Y(new_new_n198_));
  AOI210     g176(.A0(new_new_n198_), .A1(new_new_n196_), .B0(new_new_n194_), .Y(new_new_n199_));
  NO2        g177(.A(i_3_), .B(i_8_), .Y(new_new_n200_));
  NO3        g178(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n201_));
  NA3        g179(.A(new_new_n201_), .B(new_new_n200_), .C(new_new_n40_), .Y(new_new_n202_));
  NO2        g180(.A(new_new_n98_), .B(new_new_n58_), .Y(new_new_n203_));
  INV        g181(.A(new_new_n203_), .Y(new_new_n204_));
  NO2        g182(.A(i_13_), .B(i_9_), .Y(new_new_n205_));
  NA3        g183(.A(new_new_n205_), .B(i_6_), .C(new_new_n190_), .Y(new_new_n206_));
  NAi21      g184(.An(i_12_), .B(i_3_), .Y(new_new_n207_));
  OR2        g185(.A(new_new_n207_), .B(new_new_n206_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n45_), .B(i_5_), .Y(new_new_n209_));
  NO3        g187(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n210_));
  NA2        g188(.A(new_new_n210_), .B(i_10_), .Y(new_new_n211_));
  OAI220     g189(.A0(new_new_n211_), .A1(new_new_n208_), .B0(new_new_n204_), .B1(new_new_n202_), .Y(new_new_n212_));
  AOI210     g190(.A0(new_new_n212_), .A1(i_7_), .B0(new_new_n199_), .Y(new_new_n213_));
  OAI220     g191(.A0(new_new_n213_), .A1(i_4_), .B0(new_new_n192_), .B1(new_new_n189_), .Y(new_new_n214_));
  NAi21      g192(.An(i_12_), .B(i_7_), .Y(new_new_n215_));
  NA3        g193(.A(i_13_), .B(new_new_n190_), .C(i_10_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  NA2        g195(.A(i_0_), .B(i_5_), .Y(new_new_n218_));
  OAI220     g196(.A0(new_new_n79_), .A1(new_new_n186_), .B0(new_new_n176_), .B1(new_new_n129_), .Y(new_new_n219_));
  NAi31      g197(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n47_), .B(new_new_n61_), .Y(new_new_n221_));
  NA3        g199(.A(new_new_n221_), .B(i_0_), .C(i_4_), .Y(new_new_n222_));
  INV        g200(.A(i_13_), .Y(new_new_n223_));
  NO2        g201(.A(i_12_), .B(new_new_n223_), .Y(new_new_n224_));
  NA3        g202(.A(new_new_n224_), .B(new_new_n195_), .C(new_new_n193_), .Y(new_new_n225_));
  OAI210     g203(.A0(new_new_n222_), .A1(new_new_n220_), .B0(new_new_n225_), .Y(new_new_n226_));
  AOI220     g204(.A0(new_new_n226_), .A1(new_new_n138_), .B0(new_new_n219_), .B1(new_new_n217_), .Y(new_new_n227_));
  NO2        g205(.A(i_12_), .B(new_new_n37_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n179_), .B(i_4_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n229_), .B(new_new_n228_), .Y(new_new_n230_));
  OR2        g208(.A(i_8_), .B(i_7_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n231_), .B(new_new_n79_), .Y(new_new_n232_));
  NO2        g210(.A(new_new_n54_), .B(i_1_), .Y(new_new_n233_));
  NA2        g211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  INV        g212(.A(i_12_), .Y(new_new_n235_));
  NO3        g213(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n236_));
  NA2        g214(.A(i_2_), .B(i_1_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n234_), .B(new_new_n230_), .Y(new_new_n238_));
  NO3        g216(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n239_));
  NAi21      g217(.An(i_4_), .B(i_3_), .Y(new_new_n240_));
  NO2        g218(.A(i_0_), .B(i_6_), .Y(new_new_n241_));
  NOi41      g219(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n242_));
  NA2        g220(.A(new_new_n242_), .B(new_new_n241_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n237_), .B(new_new_n179_), .Y(new_new_n244_));
  NAi21      g222(.An(new_new_n243_), .B(new_new_n244_), .Y(new_new_n245_));
  INV        g223(.A(new_new_n245_), .Y(new_new_n246_));
  AOI220     g224(.A0(new_new_n246_), .A1(new_new_n40_), .B0(new_new_n238_), .B1(new_new_n205_), .Y(new_new_n247_));
  NO2        g225(.A(i_11_), .B(new_new_n223_), .Y(new_new_n248_));
  NOi21      g226(.An(i_1_), .B(i_6_), .Y(new_new_n249_));
  NAi21      g227(.An(i_3_), .B(i_7_), .Y(new_new_n250_));
  NO2        g228(.A(i_12_), .B(i_3_), .Y(new_new_n251_));
  NA3        g229(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n252_));
  INV        g230(.A(new_new_n139_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n235_), .B(i_13_), .Y(new_new_n254_));
  NO2        g232(.A(new_new_n254_), .B(new_new_n69_), .Y(new_new_n255_));
  NA2        g233(.A(new_new_n255_), .B(new_new_n253_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n231_), .B(new_new_n37_), .Y(new_new_n257_));
  NA2        g235(.A(i_12_), .B(i_6_), .Y(new_new_n258_));
  OR2        g236(.A(i_13_), .B(i_9_), .Y(new_new_n259_));
  NO3        g237(.A(new_new_n259_), .B(new_new_n258_), .C(new_new_n49_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n240_), .B(i_2_), .Y(new_new_n261_));
  NA3        g239(.A(new_new_n261_), .B(new_new_n260_), .C(new_new_n45_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n248_), .B(i_9_), .Y(new_new_n263_));
  NA2        g241(.A(i_0_), .B(new_new_n62_), .Y(new_new_n264_));
  OAI210     g242(.A0(new_new_n264_), .A1(new_new_n263_), .B0(new_new_n262_), .Y(new_new_n265_));
  NA2        g243(.A(new_new_n151_), .B(new_new_n61_), .Y(new_new_n266_));
  NO3        g244(.A(i_11_), .B(new_new_n223_), .C(new_new_n25_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n250_), .B(i_8_), .Y(new_new_n268_));
  NA3        g246(.A(i_5_), .B(new_new_n268_), .C(new_new_n267_), .Y(new_new_n269_));
  NO3        g247(.A(new_new_n26_), .B(new_new_n79_), .C(i_5_), .Y(new_new_n270_));
  NA3        g248(.A(new_new_n270_), .B(new_new_n257_), .C(new_new_n224_), .Y(new_new_n271_));
  AOI210     g249(.A0(new_new_n271_), .A1(new_new_n269_), .B0(new_new_n266_), .Y(new_new_n272_));
  AOI210     g250(.A0(new_new_n265_), .A1(new_new_n257_), .B0(new_new_n272_), .Y(new_new_n273_));
  NA4        g251(.A(new_new_n273_), .B(new_new_n256_), .C(new_new_n247_), .D(new_new_n227_), .Y(new_new_n274_));
  NO3        g252(.A(i_12_), .B(new_new_n223_), .C(new_new_n37_), .Y(new_new_n275_));
  INV        g253(.A(new_new_n275_), .Y(new_new_n276_));
  NO3        g254(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n277_));
  AOI220     g255(.A0(new_new_n277_), .A1(new_new_n193_), .B0(new_new_n160_), .B1(new_new_n233_), .Y(new_new_n278_));
  NO2        g256(.A(new_new_n278_), .B(new_new_n969_), .Y(new_new_n279_));
  NO3        g257(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n237_), .B(i_0_), .Y(new_new_n281_));
  AOI220     g259(.A0(new_new_n281_), .A1(new_new_n191_), .B0(new_new_n280_), .B1(new_new_n138_), .Y(new_new_n282_));
  NO2        g260(.A(i_3_), .B(new_new_n282_), .Y(new_new_n283_));
  NA2        g261(.A(i_0_), .B(i_1_), .Y(new_new_n284_));
  NO2        g262(.A(new_new_n284_), .B(i_2_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n59_), .B(i_6_), .Y(new_new_n286_));
  NA3        g264(.A(new_new_n286_), .B(new_new_n285_), .C(new_new_n160_), .Y(new_new_n287_));
  OAI210     g265(.A0(i_3_), .A1(new_new_n139_), .B0(new_new_n287_), .Y(new_new_n288_));
  NO3        g266(.A(new_new_n288_), .B(new_new_n283_), .C(new_new_n279_), .Y(new_new_n289_));
  NO2        g267(.A(i_3_), .B(i_10_), .Y(new_new_n290_));
  NA3        g268(.A(new_new_n290_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n291_));
  NO2        g269(.A(i_2_), .B(new_new_n96_), .Y(new_new_n292_));
  NOi21      g270(.An(new_new_n218_), .B(new_new_n98_), .Y(new_new_n293_));
  NA2        g271(.A(new_new_n293_), .B(new_new_n292_), .Y(new_new_n294_));
  AN2        g272(.A(i_3_), .B(i_10_), .Y(new_new_n295_));
  NA4        g273(.A(new_new_n295_), .B(new_new_n195_), .C(new_new_n172_), .D(new_new_n170_), .Y(new_new_n296_));
  NO2        g274(.A(i_5_), .B(new_new_n37_), .Y(new_new_n297_));
  NO2        g275(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n298_));
  OR2        g276(.A(new_new_n294_), .B(new_new_n291_), .Y(new_new_n299_));
  OAI220     g277(.A0(new_new_n299_), .A1(i_6_), .B0(new_new_n289_), .B1(new_new_n276_), .Y(new_new_n300_));
  NO4        g278(.A(new_new_n300_), .B(new_new_n274_), .C(new_new_n214_), .D(new_new_n164_), .Y(new_new_n301_));
  NO3        g279(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n302_));
  NA2        g280(.A(new_new_n281_), .B(i_8_), .Y(new_new_n303_));
  NO3        g281(.A(i_6_), .B(new_new_n190_), .C(i_7_), .Y(new_new_n304_));
  AOI210     g282(.A0(new_new_n971_), .A1(new_new_n303_), .B0(new_new_n165_), .Y(new_new_n305_));
  NO2        g283(.A(i_2_), .B(i_3_), .Y(new_new_n306_));
  OR2        g284(.A(i_0_), .B(i_5_), .Y(new_new_n307_));
  NA3        g285(.A(new_new_n232_), .B(new_new_n306_), .C(i_1_), .Y(new_new_n308_));
  NA3        g286(.A(new_new_n281_), .B(new_new_n160_), .C(new_new_n108_), .Y(new_new_n309_));
  NAi21      g287(.An(i_8_), .B(i_7_), .Y(new_new_n310_));
  NO2        g288(.A(new_new_n310_), .B(i_6_), .Y(new_new_n311_));
  NO2        g289(.A(new_new_n154_), .B(new_new_n47_), .Y(new_new_n312_));
  NA3        g290(.A(new_new_n312_), .B(new_new_n311_), .C(new_new_n160_), .Y(new_new_n313_));
  NA3        g291(.A(new_new_n313_), .B(new_new_n309_), .C(new_new_n308_), .Y(new_new_n314_));
  OAI210     g292(.A0(new_new_n314_), .A1(new_new_n305_), .B0(i_4_), .Y(new_new_n315_));
  NO2        g293(.A(i_12_), .B(i_10_), .Y(new_new_n316_));
  NOi21      g294(.An(i_5_), .B(i_0_), .Y(new_new_n317_));
  AOI210     g295(.A0(i_2_), .A1(new_new_n49_), .B0(new_new_n96_), .Y(new_new_n318_));
  NO3        g296(.A(new_new_n318_), .B(i_4_), .C(new_new_n124_), .Y(new_new_n319_));
  NA4        g297(.A(new_new_n77_), .B(new_new_n36_), .C(new_new_n79_), .D(i_8_), .Y(new_new_n320_));
  NA2        g298(.A(new_new_n319_), .B(new_new_n316_), .Y(new_new_n321_));
  NO2        g299(.A(i_6_), .B(i_8_), .Y(new_new_n322_));
  NO2        g300(.A(i_1_), .B(i_7_), .Y(new_new_n323_));
  AO220      g301(.A0(new_new_n323_), .A1(new_new_n322_), .B0(new_new_n311_), .B1(new_new_n233_), .Y(new_new_n324_));
  NA2        g302(.A(new_new_n324_), .B(new_new_n42_), .Y(new_new_n325_));
  NA3        g303(.A(new_new_n325_), .B(new_new_n321_), .C(new_new_n315_), .Y(new_new_n326_));
  NO3        g304(.A(new_new_n231_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n327_));
  NO3        g305(.A(new_new_n310_), .B(i_2_), .C(i_1_), .Y(new_new_n328_));
  OAI210     g306(.A0(new_new_n328_), .A1(new_new_n327_), .B0(i_6_), .Y(new_new_n329_));
  NA3        g307(.A(new_new_n249_), .B(new_new_n292_), .C(new_new_n190_), .Y(new_new_n330_));
  NA2        g308(.A(new_new_n330_), .B(new_new_n329_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n331_), .B(i_3_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n284_), .B(new_new_n75_), .Y(new_new_n333_));
  NA2        g311(.A(new_new_n333_), .B(new_new_n128_), .Y(new_new_n334_));
  NO2        g312(.A(new_new_n87_), .B(new_new_n190_), .Y(new_new_n335_));
  NA3        g313(.A(new_new_n293_), .B(new_new_n335_), .C(new_new_n61_), .Y(new_new_n336_));
  AOI210     g314(.A0(new_new_n336_), .A1(new_new_n334_), .B0(i_7_), .Y(new_new_n337_));
  NO2        g315(.A(new_new_n190_), .B(i_9_), .Y(new_new_n338_));
  NA2        g316(.A(new_new_n338_), .B(new_new_n203_), .Y(new_new_n339_));
  NO2        g317(.A(new_new_n337_), .B(new_new_n283_), .Y(new_new_n340_));
  AOI210     g318(.A0(new_new_n340_), .A1(new_new_n332_), .B0(new_new_n159_), .Y(new_new_n341_));
  AOI210     g319(.A0(new_new_n326_), .A1(new_new_n302_), .B0(new_new_n341_), .Y(new_new_n342_));
  NOi32      g320(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n343_));
  INV        g321(.A(new_new_n343_), .Y(new_new_n344_));
  NAi21      g322(.An(i_0_), .B(i_6_), .Y(new_new_n345_));
  NAi21      g323(.An(i_1_), .B(i_5_), .Y(new_new_n346_));
  NAi41      g324(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n347_));
  OAI220     g325(.A0(new_new_n347_), .A1(new_new_n346_), .B0(new_new_n220_), .B1(new_new_n156_), .Y(new_new_n348_));
  AOI210     g326(.A0(new_new_n347_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n349_));
  NOi32      g327(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n350_));
  NA2        g328(.A(new_new_n350_), .B(new_new_n47_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n351_), .B(i_0_), .Y(new_new_n352_));
  OR3        g330(.A(new_new_n352_), .B(new_new_n349_), .C(new_new_n348_), .Y(new_new_n353_));
  NO2        g331(.A(i_1_), .B(new_new_n96_), .Y(new_new_n354_));
  NAi21      g332(.An(i_3_), .B(i_4_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n355_), .B(i_9_), .Y(new_new_n356_));
  AN2        g334(.A(i_6_), .B(i_7_), .Y(new_new_n357_));
  OAI210     g335(.A0(new_new_n357_), .A1(new_new_n354_), .B0(new_new_n356_), .Y(new_new_n358_));
  NA2        g336(.A(i_2_), .B(i_7_), .Y(new_new_n359_));
  NO2        g337(.A(new_new_n355_), .B(i_10_), .Y(new_new_n360_));
  NA3        g338(.A(new_new_n360_), .B(new_new_n359_), .C(new_new_n241_), .Y(new_new_n361_));
  AOI210     g339(.A0(new_new_n361_), .A1(new_new_n358_), .B0(new_new_n182_), .Y(new_new_n362_));
  AOI210     g340(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n363_));
  OAI210     g341(.A0(new_new_n363_), .A1(new_new_n185_), .B0(new_new_n360_), .Y(new_new_n364_));
  AOI220     g342(.A0(new_new_n360_), .A1(new_new_n323_), .B0(new_new_n236_), .B1(new_new_n185_), .Y(new_new_n365_));
  AOI210     g343(.A0(new_new_n365_), .A1(new_new_n364_), .B0(i_5_), .Y(new_new_n366_));
  NO3        g344(.A(new_new_n366_), .B(new_new_n362_), .C(new_new_n353_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n367_), .B(new_new_n344_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n369_));
  AN2        g347(.A(i_12_), .B(i_5_), .Y(new_new_n370_));
  NO2        g348(.A(i_4_), .B(new_new_n26_), .Y(new_new_n371_));
  NA2        g349(.A(new_new_n371_), .B(new_new_n370_), .Y(new_new_n372_));
  NO2        g350(.A(i_11_), .B(i_6_), .Y(new_new_n373_));
  NA3        g351(.A(new_new_n373_), .B(new_new_n312_), .C(new_new_n223_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n374_), .B(new_new_n372_), .Y(new_new_n375_));
  NO2        g353(.A(new_new_n240_), .B(i_5_), .Y(new_new_n376_));
  NO2        g354(.A(i_5_), .B(i_10_), .Y(new_new_n377_));
  AOI220     g355(.A0(new_new_n377_), .A1(new_new_n261_), .B0(new_new_n376_), .B1(new_new_n195_), .Y(new_new_n378_));
  NA2        g356(.A(new_new_n140_), .B(new_new_n46_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(new_new_n378_), .Y(new_new_n380_));
  OAI210     g358(.A0(new_new_n380_), .A1(new_new_n375_), .B0(new_new_n369_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n382_));
  NO2        g360(.A(new_new_n146_), .B(new_new_n79_), .Y(new_new_n383_));
  OAI210     g361(.A0(new_new_n383_), .A1(new_new_n375_), .B0(new_new_n382_), .Y(new_new_n384_));
  NO3        g362(.A(new_new_n79_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n385_));
  NO2        g363(.A(i_11_), .B(i_12_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n377_), .B(new_new_n235_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n42_), .B(i_11_), .Y(new_new_n388_));
  OAI220     g366(.A0(new_new_n388_), .A1(new_new_n220_), .B0(new_new_n387_), .B1(new_new_n320_), .Y(new_new_n389_));
  NAi21      g367(.An(i_13_), .B(i_0_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n390_), .B(new_new_n237_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n389_), .B(new_new_n391_), .Y(new_new_n392_));
  NA3        g370(.A(new_new_n392_), .B(new_new_n384_), .C(new_new_n381_), .Y(new_new_n393_));
  NA2        g371(.A(new_new_n45_), .B(new_new_n223_), .Y(new_new_n394_));
  NO3        g372(.A(i_1_), .B(i_12_), .C(new_new_n79_), .Y(new_new_n395_));
  NO2        g373(.A(i_0_), .B(i_11_), .Y(new_new_n396_));
  INV        g374(.A(i_5_), .Y(new_new_n397_));
  AN2        g375(.A(i_1_), .B(i_6_), .Y(new_new_n398_));
  NOi21      g376(.An(i_2_), .B(i_12_), .Y(new_new_n399_));
  NA2        g377(.A(new_new_n399_), .B(new_new_n398_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n400_), .B(new_new_n397_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n138_), .B(i_9_), .Y(new_new_n402_));
  NO2        g380(.A(new_new_n402_), .B(i_4_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n401_), .B(new_new_n403_), .Y(new_new_n404_));
  OR2        g382(.A(i_13_), .B(i_10_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n168_), .B(new_new_n119_), .Y(new_new_n406_));
  OR2        g384(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n96_), .B(new_new_n25_), .Y(new_new_n408_));
  NA2        g386(.A(i_5_), .B(new_new_n210_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n409_), .B(new_new_n407_), .Y(new_new_n410_));
  INV        g388(.A(new_new_n410_), .Y(new_new_n411_));
  AOI210     g389(.A0(new_new_n411_), .A1(new_new_n404_), .B0(new_new_n26_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n309_), .B(new_new_n308_), .Y(new_new_n413_));
  AOI220     g391(.A0(new_new_n286_), .A1(new_new_n277_), .B0(new_new_n281_), .B1(i_8_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n414_), .B(new_new_n165_), .Y(new_new_n415_));
  NO2        g393(.A(new_new_n179_), .B(new_new_n79_), .Y(new_new_n416_));
  AOI220     g394(.A0(new_new_n416_), .A1(new_new_n285_), .B0(new_new_n270_), .B1(new_new_n210_), .Y(new_new_n417_));
  INV        g395(.A(new_new_n417_), .Y(new_new_n418_));
  NO3        g396(.A(new_new_n418_), .B(new_new_n415_), .C(new_new_n413_), .Y(new_new_n419_));
  INV        g397(.A(new_new_n91_), .Y(new_new_n420_));
  AOI210     g398(.A0(new_new_n154_), .A1(new_new_n420_), .B0(new_new_n310_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n286_), .B(new_new_n233_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n422_), .B(new_new_n179_), .Y(new_new_n423_));
  NO2        g401(.A(i_3_), .B(new_new_n49_), .Y(new_new_n424_));
  NA3        g402(.A(new_new_n323_), .B(new_new_n322_), .C(new_new_n424_), .Y(new_new_n425_));
  OAI210     g403(.A0(new_new_n190_), .A1(new_new_n186_), .B0(new_new_n425_), .Y(new_new_n426_));
  NO3        g404(.A(new_new_n426_), .B(new_new_n423_), .C(new_new_n421_), .Y(new_new_n427_));
  AOI210     g405(.A0(new_new_n427_), .A1(new_new_n419_), .B0(new_new_n263_), .Y(new_new_n428_));
  NO4        g406(.A(new_new_n428_), .B(new_new_n412_), .C(new_new_n393_), .D(new_new_n368_), .Y(new_new_n429_));
  NO2        g407(.A(new_new_n67_), .B(i_13_), .Y(new_new_n430_));
  NA3        g408(.A(new_new_n430_), .B(i_1_), .C(i_2_), .Y(new_new_n431_));
  NO2        g409(.A(i_10_), .B(i_9_), .Y(new_new_n432_));
  NAi21      g410(.An(i_12_), .B(i_8_), .Y(new_new_n433_));
  NO2        g411(.A(new_new_n433_), .B(i_3_), .Y(new_new_n434_));
  NA2        g412(.A(new_new_n434_), .B(new_new_n432_), .Y(new_new_n435_));
  NO2        g413(.A(new_new_n47_), .B(i_4_), .Y(new_new_n436_));
  NA2        g414(.A(new_new_n436_), .B(new_new_n99_), .Y(new_new_n437_));
  OAI220     g415(.A0(new_new_n437_), .A1(new_new_n202_), .B0(new_new_n435_), .B1(new_new_n431_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n298_), .B(i_0_), .Y(new_new_n439_));
  NO3        g417(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n258_), .B(new_new_n92_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n441_), .B(new_new_n440_), .Y(new_new_n442_));
  NA2        g420(.A(i_8_), .B(i_9_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n275_), .B(new_new_n203_), .Y(new_new_n444_));
  OAI220     g422(.A0(new_new_n444_), .A1(new_new_n443_), .B0(new_new_n442_), .B1(new_new_n439_), .Y(new_new_n445_));
  NA2        g423(.A(new_new_n248_), .B(new_new_n297_), .Y(new_new_n446_));
  NO3        g424(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n447_));
  INV        g425(.A(new_new_n447_), .Y(new_new_n448_));
  NA3        g426(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n449_));
  NA4        g427(.A(new_new_n141_), .B(new_new_n111_), .C(new_new_n74_), .D(new_new_n23_), .Y(new_new_n450_));
  OAI220     g428(.A0(new_new_n450_), .A1(new_new_n449_), .B0(new_new_n448_), .B1(new_new_n446_), .Y(new_new_n451_));
  NO3        g429(.A(new_new_n451_), .B(new_new_n445_), .C(new_new_n438_), .Y(new_new_n452_));
  NA2        g430(.A(new_new_n285_), .B(new_new_n103_), .Y(new_new_n453_));
  OR2        g431(.A(new_new_n453_), .B(new_new_n206_), .Y(new_new_n454_));
  OA220      g432(.A0(new_new_n339_), .A1(new_new_n159_), .B0(new_new_n454_), .B1(new_new_n230_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n91_), .B(i_13_), .Y(new_new_n456_));
  NA2        g434(.A(new_new_n416_), .B(new_new_n369_), .Y(new_new_n457_));
  NO2        g435(.A(i_2_), .B(i_13_), .Y(new_new_n458_));
  NA3        g436(.A(new_new_n458_), .B(new_new_n158_), .C(new_new_n94_), .Y(new_new_n459_));
  NO2        g437(.A(new_new_n457_), .B(new_new_n456_), .Y(new_new_n460_));
  NO2        g438(.A(i_6_), .B(i_7_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n461_), .B(i_5_), .Y(new_new_n462_));
  NO2        g440(.A(i_11_), .B(i_1_), .Y(new_new_n463_));
  OR2        g441(.A(i_11_), .B(i_8_), .Y(new_new_n464_));
  NOi21      g442(.An(i_2_), .B(i_7_), .Y(new_new_n465_));
  NAi31      g443(.An(new_new_n464_), .B(new_new_n465_), .C(i_0_), .Y(new_new_n466_));
  NO2        g444(.A(new_new_n405_), .B(i_6_), .Y(new_new_n467_));
  NA3        g445(.A(new_new_n467_), .B(i_1_), .C(new_new_n69_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n468_), .B(new_new_n466_), .Y(new_new_n469_));
  NO2        g447(.A(i_3_), .B(new_new_n190_), .Y(new_new_n470_));
  NO2        g448(.A(i_6_), .B(i_10_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n154_), .B(i_3_), .Y(new_new_n473_));
  NAi31      g451(.An(new_new_n472_), .B(new_new_n473_), .C(new_new_n224_), .Y(new_new_n474_));
  NA3        g452(.A(new_new_n382_), .B(new_new_n175_), .C(new_new_n145_), .Y(new_new_n475_));
  NA2        g453(.A(new_new_n475_), .B(new_new_n474_), .Y(new_new_n476_));
  NO3        g454(.A(new_new_n476_), .B(new_new_n469_), .C(new_new_n460_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n440_), .B(new_new_n370_), .Y(new_new_n478_));
  NA2        g456(.A(new_new_n447_), .B(new_new_n377_), .Y(new_new_n479_));
  NO2        g457(.A(new_new_n479_), .B(new_new_n222_), .Y(new_new_n480_));
  NAi21      g458(.An(new_new_n216_), .B(new_new_n386_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n323_), .B(new_new_n218_), .Y(new_new_n482_));
  NO2        g460(.A(new_new_n26_), .B(i_5_), .Y(new_new_n483_));
  NO2        g461(.A(i_0_), .B(new_new_n79_), .Y(new_new_n484_));
  NA3        g462(.A(new_new_n484_), .B(new_new_n483_), .C(new_new_n138_), .Y(new_new_n485_));
  OAI220     g463(.A0(new_new_n38_), .A1(new_new_n485_), .B0(new_new_n482_), .B1(new_new_n481_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n27_), .B(i_10_), .Y(new_new_n487_));
  NO2        g465(.A(new_new_n487_), .B(new_new_n456_), .Y(new_new_n488_));
  NA4        g466(.A(new_new_n295_), .B(new_new_n221_), .C(new_new_n67_), .D(new_new_n235_), .Y(new_new_n489_));
  NO2        g467(.A(new_new_n489_), .B(new_new_n462_), .Y(new_new_n490_));
  NO4        g468(.A(new_new_n490_), .B(new_new_n488_), .C(new_new_n486_), .D(new_new_n480_), .Y(new_new_n491_));
  NA4        g469(.A(new_new_n491_), .B(new_new_n477_), .C(new_new_n455_), .D(new_new_n452_), .Y(new_new_n492_));
  AN2        g470(.A(new_new_n277_), .B(new_new_n232_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n493_), .B(new_new_n172_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n118_), .B(new_new_n107_), .Y(new_new_n495_));
  AN2        g473(.A(new_new_n495_), .B(new_new_n440_), .Y(new_new_n496_));
  OAI210     g474(.A0(i_2_), .A1(new_new_n230_), .B0(new_new_n296_), .Y(new_new_n497_));
  AOI220     g475(.A0(new_new_n497_), .A1(new_new_n311_), .B0(new_new_n496_), .B1(new_new_n298_), .Y(new_new_n498_));
  NA4        g476(.A(new_new_n430_), .B(i_1_), .C(new_new_n200_), .D(i_2_), .Y(new_new_n499_));
  INV        g477(.A(new_new_n499_), .Y(new_new_n500_));
  NA2        g478(.A(new_new_n343_), .B(new_new_n67_), .Y(new_new_n501_));
  NA2        g479(.A(new_new_n357_), .B(new_new_n350_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n36_), .B(i_8_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n39_), .B(i_13_), .Y(new_new_n504_));
  INV        g482(.A(new_new_n504_), .Y(new_new_n505_));
  AOI210     g483(.A0(new_new_n500_), .A1(new_new_n201_), .B0(new_new_n505_), .Y(new_new_n506_));
  OAI210     g484(.A0(i_8_), .A1(new_new_n61_), .B0(new_new_n130_), .Y(new_new_n507_));
  AOI210     g485(.A0(new_new_n191_), .A1(i_9_), .B0(new_new_n257_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n508_), .B(new_new_n196_), .Y(new_new_n509_));
  AOI220     g487(.A0(i_6_), .A1(new_new_n509_), .B0(new_new_n507_), .B1(new_new_n406_), .Y(new_new_n510_));
  NA4        g488(.A(new_new_n510_), .B(new_new_n506_), .C(new_new_n498_), .D(new_new_n494_), .Y(new_new_n511_));
  INV        g489(.A(new_new_n376_), .Y(new_new_n512_));
  OAI210     g490(.A0(new_new_n372_), .A1(i_0_), .B0(new_new_n512_), .Y(new_new_n513_));
  NO2        g491(.A(i_12_), .B(new_new_n190_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n514_), .B(new_new_n223_), .Y(new_new_n515_));
  NO3        g493(.A(i_10_), .B(new_new_n515_), .C(new_new_n453_), .Y(new_new_n516_));
  NOi21      g494(.An(new_new_n304_), .B(new_new_n38_), .Y(new_new_n517_));
  OAI210     g495(.A0(new_new_n517_), .A1(new_new_n516_), .B0(new_new_n513_), .Y(new_new_n518_));
  NO2        g496(.A(i_8_), .B(i_7_), .Y(new_new_n519_));
  OAI210     g497(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n520_), .B(new_new_n221_), .Y(new_new_n521_));
  AOI220     g499(.A0(new_new_n312_), .A1(new_new_n40_), .B0(new_new_n233_), .B1(new_new_n205_), .Y(new_new_n522_));
  OAI220     g500(.A0(new_new_n522_), .A1(new_new_n179_), .B0(new_new_n521_), .B1(new_new_n240_), .Y(new_new_n523_));
  NO2        g501(.A(new_new_n974_), .B(i_6_), .Y(new_new_n524_));
  NA3        g502(.A(new_new_n524_), .B(new_new_n523_), .C(new_new_n519_), .Y(new_new_n525_));
  NA2        g503(.A(new_new_n416_), .B(new_new_n312_), .Y(new_new_n526_));
  OAI220     g504(.A0(new_new_n526_), .A1(new_new_n254_), .B0(new_new_n456_), .B1(new_new_n129_), .Y(new_new_n527_));
  NA2        g505(.A(new_new_n527_), .B(new_new_n257_), .Y(new_new_n528_));
  NOi31      g506(.An(new_new_n281_), .B(new_new_n291_), .C(new_new_n177_), .Y(new_new_n529_));
  NA3        g507(.A(new_new_n295_), .B(new_new_n170_), .C(new_new_n91_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n154_), .B(i_5_), .Y(new_new_n531_));
  NA3        g509(.A(new_new_n531_), .B(new_new_n394_), .C(new_new_n306_), .Y(new_new_n532_));
  INV        g510(.A(new_new_n532_), .Y(new_new_n533_));
  OAI210     g511(.A0(new_new_n533_), .A1(new_new_n529_), .B0(new_new_n447_), .Y(new_new_n534_));
  NA4        g512(.A(new_new_n534_), .B(new_new_n528_), .C(new_new_n525_), .D(new_new_n518_), .Y(new_new_n535_));
  NA2        g513(.A(new_new_n275_), .B(new_new_n77_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n334_), .B(new_new_n536_), .Y(new_new_n537_));
  INV        g515(.A(new_new_n277_), .Y(new_new_n538_));
  NO2        g516(.A(new_new_n538_), .B(new_new_n169_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n47_), .B(new_new_n354_), .Y(new_new_n540_));
  NA2        g518(.A(new_new_n514_), .B(new_new_n267_), .Y(new_new_n541_));
  NO2        g519(.A(new_new_n540_), .B(new_new_n541_), .Y(new_new_n542_));
  NO3        g520(.A(new_new_n542_), .B(new_new_n539_), .C(new_new_n537_), .Y(new_new_n543_));
  NO3        g521(.A(new_new_n43_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n544_));
  NO3        g522(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n231_), .B(new_new_n36_), .Y(new_new_n546_));
  AN2        g524(.A(new_new_n546_), .B(new_new_n545_), .Y(new_new_n547_));
  OA210      g525(.A0(new_new_n547_), .A1(new_new_n544_), .B0(new_new_n343_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n405_), .B(i_1_), .Y(new_new_n549_));
  NOi31      g527(.An(new_new_n549_), .B(new_new_n441_), .C(new_new_n67_), .Y(new_new_n550_));
  AN4        g528(.A(new_new_n550_), .B(new_new_n403_), .C(new_new_n483_), .D(i_2_), .Y(new_new_n551_));
  NO2        g529(.A(new_new_n414_), .B(new_new_n173_), .Y(new_new_n552_));
  NO3        g530(.A(new_new_n552_), .B(new_new_n551_), .C(new_new_n548_), .Y(new_new_n553_));
  NOi21      g531(.An(i_10_), .B(i_6_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n79_), .B(new_new_n25_), .Y(new_new_n555_));
  AOI220     g533(.A0(new_new_n275_), .A1(new_new_n555_), .B0(new_new_n267_), .B1(new_new_n554_), .Y(new_new_n556_));
  NO2        g534(.A(new_new_n556_), .B(new_new_n439_), .Y(new_new_n557_));
  NO2        g535(.A(new_new_n110_), .B(new_new_n23_), .Y(new_new_n558_));
  NA2        g536(.A(new_new_n304_), .B(new_new_n161_), .Y(new_new_n559_));
  AOI220     g537(.A0(new_new_n559_), .A1(new_new_n422_), .B0(new_new_n180_), .B1(new_new_n178_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n195_), .B(new_new_n37_), .Y(new_new_n561_));
  NOi31      g539(.An(new_new_n142_), .B(new_new_n561_), .C(new_new_n320_), .Y(new_new_n562_));
  NO3        g540(.A(new_new_n562_), .B(new_new_n560_), .C(new_new_n557_), .Y(new_new_n563_));
  NO2        g541(.A(new_new_n501_), .B(new_new_n365_), .Y(new_new_n564_));
  INV        g542(.A(new_new_n306_), .Y(new_new_n565_));
  NA2        g543(.A(new_new_n973_), .B(new_new_n267_), .Y(new_new_n566_));
  NA3        g544(.A(new_new_n373_), .B(new_new_n275_), .C(new_new_n218_), .Y(new_new_n567_));
  AOI210     g545(.A0(new_new_n567_), .A1(new_new_n566_), .B0(new_new_n565_), .Y(new_new_n568_));
  NO3        g546(.A(i_4_), .B(new_new_n329_), .C(new_new_n291_), .Y(new_new_n569_));
  OR2        g547(.A(i_2_), .B(i_5_), .Y(new_new_n570_));
  BUFFER     g548(.A(new_new_n570_), .Y(new_new_n571_));
  NO3        g549(.A(new_new_n569_), .B(new_new_n568_), .C(new_new_n564_), .Y(new_new_n572_));
  NA4        g550(.A(new_new_n572_), .B(new_new_n563_), .C(new_new_n553_), .D(new_new_n543_), .Y(new_new_n573_));
  NO4        g551(.A(new_new_n573_), .B(new_new_n535_), .C(new_new_n511_), .D(new_new_n492_), .Y(new_new_n574_));
  NA4        g552(.A(new_new_n574_), .B(new_new_n429_), .C(new_new_n342_), .D(new_new_n301_), .Y(men7));
  NO2        g553(.A(new_new_n103_), .B(new_new_n84_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n371_), .B(new_new_n576_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n471_), .B(new_new_n77_), .Y(new_new_n578_));
  NA2        g556(.A(i_11_), .B(new_new_n190_), .Y(new_new_n579_));
  OAI210     g557(.A0(new_new_n970_), .A1(new_new_n578_), .B0(new_new_n577_), .Y(new_new_n580_));
  NA3        g558(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n235_), .B(i_4_), .Y(new_new_n582_));
  NA2        g560(.A(new_new_n582_), .B(i_8_), .Y(new_new_n583_));
  NO2        g561(.A(new_new_n100_), .B(new_new_n581_), .Y(new_new_n584_));
  NA2        g562(.A(i_2_), .B(new_new_n79_), .Y(new_new_n585_));
  OAI210     g563(.A0(new_new_n82_), .A1(new_new_n200_), .B0(new_new_n201_), .Y(new_new_n586_));
  NO2        g564(.A(i_7_), .B(new_new_n37_), .Y(new_new_n587_));
  NA2        g565(.A(i_4_), .B(i_8_), .Y(new_new_n588_));
  AOI210     g566(.A0(new_new_n588_), .A1(new_new_n295_), .B0(new_new_n587_), .Y(new_new_n589_));
  OAI220     g567(.A0(new_new_n589_), .A1(new_new_n585_), .B0(new_new_n586_), .B1(i_13_), .Y(new_new_n590_));
  NO3        g568(.A(new_new_n590_), .B(new_new_n584_), .C(new_new_n580_), .Y(new_new_n591_));
  AOI210     g569(.A0(new_new_n124_), .A1(new_new_n60_), .B0(i_10_), .Y(new_new_n592_));
  AOI210     g570(.A0(new_new_n592_), .A1(new_new_n235_), .B0(new_new_n158_), .Y(new_new_n593_));
  NO2        g571(.A(i_10_), .B(new_new_n23_), .Y(new_new_n594_));
  OR3        g572(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n595_));
  NO3        g573(.A(new_new_n595_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n596_));
  INV        g574(.A(new_new_n197_), .Y(new_new_n597_));
  OA220      g575(.A0(new_new_n595_), .A1(new_new_n565_), .B0(new_new_n593_), .B1(new_new_n259_), .Y(new_new_n598_));
  AOI210     g576(.A0(new_new_n598_), .A1(new_new_n591_), .B0(new_new_n61_), .Y(new_new_n599_));
  NOi21      g577(.An(i_11_), .B(i_7_), .Y(new_new_n600_));
  AO210      g578(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n601_));
  NO2        g579(.A(new_new_n601_), .B(new_new_n600_), .Y(new_new_n602_));
  NA3        g580(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n603_), .B(new_new_n61_), .Y(new_new_n604_));
  AO210      g582(.A0(new_new_n80_), .A1(new_new_n365_), .B0(new_new_n41_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n61_), .B(new_new_n977_), .Y(new_new_n606_));
  NA2        g584(.A(new_new_n606_), .B(new_new_n605_), .Y(new_new_n607_));
  OAI210     g585(.A0(new_new_n607_), .A1(new_new_n604_), .B0(i_6_), .Y(new_new_n608_));
  NO2        g586(.A(i_6_), .B(i_11_), .Y(new_new_n609_));
  NO4        g587(.A(new_new_n215_), .B(new_new_n124_), .C(i_13_), .D(new_new_n79_), .Y(new_new_n610_));
  NA3        g588(.A(new_new_n519_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n134_), .B(i_9_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n612_), .B(new_new_n964_), .Y(new_new_n613_));
  NA3        g591(.A(i_1_), .B(new_new_n306_), .C(i_6_), .Y(new_new_n614_));
  AOI210     g592(.A0(new_new_n463_), .A1(new_new_n408_), .B0(new_new_n239_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n615_), .B(new_new_n585_), .Y(new_new_n616_));
  NAi21      g594(.An(new_new_n611_), .B(new_new_n86_), .Y(new_new_n617_));
  NO2        g595(.A(i_11_), .B(new_new_n37_), .Y(new_new_n618_));
  NA2        g596(.A(new_new_n618_), .B(new_new_n24_), .Y(new_new_n619_));
  OAI210     g597(.A0(new_new_n619_), .A1(i_6_), .B0(new_new_n617_), .Y(new_new_n620_));
  OR3        g598(.A(new_new_n620_), .B(new_new_n616_), .C(new_new_n613_), .Y(new_new_n621_));
  NO2        g599(.A(new_new_n621_), .B(new_new_n610_), .Y(new_new_n622_));
  NA2        g600(.A(i_3_), .B(new_new_n190_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n113_), .B(new_new_n37_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n79_), .B(i_9_), .Y(new_new_n625_));
  NA2        g603(.A(i_1_), .B(i_3_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n622_), .B(new_new_n608_), .Y(new_new_n627_));
  NO3        g605(.A(new_new_n464_), .B(i_3_), .C(i_7_), .Y(new_new_n628_));
  OA210      g606(.A0(new_new_n628_), .A1(new_new_n242_), .B0(new_new_n79_), .Y(new_new_n629_));
  NA3        g607(.A(new_new_n471_), .B(new_new_n503_), .C(new_new_n47_), .Y(new_new_n630_));
  NO3        g608(.A(new_new_n465_), .B(new_new_n588_), .C(new_new_n79_), .Y(new_new_n631_));
  NA2        g609(.A(new_new_n631_), .B(new_new_n25_), .Y(new_new_n632_));
  NA3        g610(.A(new_new_n158_), .B(new_new_n77_), .C(new_new_n79_), .Y(new_new_n633_));
  NA3        g611(.A(new_new_n633_), .B(new_new_n632_), .C(new_new_n630_), .Y(new_new_n634_));
  OAI210     g612(.A0(new_new_n634_), .A1(new_new_n629_), .B0(i_1_), .Y(new_new_n635_));
  AOI210     g613(.A0(new_new_n258_), .A1(new_new_n92_), .B0(i_1_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n355_), .B(i_2_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n637_), .B(new_new_n636_), .Y(new_new_n638_));
  NA2        g616(.A(new_new_n614_), .B(new_new_n638_), .Y(new_new_n639_));
  INV        g617(.A(new_new_n639_), .Y(new_new_n640_));
  AOI210     g618(.A0(new_new_n640_), .A1(new_new_n635_), .B0(i_13_), .Y(new_new_n641_));
  OR2        g619(.A(i_11_), .B(i_7_), .Y(new_new_n642_));
  NA2        g620(.A(new_new_n101_), .B(new_new_n134_), .Y(new_new_n643_));
  AOI220     g621(.A0(new_new_n458_), .A1(new_new_n158_), .B0(new_new_n436_), .B1(new_new_n134_), .Y(new_new_n644_));
  OAI210     g622(.A0(new_new_n644_), .A1(new_new_n45_), .B0(new_new_n643_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n55_), .B(i_12_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n465_), .B(new_new_n24_), .Y(new_new_n647_));
  NO2        g625(.A(new_new_n963_), .B(new_new_n87_), .Y(new_new_n648_));
  AOI210     g626(.A0(new_new_n645_), .A1(new_new_n322_), .B0(new_new_n648_), .Y(new_new_n649_));
  AOI220     g627(.A0(i_12_), .A1(new_new_n66_), .B0(new_new_n373_), .B1(new_new_n975_), .Y(new_new_n650_));
  NO2        g628(.A(new_new_n650_), .B(new_new_n240_), .Y(new_new_n651_));
  AOI210     g629(.A0(new_new_n433_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n652_));
  NOi31      g630(.An(new_new_n652_), .B(new_new_n578_), .C(new_new_n45_), .Y(new_new_n653_));
  NA2        g631(.A(new_new_n123_), .B(i_13_), .Y(new_new_n654_));
  NO2        g632(.A(new_new_n654_), .B(new_new_n636_), .Y(new_new_n655_));
  NO3        g633(.A(new_new_n65_), .B(new_new_n32_), .C(new_new_n96_), .Y(new_new_n656_));
  NA2        g634(.A(new_new_n26_), .B(new_new_n190_), .Y(new_new_n657_));
  NA2        g635(.A(new_new_n657_), .B(i_7_), .Y(new_new_n658_));
  NO3        g636(.A(new_new_n465_), .B(new_new_n235_), .C(new_new_n79_), .Y(new_new_n659_));
  AOI210     g637(.A0(new_new_n659_), .A1(new_new_n658_), .B0(new_new_n656_), .Y(new_new_n660_));
  AOI220     g638(.A0(new_new_n373_), .A1(new_new_n975_), .B0(new_new_n86_), .B1(new_new_n97_), .Y(new_new_n661_));
  OAI220     g639(.A0(new_new_n661_), .A1(new_new_n583_), .B0(new_new_n660_), .B1(new_new_n597_), .Y(new_new_n662_));
  NO4        g640(.A(new_new_n662_), .B(new_new_n655_), .C(new_new_n653_), .D(new_new_n651_), .Y(new_new_n663_));
  NA2        g641(.A(new_new_n609_), .B(i_13_), .Y(new_new_n664_));
  NAi21      g642(.An(i_11_), .B(i_12_), .Y(new_new_n665_));
  NA2        g643(.A(new_new_n972_), .B(new_new_n302_), .Y(new_new_n666_));
  NA2        g644(.A(new_new_n666_), .B(new_new_n664_), .Y(new_new_n667_));
  NA2        g645(.A(new_new_n667_), .B(new_new_n61_), .Y(new_new_n668_));
  NO2        g646(.A(i_2_), .B(i_12_), .Y(new_new_n669_));
  NA2        g647(.A(new_new_n354_), .B(new_new_n669_), .Y(new_new_n670_));
  NA2        g648(.A(i_8_), .B(new_new_n25_), .Y(new_new_n671_));
  NO3        g649(.A(new_new_n671_), .B(new_new_n371_), .C(new_new_n582_), .Y(new_new_n672_));
  OAI210     g650(.A0(new_new_n672_), .A1(new_new_n356_), .B0(new_new_n354_), .Y(new_new_n673_));
  NA2        g651(.A(new_new_n673_), .B(new_new_n670_), .Y(new_new_n674_));
  NA3        g652(.A(new_new_n674_), .B(new_new_n46_), .C(new_new_n223_), .Y(new_new_n675_));
  NA4        g653(.A(new_new_n675_), .B(new_new_n668_), .C(new_new_n663_), .D(new_new_n649_), .Y(new_new_n676_));
  OR4        g654(.A(new_new_n676_), .B(new_new_n641_), .C(new_new_n627_), .D(new_new_n599_), .Y(men5));
  AN2        g655(.A(new_new_n24_), .B(i_10_), .Y(new_new_n678_));
  NA3        g656(.A(new_new_n678_), .B(new_new_n669_), .C(new_new_n103_), .Y(new_new_n679_));
  NO2        g657(.A(new_new_n583_), .B(i_11_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n82_), .B(new_new_n680_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n681_), .B(new_new_n679_), .Y(new_new_n682_));
  NO3        g660(.A(i_11_), .B(new_new_n235_), .C(i_13_), .Y(new_new_n683_));
  NO2        g661(.A(new_new_n120_), .B(new_new_n23_), .Y(new_new_n684_));
  NA2        g662(.A(i_12_), .B(i_8_), .Y(new_new_n685_));
  OAI210     g663(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n685_), .Y(new_new_n686_));
  INV        g664(.A(new_new_n432_), .Y(new_new_n687_));
  AOI220     g665(.A0(new_new_n306_), .A1(new_new_n558_), .B0(new_new_n686_), .B1(new_new_n684_), .Y(new_new_n688_));
  INV        g666(.A(new_new_n688_), .Y(new_new_n689_));
  NO2        g667(.A(new_new_n689_), .B(new_new_n682_), .Y(new_new_n690_));
  INV        g668(.A(new_new_n167_), .Y(new_new_n691_));
  OAI210     g669(.A0(new_new_n637_), .A1(new_new_n434_), .B0(new_new_n106_), .Y(new_new_n692_));
  NO2        g670(.A(new_new_n692_), .B(new_new_n691_), .Y(new_new_n693_));
  NO2        g671(.A(new_new_n443_), .B(new_new_n26_), .Y(new_new_n694_));
  NO2        g672(.A(new_new_n187_), .B(new_new_n121_), .Y(new_new_n695_));
  OAI210     g673(.A0(new_new_n695_), .A1(new_new_n684_), .B0(i_2_), .Y(new_new_n696_));
  INV        g674(.A(new_new_n168_), .Y(new_new_n697_));
  NO3        g675(.A(new_new_n601_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n698_));
  AOI210     g676(.A0(new_new_n697_), .A1(new_new_n82_), .B0(new_new_n698_), .Y(new_new_n699_));
  AOI210     g677(.A0(new_new_n699_), .A1(new_new_n696_), .B0(new_new_n190_), .Y(new_new_n700_));
  OA210      g678(.A0(new_new_n602_), .A1(new_new_n122_), .B0(i_13_), .Y(new_new_n701_));
  NA2        g679(.A(new_new_n197_), .B(new_new_n200_), .Y(new_new_n702_));
  NA2        g680(.A(new_new_n148_), .B(new_new_n579_), .Y(new_new_n703_));
  AOI210     g681(.A0(new_new_n703_), .A1(new_new_n702_), .B0(new_new_n359_), .Y(new_new_n704_));
  AOI210     g682(.A0(new_new_n207_), .A1(new_new_n144_), .B0(new_new_n503_), .Y(new_new_n705_));
  NA2        g683(.A(new_new_n705_), .B(new_new_n408_), .Y(new_new_n706_));
  NO2        g684(.A(new_new_n97_), .B(new_new_n45_), .Y(new_new_n707_));
  INV        g685(.A(new_new_n292_), .Y(new_new_n708_));
  NA4        g686(.A(new_new_n708_), .B(new_new_n295_), .C(new_new_n120_), .D(new_new_n43_), .Y(new_new_n709_));
  OAI210     g687(.A0(new_new_n709_), .A1(new_new_n707_), .B0(new_new_n706_), .Y(new_new_n710_));
  NO4        g688(.A(new_new_n710_), .B(new_new_n704_), .C(new_new_n701_), .D(new_new_n700_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n558_), .B(new_new_n28_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n683_), .B(new_new_n268_), .Y(new_new_n713_));
  NA2        g691(.A(new_new_n713_), .B(new_new_n712_), .Y(new_new_n714_));
  NO2        g692(.A(new_new_n60_), .B(i_12_), .Y(new_new_n715_));
  NO2        g693(.A(new_new_n715_), .B(new_new_n122_), .Y(new_new_n716_));
  NO2        g694(.A(new_new_n716_), .B(new_new_n579_), .Y(new_new_n717_));
  AOI220     g695(.A0(new_new_n717_), .A1(new_new_n36_), .B0(new_new_n714_), .B1(new_new_n47_), .Y(new_new_n718_));
  NA4        g696(.A(new_new_n718_), .B(new_new_n711_), .C(new_new_n976_), .D(new_new_n690_), .Y(men6));
  NO3        g697(.A(i_9_), .B(new_new_n297_), .C(i_1_), .Y(new_new_n720_));
  NO2        g698(.A(new_new_n182_), .B(new_new_n135_), .Y(new_new_n721_));
  OAI210     g699(.A0(new_new_n721_), .A1(new_new_n720_), .B0(new_new_n967_), .Y(new_new_n722_));
  NA4        g700(.A(new_new_n377_), .B(new_new_n470_), .C(new_new_n65_), .D(new_new_n96_), .Y(new_new_n723_));
  INV        g701(.A(new_new_n723_), .Y(new_new_n724_));
  NO2        g702(.A(new_new_n220_), .B(new_new_n472_), .Y(new_new_n725_));
  NO2        g703(.A(i_11_), .B(i_9_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n724_), .B(new_new_n317_), .Y(new_new_n727_));
  AO210      g705(.A0(new_new_n727_), .A1(new_new_n722_), .B0(i_12_), .Y(new_new_n728_));
  NA2        g706(.A(new_new_n360_), .B(new_new_n323_), .Y(new_new_n729_));
  NA2        g707(.A(new_new_n628_), .B(new_new_n65_), .Y(new_new_n730_));
  NA3        g708(.A(new_new_n80_), .B(new_new_n730_), .C(new_new_n729_), .Y(new_new_n731_));
  INV        g709(.A(new_new_n194_), .Y(new_new_n732_));
  AOI220     g710(.A0(new_new_n732_), .A1(new_new_n726_), .B0(new_new_n731_), .B1(new_new_n67_), .Y(new_new_n733_));
  INV        g711(.A(new_new_n316_), .Y(new_new_n734_));
  NA2        g712(.A(new_new_n69_), .B(new_new_n127_), .Y(new_new_n735_));
  NA2        g713(.A(new_new_n25_), .B(new_new_n47_), .Y(new_new_n736_));
  AOI210     g714(.A0(new_new_n736_), .A1(new_new_n735_), .B0(new_new_n734_), .Y(new_new_n737_));
  NO2        g715(.A(new_new_n32_), .B(i_11_), .Y(new_new_n738_));
  NA3        g716(.A(new_new_n738_), .B(new_new_n461_), .C(new_new_n377_), .Y(new_new_n739_));
  OAI210     g717(.A0(new_new_n628_), .A1(new_new_n546_), .B0(new_new_n545_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n740_), .B(new_new_n739_), .Y(new_new_n741_));
  OR2        g719(.A(new_new_n741_), .B(new_new_n737_), .Y(new_new_n742_));
  NO2        g720(.A(new_new_n642_), .B(i_2_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n37_), .B(new_new_n743_), .Y(new_new_n744_));
  NA3        g722(.A(new_new_n338_), .B(new_new_n251_), .C(i_7_), .Y(new_new_n745_));
  BUFFER     g723(.A(new_new_n602_), .Y(new_new_n746_));
  NA2        g724(.A(new_new_n746_), .B(new_new_n143_), .Y(new_new_n747_));
  AO210      g725(.A0(new_new_n479_), .A1(new_new_n687_), .B0(new_new_n36_), .Y(new_new_n748_));
  NA4        g726(.A(new_new_n748_), .B(new_new_n747_), .C(new_new_n745_), .D(new_new_n744_), .Y(new_new_n749_));
  OAI210     g727(.A0(i_6_), .A1(i_11_), .B0(new_new_n80_), .Y(new_new_n750_));
  AOI220     g728(.A0(new_new_n750_), .A1(new_new_n545_), .B0(new_new_n725_), .B1(new_new_n658_), .Y(new_new_n751_));
  NA3        g729(.A(new_new_n359_), .B(new_new_n236_), .C(new_new_n143_), .Y(new_new_n752_));
  NA2        g730(.A(new_new_n385_), .B(new_new_n64_), .Y(new_new_n753_));
  NA3        g731(.A(new_new_n753_), .B(new_new_n752_), .C(new_new_n751_), .Y(new_new_n754_));
  AO210      g732(.A0(new_new_n503_), .A1(new_new_n47_), .B0(new_new_n81_), .Y(new_new_n755_));
  NA3        g733(.A(new_new_n755_), .B(new_new_n471_), .C(new_new_n218_), .Y(new_new_n756_));
  INV        g734(.A(new_new_n544_), .Y(new_new_n757_));
  NA2        g735(.A(new_new_n107_), .B(new_new_n396_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n241_), .B(new_new_n47_), .Y(new_new_n759_));
  INV        g737(.A(new_new_n571_), .Y(new_new_n760_));
  NA3        g738(.A(new_new_n760_), .B(new_new_n316_), .C(i_7_), .Y(new_new_n761_));
  NA4        g739(.A(new_new_n761_), .B(new_new_n758_), .C(new_new_n757_), .D(new_new_n756_), .Y(new_new_n762_));
  NO4        g740(.A(new_new_n762_), .B(new_new_n754_), .C(new_new_n749_), .D(new_new_n742_), .Y(new_new_n763_));
  NA4        g741(.A(new_new_n763_), .B(new_new_n733_), .C(new_new_n728_), .D(new_new_n367_), .Y(men3));
  NA2        g742(.A(i_6_), .B(i_7_), .Y(new_new_n765_));
  NO2        g743(.A(new_new_n765_), .B(i_0_), .Y(new_new_n766_));
  NO2        g744(.A(i_11_), .B(new_new_n235_), .Y(new_new_n767_));
  OAI210     g745(.A0(new_new_n766_), .A1(new_new_n281_), .B0(new_new_n767_), .Y(new_new_n768_));
  NO2        g746(.A(new_new_n768_), .B(new_new_n190_), .Y(new_new_n769_));
  NO3        g747(.A(new_new_n439_), .B(new_new_n84_), .C(new_new_n45_), .Y(new_new_n770_));
  OA210      g748(.A0(new_new_n770_), .A1(new_new_n769_), .B0(new_new_n170_), .Y(new_new_n771_));
  NA3        g749(.A(new_new_n752_), .B(new_new_n586_), .C(new_new_n358_), .Y(new_new_n772_));
  NA2        g750(.A(new_new_n772_), .B(new_new_n40_), .Y(new_new_n773_));
  AN2        g751(.A(new_new_n441_), .B(new_new_n56_), .Y(new_new_n774_));
  AOI210     g752(.A0(new_new_n965_), .A1(new_new_n773_), .B0(new_new_n49_), .Y(new_new_n775_));
  NO4        g753(.A(new_new_n363_), .B(new_new_n370_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n776_));
  NA2        g754(.A(new_new_n182_), .B(new_new_n554_), .Y(new_new_n777_));
  NOi21      g755(.An(new_new_n777_), .B(new_new_n776_), .Y(new_new_n778_));
  NA2        g756(.A(new_new_n652_), .B(new_new_n625_), .Y(new_new_n779_));
  NA2        g757(.A(i_0_), .B(new_new_n424_), .Y(new_new_n780_));
  OAI220     g758(.A0(new_new_n780_), .A1(new_new_n779_), .B0(new_new_n778_), .B1(new_new_n61_), .Y(new_new_n781_));
  NOi21      g759(.An(i_5_), .B(i_9_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n782_), .B(new_new_n430_), .Y(new_new_n783_));
  NO3        g761(.A(new_new_n402_), .B(new_new_n258_), .C(new_new_n67_), .Y(new_new_n784_));
  INV        g762(.A(new_new_n784_), .Y(new_new_n785_));
  OAI220     g763(.A0(new_new_n785_), .A1(new_new_n177_), .B0(new_new_n588_), .B1(new_new_n783_), .Y(new_new_n786_));
  NO4        g764(.A(new_new_n786_), .B(new_new_n781_), .C(new_new_n775_), .D(new_new_n771_), .Y(new_new_n787_));
  NA2        g765(.A(new_new_n182_), .B(new_new_n24_), .Y(new_new_n788_));
  NO2        g766(.A(new_new_n624_), .B(new_new_n576_), .Y(new_new_n789_));
  NO2        g767(.A(new_new_n789_), .B(new_new_n788_), .Y(new_new_n790_));
  NA2        g768(.A(new_new_n302_), .B(new_new_n125_), .Y(new_new_n791_));
  NAi21      g769(.An(new_new_n159_), .B(new_new_n424_), .Y(new_new_n792_));
  OAI220     g770(.A0(new_new_n792_), .A1(new_new_n759_), .B0(new_new_n791_), .B1(new_new_n387_), .Y(new_new_n793_));
  NO2        g771(.A(new_new_n793_), .B(new_new_n790_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n555_), .B(i_0_), .Y(new_new_n795_));
  NO3        g773(.A(new_new_n795_), .B(new_new_n372_), .C(new_new_n82_), .Y(new_new_n796_));
  NO3        g774(.A(new_new_n570_), .B(new_new_n215_), .C(new_new_n405_), .Y(new_new_n797_));
  AOI210     g775(.A0(new_new_n797_), .A1(i_11_), .B0(new_new_n796_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n683_), .B(new_new_n317_), .Y(new_new_n799_));
  NO2        g777(.A(new_new_n619_), .B(new_new_n521_), .Y(new_new_n800_));
  NA2        g778(.A(i_0_), .B(i_10_), .Y(new_new_n801_));
  NO4        g779(.A(new_new_n110_), .B(new_new_n58_), .C(new_new_n623_), .D(i_5_), .Y(new_new_n802_));
  AN2        g780(.A(new_new_n802_), .B(new_new_n45_), .Y(new_new_n803_));
  NA2        g781(.A(new_new_n182_), .B(new_new_n77_), .Y(new_new_n804_));
  NA2        g782(.A(new_new_n549_), .B(i_4_), .Y(new_new_n805_));
  NA2        g783(.A(new_new_n185_), .B(new_new_n200_), .Y(new_new_n806_));
  OAI220     g784(.A0(new_new_n806_), .A1(new_new_n799_), .B0(new_new_n805_), .B1(new_new_n804_), .Y(new_new_n807_));
  NO3        g785(.A(new_new_n807_), .B(new_new_n803_), .C(new_new_n800_), .Y(new_new_n808_));
  NA3        g786(.A(new_new_n808_), .B(new_new_n798_), .C(new_new_n794_), .Y(new_new_n809_));
  NA2        g787(.A(i_11_), .B(i_9_), .Y(new_new_n810_));
  NO3        g788(.A(i_12_), .B(new_new_n810_), .C(new_new_n585_), .Y(new_new_n811_));
  AN2        g789(.A(new_new_n811_), .B(i_0_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n49_), .B(i_7_), .Y(new_new_n813_));
  NA2        g791(.A(new_new_n382_), .B(new_new_n175_), .Y(new_new_n814_));
  NA2        g792(.A(new_new_n814_), .B(new_new_n157_), .Y(new_new_n815_));
  NO2        g793(.A(new_new_n810_), .B(new_new_n67_), .Y(new_new_n816_));
  NO2        g794(.A(new_new_n171_), .B(i_0_), .Y(new_new_n817_));
  INV        g795(.A(new_new_n817_), .Y(new_new_n818_));
  NA2        g796(.A(new_new_n461_), .B(new_new_n229_), .Y(new_new_n819_));
  AOI210     g797(.A0(new_new_n357_), .A1(new_new_n42_), .B0(new_new_n395_), .Y(new_new_n820_));
  OAI220     g798(.A0(new_new_n820_), .A1(new_new_n783_), .B0(new_new_n819_), .B1(new_new_n818_), .Y(new_new_n821_));
  NO3        g799(.A(new_new_n821_), .B(new_new_n815_), .C(new_new_n812_), .Y(new_new_n822_));
  NA2        g800(.A(new_new_n618_), .B(new_new_n117_), .Y(new_new_n823_));
  NO2        g801(.A(i_6_), .B(new_new_n823_), .Y(new_new_n824_));
  AOI210     g802(.A0(new_new_n433_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n825_));
  NA2        g803(.A(new_new_n167_), .B(new_new_n98_), .Y(new_new_n826_));
  NOi32      g804(.An(new_new_n825_), .Bn(new_new_n185_), .C(new_new_n826_), .Y(new_new_n827_));
  NO2        g805(.A(new_new_n827_), .B(new_new_n824_), .Y(new_new_n828_));
  OR2        g806(.A(new_new_n826_), .B(new_new_n502_), .Y(new_new_n829_));
  NO2        g807(.A(new_new_n252_), .B(new_new_n307_), .Y(new_new_n830_));
  INV        g808(.A(new_new_n665_), .Y(new_new_n831_));
  NA2        g809(.A(new_new_n831_), .B(new_new_n830_), .Y(new_new_n832_));
  NA4        g810(.A(new_new_n832_), .B(new_new_n829_), .C(new_new_n828_), .D(new_new_n822_), .Y(new_new_n833_));
  NO2        g811(.A(new_new_n788_), .B(new_new_n237_), .Y(new_new_n834_));
  AN2        g812(.A(new_new_n322_), .B(new_new_n317_), .Y(new_new_n835_));
  NA2        g813(.A(new_new_n834_), .B(i_10_), .Y(new_new_n836_));
  NA3        g814(.A(i_5_), .B(new_new_n399_), .C(new_new_n46_), .Y(new_new_n837_));
  OAI210     g815(.A0(new_new_n792_), .A1(i_7_), .B0(new_new_n837_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n816_), .B(new_new_n295_), .Y(new_new_n839_));
  NA2        g817(.A(new_new_n184_), .B(new_new_n839_), .Y(new_new_n840_));
  AOI220     g818(.A0(new_new_n840_), .A1(new_new_n461_), .B0(new_new_n838_), .B1(new_new_n67_), .Y(new_new_n841_));
  NO2        g819(.A(new_new_n69_), .B(new_new_n685_), .Y(new_new_n842_));
  AOI210     g820(.A0(new_new_n170_), .A1(new_new_n576_), .B0(new_new_n842_), .Y(new_new_n843_));
  NO2        g821(.A(new_new_n843_), .B(new_new_n48_), .Y(new_new_n844_));
  NO3        g822(.A(new_new_n570_), .B(new_new_n345_), .C(new_new_n24_), .Y(new_new_n845_));
  AOI210     g823(.A0(new_new_n647_), .A1(new_new_n531_), .B0(new_new_n845_), .Y(new_new_n846_));
  NAi21      g824(.An(i_9_), .B(i_5_), .Y(new_new_n847_));
  NO2        g825(.A(new_new_n847_), .B(new_new_n390_), .Y(new_new_n848_));
  NO2        g826(.A(new_new_n581_), .B(new_new_n100_), .Y(new_new_n849_));
  AOI220     g827(.A0(new_new_n849_), .A1(i_0_), .B0(new_new_n848_), .B1(new_new_n602_), .Y(new_new_n850_));
  OAI220     g828(.A0(new_new_n850_), .A1(new_new_n79_), .B0(new_new_n846_), .B1(new_new_n168_), .Y(new_new_n851_));
  NO2        g829(.A(new_new_n851_), .B(new_new_n844_), .Y(new_new_n852_));
  NA3        g830(.A(new_new_n852_), .B(new_new_n841_), .C(new_new_n836_), .Y(new_new_n853_));
  NO3        g831(.A(new_new_n853_), .B(new_new_n833_), .C(new_new_n809_), .Y(new_new_n854_));
  NO2        g832(.A(i_0_), .B(new_new_n665_), .Y(new_new_n855_));
  NA2        g833(.A(new_new_n67_), .B(new_new_n45_), .Y(new_new_n856_));
  NA2        g834(.A(new_new_n801_), .B(new_new_n856_), .Y(new_new_n857_));
  NO3        g835(.A(new_new_n100_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n858_));
  AO220      g836(.A0(new_new_n858_), .A1(new_new_n857_), .B0(new_new_n855_), .B1(new_new_n170_), .Y(new_new_n859_));
  NA2        g837(.A(new_new_n859_), .B(new_new_n335_), .Y(new_new_n860_));
  NA2        g838(.A(new_new_n967_), .B(new_new_n142_), .Y(new_new_n861_));
  INV        g839(.A(new_new_n861_), .Y(new_new_n862_));
  NA3        g840(.A(new_new_n862_), .B(new_new_n625_), .C(new_new_n67_), .Y(new_new_n863_));
  NO2        g841(.A(new_new_n740_), .B(new_new_n390_), .Y(new_new_n864_));
  NA3        g842(.A(new_new_n766_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n865_));
  NA2        g843(.A(new_new_n767_), .B(i_9_), .Y(new_new_n866_));
  AOI210     g844(.A0(new_new_n865_), .A1(new_new_n485_), .B0(new_new_n866_), .Y(new_new_n867_));
  OAI210     g845(.A0(new_new_n241_), .A1(i_9_), .B0(new_new_n228_), .Y(new_new_n868_));
  AOI210     g846(.A0(new_new_n868_), .A1(new_new_n795_), .B0(new_new_n150_), .Y(new_new_n869_));
  NO3        g847(.A(new_new_n869_), .B(new_new_n867_), .C(new_new_n864_), .Y(new_new_n870_));
  NA3        g848(.A(new_new_n870_), .B(new_new_n863_), .C(new_new_n860_), .Y(new_new_n871_));
  NA2        g849(.A(new_new_n835_), .B(new_new_n359_), .Y(new_new_n872_));
  AOI210     g850(.A0(new_new_n291_), .A1(new_new_n159_), .B0(new_new_n872_), .Y(new_new_n873_));
  NA3        g851(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n874_));
  NA2        g852(.A(new_new_n813_), .B(new_new_n473_), .Y(new_new_n875_));
  AOI210     g853(.A0(new_new_n874_), .A1(new_new_n159_), .B0(new_new_n875_), .Y(new_new_n876_));
  NO2        g854(.A(new_new_n876_), .B(new_new_n873_), .Y(new_new_n877_));
  NO3        g855(.A(new_new_n801_), .B(new_new_n782_), .C(new_new_n187_), .Y(new_new_n878_));
  AOI220     g856(.A0(new_new_n878_), .A1(i_11_), .B0(new_new_n550_), .B1(new_new_n69_), .Y(new_new_n879_));
  NO3        g857(.A(new_new_n209_), .B(new_new_n370_), .C(i_0_), .Y(new_new_n880_));
  OAI210     g858(.A0(new_new_n880_), .A1(new_new_n70_), .B0(i_13_), .Y(new_new_n881_));
  INV        g859(.A(new_new_n218_), .Y(new_new_n882_));
  NO2        g860(.A(i_12_), .B(new_new_n597_), .Y(new_new_n883_));
  NA3        g861(.A(new_new_n883_), .B(new_new_n968_), .C(new_new_n882_), .Y(new_new_n884_));
  NA4        g862(.A(new_new_n884_), .B(new_new_n881_), .C(new_new_n879_), .D(new_new_n877_), .Y(new_new_n885_));
  NO2        g863(.A(new_new_n240_), .B(new_new_n87_), .Y(new_new_n886_));
  AOI210     g864(.A0(new_new_n886_), .A1(new_new_n855_), .B0(new_new_n104_), .Y(new_new_n887_));
  AOI220     g865(.A0(i_7_), .A1(new_new_n473_), .B0(new_new_n766_), .B1(new_new_n160_), .Y(new_new_n888_));
  NA2        g866(.A(new_new_n338_), .B(new_new_n172_), .Y(new_new_n889_));
  OA220      g867(.A0(new_new_n889_), .A1(new_new_n888_), .B0(new_new_n887_), .B1(i_5_), .Y(new_new_n890_));
  AOI210     g868(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n171_), .Y(new_new_n891_));
  INV        g869(.A(new_new_n530_), .Y(new_new_n892_));
  NA2        g870(.A(new_new_n478_), .B(new_new_n459_), .Y(new_new_n893_));
  NO2        g871(.A(new_new_n893_), .B(new_new_n892_), .Y(new_new_n894_));
  NA3        g872(.A(new_new_n377_), .B(new_new_n167_), .C(new_new_n166_), .Y(new_new_n895_));
  NA3        g873(.A(new_new_n813_), .B(new_new_n281_), .C(new_new_n228_), .Y(new_new_n896_));
  NA2        g874(.A(new_new_n896_), .B(new_new_n895_), .Y(new_new_n897_));
  NOi31      g875(.An(new_new_n376_), .B(new_new_n856_), .C(new_new_n237_), .Y(new_new_n898_));
  NO2        g876(.A(new_new_n898_), .B(new_new_n897_), .Y(new_new_n899_));
  NA3        g877(.A(new_new_n899_), .B(new_new_n894_), .C(new_new_n890_), .Y(new_new_n900_));
  NO2        g878(.A(new_new_n79_), .B(i_5_), .Y(new_new_n901_));
  NA3        g879(.A(new_new_n767_), .B(new_new_n105_), .C(new_new_n120_), .Y(new_new_n902_));
  INV        g880(.A(new_new_n902_), .Y(new_new_n903_));
  NA2        g881(.A(new_new_n903_), .B(new_new_n901_), .Y(new_new_n904_));
  NA3        g882(.A(new_new_n295_), .B(i_5_), .C(new_new_n190_), .Y(new_new_n905_));
  INV        g883(.A(new_new_n240_), .Y(new_new_n906_));
  NO4        g884(.A(new_new_n237_), .B(new_new_n209_), .C(i_0_), .D(i_12_), .Y(new_new_n907_));
  AOI220     g885(.A0(new_new_n907_), .A1(new_new_n906_), .B0(new_new_n724_), .B1(new_new_n172_), .Y(new_new_n908_));
  AN2        g886(.A(new_new_n801_), .B(new_new_n150_), .Y(new_new_n909_));
  NO3        g887(.A(new_new_n909_), .B(i_12_), .C(new_new_n611_), .Y(new_new_n910_));
  NA2        g888(.A(new_new_n910_), .B(new_new_n218_), .Y(new_new_n911_));
  NA3        g889(.A(new_new_n93_), .B(new_new_n554_), .C(i_11_), .Y(new_new_n912_));
  NO2        g890(.A(new_new_n912_), .B(new_new_n152_), .Y(new_new_n913_));
  INV        g891(.A(new_new_n62_), .Y(new_new_n914_));
  NO2        g892(.A(new_new_n914_), .B(new_new_n905_), .Y(new_new_n915_));
  AOI210     g893(.A0(new_new_n915_), .A1(new_new_n817_), .B0(new_new_n913_), .Y(new_new_n916_));
  NA4        g894(.A(new_new_n916_), .B(new_new_n911_), .C(new_new_n908_), .D(new_new_n904_), .Y(new_new_n917_));
  NO4        g895(.A(new_new_n917_), .B(new_new_n900_), .C(new_new_n885_), .D(new_new_n871_), .Y(new_new_n918_));
  OAI210     g896(.A0(new_new_n743_), .A1(new_new_n738_), .B0(new_new_n37_), .Y(new_new_n919_));
  NA3        g897(.A(new_new_n825_), .B(new_new_n354_), .C(i_5_), .Y(new_new_n920_));
  NA3        g898(.A(new_new_n920_), .B(new_new_n919_), .C(new_new_n593_), .Y(new_new_n921_));
  NA2        g899(.A(new_new_n921_), .B(new_new_n205_), .Y(new_new_n922_));
  NA2        g900(.A(new_new_n183_), .B(new_new_n185_), .Y(new_new_n923_));
  AO210      g901(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n923_), .Y(new_new_n924_));
  OAI210     g902(.A0(new_new_n596_), .A1(new_new_n594_), .B0(new_new_n306_), .Y(new_new_n925_));
  NA2        g903(.A(new_new_n925_), .B(new_new_n924_), .Y(new_new_n926_));
  NO2        g904(.A(new_new_n449_), .B(new_new_n258_), .Y(new_new_n927_));
  NO4        g905(.A(new_new_n231_), .B(new_new_n141_), .C(new_new_n626_), .D(new_new_n37_), .Y(new_new_n928_));
  NO3        g906(.A(new_new_n928_), .B(new_new_n927_), .C(new_new_n797_), .Y(new_new_n929_));
  OAI210     g907(.A0(new_new_n912_), .A1(new_new_n144_), .B0(new_new_n929_), .Y(new_new_n930_));
  AOI210     g908(.A0(new_new_n926_), .A1(new_new_n49_), .B0(new_new_n930_), .Y(new_new_n931_));
  AOI210     g909(.A0(new_new_n931_), .A1(new_new_n922_), .B0(new_new_n67_), .Y(new_new_n932_));
  NO2        g910(.A(new_new_n547_), .B(new_new_n366_), .Y(new_new_n933_));
  NO2        g911(.A(new_new_n933_), .B(new_new_n691_), .Y(new_new_n934_));
  NA2        g912(.A(new_new_n966_), .B(new_new_n70_), .Y(new_new_n935_));
  NA2        g913(.A(new_new_n891_), .B(new_new_n813_), .Y(new_new_n936_));
  AOI210     g914(.A0(new_new_n936_), .A1(new_new_n935_), .B0(new_new_n626_), .Y(new_new_n937_));
  NA2        g915(.A(i_1_), .B(new_new_n70_), .Y(new_new_n938_));
  NO2        g916(.A(new_new_n938_), .B(new_new_n235_), .Y(new_new_n939_));
  NA3        g917(.A(new_new_n91_), .B(new_new_n297_), .C(new_new_n31_), .Y(new_new_n940_));
  INV        g918(.A(new_new_n940_), .Y(new_new_n941_));
  NO3        g919(.A(new_new_n941_), .B(new_new_n939_), .C(new_new_n937_), .Y(new_new_n942_));
  OAI210     g920(.A0(new_new_n260_), .A1(new_new_n155_), .B0(new_new_n82_), .Y(new_new_n943_));
  NA3        g921(.A(new_new_n694_), .B(new_new_n281_), .C(new_new_n74_), .Y(new_new_n944_));
  AOI210     g922(.A0(new_new_n944_), .A1(new_new_n943_), .B0(i_11_), .Y(new_new_n945_));
  NA2        g923(.A(new_new_n588_), .B(new_new_n215_), .Y(new_new_n946_));
  OAI210     g924(.A0(new_new_n946_), .A1(new_new_n825_), .B0(new_new_n205_), .Y(new_new_n947_));
  NA2        g925(.A(new_new_n161_), .B(i_5_), .Y(new_new_n948_));
  NO2        g926(.A(new_new_n947_), .B(new_new_n948_), .Y(new_new_n949_));
  NO3        g927(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n950_));
  NA2        g928(.A(new_new_n297_), .B(new_new_n950_), .Y(new_new_n951_));
  NO2        g929(.A(new_new_n951_), .B(new_new_n665_), .Y(new_new_n952_));
  NO3        g930(.A(new_new_n847_), .B(new_new_n464_), .C(new_new_n250_), .Y(new_new_n953_));
  NO2        g931(.A(new_new_n953_), .B(new_new_n544_), .Y(new_new_n954_));
  INV        g932(.A(new_new_n348_), .Y(new_new_n955_));
  AOI210     g933(.A0(new_new_n955_), .A1(new_new_n954_), .B0(new_new_n41_), .Y(new_new_n956_));
  NO4        g934(.A(new_new_n956_), .B(new_new_n952_), .C(new_new_n949_), .D(new_new_n945_), .Y(new_new_n957_));
  OAI210     g935(.A0(new_new_n942_), .A1(i_4_), .B0(new_new_n957_), .Y(new_new_n958_));
  NO3        g936(.A(new_new_n958_), .B(new_new_n934_), .C(new_new_n932_), .Y(new_new_n959_));
  NA4        g937(.A(new_new_n959_), .B(new_new_n918_), .C(new_new_n854_), .D(new_new_n787_), .Y(men4));
  INV        g938(.A(new_new_n646_), .Y(new_new_n963_));
  INV        g939(.A(i_2_), .Y(new_new_n964_));
  INV        g940(.A(new_new_n774_), .Y(new_new_n965_));
  INV        g941(.A(i_7_), .Y(new_new_n966_));
  INV        g942(.A(i_2_), .Y(new_new_n967_));
  INV        g943(.A(i_3_), .Y(new_new_n968_));
  INV        g944(.A(i_8_), .Y(new_new_n969_));
  INV        g945(.A(new_new_n140_), .Y(new_new_n970_));
  INV        g946(.A(new_new_n195_), .Y(new_new_n971_));
  INV        g947(.A(new_new_n588_), .Y(new_new_n972_));
  INV        g948(.A(i_12_), .Y(new_new_n973_));
  INV        g949(.A(i_10_), .Y(new_new_n974_));
  INV        g950(.A(i_1_), .Y(new_new_n975_));
  INV        g951(.A(new_new_n693_), .Y(new_new_n976_));
  INV        g952(.A(i_12_), .Y(new_new_n977_));
endmodule


