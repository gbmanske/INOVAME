//Benchmark atmr_max1024_476_0.125

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n426_, men_men_n427_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  INV        o005(.A(ori_ori_n19_), .Y(ori_ori_n22_));
  NA2        o006(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n23_));
  INV        o007(.A(x5), .Y(ori_ori_n24_));
  NA2        o008(.A(x7), .B(x6), .Y(ori_ori_n25_));
  NA2        o009(.A(x8), .B(x3), .Y(ori_ori_n26_));
  NA2        o010(.A(x4), .B(x2), .Y(ori_ori_n27_));
  NO4        o011(.A(ori_ori_n27_), .B(ori_ori_n26_), .C(ori_ori_n25_), .D(ori_ori_n24_), .Y(ori_ori_n28_));
  NO2        o012(.A(ori_ori_n28_), .B(ori_ori_n23_), .Y(ori_ori_n29_));
  NO2        o013(.A(x4), .B(x3), .Y(ori_ori_n30_));
  INV        o014(.A(ori_ori_n30_), .Y(ori_ori_n31_));
  NOi21      o015(.An(ori_ori_n22_), .B(ori_ori_n29_), .Y(ori00));
  NO2        o016(.A(x1), .B(x0), .Y(ori_ori_n33_));
  INV        o017(.A(x6), .Y(ori_ori_n34_));
  NO2        o018(.A(ori_ori_n34_), .B(ori_ori_n24_), .Y(ori_ori_n35_));
  AN2        o019(.A(x8), .B(x7), .Y(ori_ori_n36_));
  NA3        o020(.A(ori_ori_n36_), .B(ori_ori_n35_), .C(ori_ori_n33_), .Y(ori_ori_n37_));
  NA2        o021(.A(x4), .B(x3), .Y(ori_ori_n38_));
  AOI210     o022(.A0(ori_ori_n37_), .A1(ori_ori_n22_), .B0(ori_ori_n38_), .Y(ori_ori_n39_));
  NO2        o023(.A(x2), .B(x0), .Y(ori_ori_n40_));
  INV        o024(.A(x3), .Y(ori_ori_n41_));
  NO2        o025(.A(ori_ori_n41_), .B(ori_ori_n18_), .Y(ori_ori_n42_));
  INV        o026(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n35_), .B(x4), .Y(ori_ori_n44_));
  OAI210     o028(.A0(ori_ori_n44_), .A1(ori_ori_n43_), .B0(ori_ori_n40_), .Y(ori_ori_n45_));
  INV        o029(.A(x4), .Y(ori_ori_n46_));
  NO2        o030(.A(ori_ori_n46_), .B(ori_ori_n17_), .Y(ori_ori_n47_));
  NA2        o031(.A(ori_ori_n47_), .B(x2), .Y(ori_ori_n48_));
  OAI210     o032(.A0(ori_ori_n48_), .A1(ori_ori_n20_), .B0(ori_ori_n45_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n50_));
  NA2        o034(.A(ori_ori_n50_), .B(ori_ori_n33_), .Y(ori_ori_n51_));
  INV        o035(.A(x2), .Y(ori_ori_n52_));
  NO2        o036(.A(ori_ori_n52_), .B(ori_ori_n17_), .Y(ori_ori_n53_));
  NA2        o037(.A(ori_ori_n41_), .B(ori_ori_n18_), .Y(ori_ori_n54_));
  NA2        o038(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  OAI210     o039(.A0(ori_ori_n51_), .A1(ori_ori_n31_), .B0(ori_ori_n55_), .Y(ori_ori_n56_));
  NO3        o040(.A(ori_ori_n56_), .B(ori_ori_n49_), .C(ori_ori_n39_), .Y(ori01));
  NA2        o041(.A(x8), .B(x7), .Y(ori_ori_n58_));
  NA2        o042(.A(ori_ori_n41_), .B(x1), .Y(ori_ori_n59_));
  INV        o043(.A(x9), .Y(ori_ori_n60_));
  NO2        o044(.A(x7), .B(x6), .Y(ori_ori_n61_));
  NO2        o045(.A(ori_ori_n59_), .B(x5), .Y(ori_ori_n62_));
  NO2        o046(.A(x8), .B(x2), .Y(ori_ori_n63_));
  AN2        o047(.A(ori_ori_n63_), .B(ori_ori_n61_), .Y(ori_ori_n64_));
  OAI210     o048(.A0(ori_ori_n42_), .A1(ori_ori_n24_), .B0(ori_ori_n52_), .Y(ori_ori_n65_));
  OAI210     o049(.A0(ori_ori_n54_), .A1(ori_ori_n20_), .B0(ori_ori_n65_), .Y(ori_ori_n66_));
  NO2        o050(.A(ori_ori_n66_), .B(ori_ori_n64_), .Y(ori_ori_n67_));
  NA2        o051(.A(ori_ori_n67_), .B(x4), .Y(ori_ori_n68_));
  NA2        o052(.A(ori_ori_n46_), .B(x2), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n69_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n70_));
  NA2        o054(.A(x5), .B(x3), .Y(ori_ori_n71_));
  NO2        o055(.A(x8), .B(x6), .Y(ori_ori_n72_));
  NO4        o056(.A(ori_ori_n72_), .B(ori_ori_n71_), .C(ori_ori_n61_), .D(ori_ori_n52_), .Y(ori_ori_n73_));
  NAi21      o057(.An(x4), .B(x3), .Y(ori_ori_n74_));
  INV        o058(.A(ori_ori_n74_), .Y(ori_ori_n75_));
  NO2        o059(.A(x4), .B(x2), .Y(ori_ori_n76_));
  NO2        o060(.A(ori_ori_n74_), .B(ori_ori_n18_), .Y(ori_ori_n77_));
  NO3        o061(.A(ori_ori_n77_), .B(ori_ori_n73_), .C(ori_ori_n70_), .Y(ori_ori_n78_));
  NA2        o062(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n79_));
  NO2        o063(.A(ori_ori_n79_), .B(ori_ori_n24_), .Y(ori_ori_n80_));
  INV        o064(.A(x8), .Y(ori_ori_n81_));
  NA2        o065(.A(x2), .B(x1), .Y(ori_ori_n82_));
  INV        o066(.A(ori_ori_n80_), .Y(ori_ori_n83_));
  NO2        o067(.A(ori_ori_n83_), .B(ori_ori_n25_), .Y(ori_ori_n84_));
  AOI210     o068(.A0(ori_ori_n54_), .A1(ori_ori_n24_), .B0(ori_ori_n52_), .Y(ori_ori_n85_));
  OAI210     o069(.A0(ori_ori_n43_), .A1(ori_ori_n35_), .B0(ori_ori_n46_), .Y(ori_ori_n86_));
  NO3        o070(.A(ori_ori_n86_), .B(ori_ori_n85_), .C(ori_ori_n84_), .Y(ori_ori_n87_));
  NA2        o071(.A(x4), .B(ori_ori_n41_), .Y(ori_ori_n88_));
  NO2        o072(.A(ori_ori_n46_), .B(ori_ori_n52_), .Y(ori_ori_n89_));
  OAI210     o073(.A0(ori_ori_n89_), .A1(ori_ori_n41_), .B0(ori_ori_n18_), .Y(ori_ori_n90_));
  AOI210     o074(.A0(ori_ori_n88_), .A1(ori_ori_n50_), .B0(ori_ori_n90_), .Y(ori_ori_n91_));
  NA2        o075(.A(ori_ori_n52_), .B(x1), .Y(ori_ori_n92_));
  OAI210     o076(.A0(ori_ori_n92_), .A1(ori_ori_n38_), .B0(ori_ori_n17_), .Y(ori_ori_n93_));
  NO3        o077(.A(ori_ori_n93_), .B(ori_ori_n91_), .C(ori_ori_n87_), .Y(ori_ori_n94_));
  AO210      o078(.A0(ori_ori_n78_), .A1(ori_ori_n68_), .B0(ori_ori_n94_), .Y(ori02));
  NO2        o079(.A(x3), .B(ori_ori_n52_), .Y(ori_ori_n96_));
  NA2        o080(.A(ori_ori_n41_), .B(x0), .Y(ori_ori_n97_));
  OR2        o081(.A(x8), .B(x0), .Y(ori_ori_n98_));
  INV        o082(.A(ori_ori_n98_), .Y(ori_ori_n99_));
  NO2        o083(.A(x4), .B(x1), .Y(ori_ori_n100_));
  NA3        o084(.A(ori_ori_n100_), .B(x2), .C(ori_ori_n58_), .Y(ori_ori_n101_));
  NOi21      o085(.An(x0), .B(x1), .Y(ori_ori_n102_));
  NO3        o086(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n103_));
  NOi21      o087(.An(x0), .B(x4), .Y(ori_ori_n104_));
  NAi21      o088(.An(x8), .B(x7), .Y(ori_ori_n105_));
  NO2        o089(.A(ori_ori_n105_), .B(ori_ori_n60_), .Y(ori_ori_n106_));
  AOI220     o090(.A0(ori_ori_n106_), .A1(ori_ori_n104_), .B0(ori_ori_n103_), .B1(ori_ori_n102_), .Y(ori_ori_n107_));
  AOI210     o091(.A0(ori_ori_n107_), .A1(ori_ori_n101_), .B0(ori_ori_n71_), .Y(ori_ori_n108_));
  NO2        o092(.A(x5), .B(ori_ori_n46_), .Y(ori_ori_n109_));
  NA2        o093(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n110_));
  AOI210     o094(.A0(ori_ori_n110_), .A1(ori_ori_n92_), .B0(ori_ori_n97_), .Y(ori_ori_n111_));
  OAI210     o095(.A0(ori_ori_n111_), .A1(ori_ori_n33_), .B0(ori_ori_n109_), .Y(ori_ori_n112_));
  NAi21      o096(.An(x0), .B(x4), .Y(ori_ori_n113_));
  NO2        o097(.A(ori_ori_n113_), .B(x1), .Y(ori_ori_n114_));
  NO2        o098(.A(x7), .B(x0), .Y(ori_ori_n115_));
  NO2        o099(.A(ori_ori_n76_), .B(ori_ori_n89_), .Y(ori_ori_n116_));
  NO2        o100(.A(ori_ori_n116_), .B(x3), .Y(ori_ori_n117_));
  OAI210     o101(.A0(ori_ori_n115_), .A1(ori_ori_n114_), .B0(ori_ori_n117_), .Y(ori_ori_n118_));
  NA2        o102(.A(x5), .B(x0), .Y(ori_ori_n119_));
  NO2        o103(.A(ori_ori_n46_), .B(x2), .Y(ori_ori_n120_));
  NA3        o104(.A(ori_ori_n118_), .B(ori_ori_n112_), .C(ori_ori_n34_), .Y(ori_ori_n121_));
  NO2        o105(.A(ori_ori_n121_), .B(ori_ori_n108_), .Y(ori_ori_n122_));
  NO3        o106(.A(ori_ori_n71_), .B(ori_ori_n69_), .C(ori_ori_n23_), .Y(ori_ori_n123_));
  NO2        o107(.A(ori_ori_n27_), .B(ori_ori_n24_), .Y(ori_ori_n124_));
  NA2        o108(.A(x7), .B(x3), .Y(ori_ori_n125_));
  NO2        o109(.A(ori_ori_n88_), .B(x5), .Y(ori_ori_n126_));
  NO2        o110(.A(x9), .B(x7), .Y(ori_ori_n127_));
  NOi21      o111(.An(x8), .B(x0), .Y(ori_ori_n128_));
  NO2        o112(.A(ori_ori_n41_), .B(x2), .Y(ori_ori_n129_));
  INV        o113(.A(x7), .Y(ori_ori_n130_));
  NA2        o114(.A(ori_ori_n130_), .B(ori_ori_n18_), .Y(ori_ori_n131_));
  AOI220     o115(.A0(ori_ori_n131_), .A1(ori_ori_n129_), .B0(ori_ori_n96_), .B1(ori_ori_n36_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n24_), .B(x4), .Y(ori_ori_n133_));
  NO2        o117(.A(ori_ori_n133_), .B(ori_ori_n104_), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n134_), .B(ori_ori_n132_), .Y(ori_ori_n135_));
  AOI210     o119(.A0(ori_ori_n127_), .A1(ori_ori_n126_), .B0(ori_ori_n135_), .Y(ori_ori_n136_));
  OAI210     o120(.A0(ori_ori_n125_), .A1(ori_ori_n48_), .B0(ori_ori_n136_), .Y(ori_ori_n137_));
  NA2        o121(.A(x5), .B(x1), .Y(ori_ori_n138_));
  INV        o122(.A(ori_ori_n138_), .Y(ori_ori_n139_));
  AOI210     o123(.A0(ori_ori_n139_), .A1(ori_ori_n104_), .B0(ori_ori_n34_), .Y(ori_ori_n140_));
  NAi21      o124(.An(x2), .B(x7), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n141_), .B(ori_ori_n46_), .Y(ori_ori_n142_));
  NA2        o126(.A(ori_ori_n142_), .B(ori_ori_n62_), .Y(ori_ori_n143_));
  NAi31      o127(.An(ori_ori_n71_), .B(ori_ori_n36_), .C(ori_ori_n33_), .Y(ori_ori_n144_));
  NA3        o128(.A(ori_ori_n144_), .B(ori_ori_n143_), .C(ori_ori_n140_), .Y(ori_ori_n145_));
  NO3        o129(.A(ori_ori_n145_), .B(ori_ori_n137_), .C(ori_ori_n123_), .Y(ori_ori_n146_));
  NO2        o130(.A(ori_ori_n146_), .B(ori_ori_n122_), .Y(ori_ori_n147_));
  NO2        o131(.A(ori_ori_n119_), .B(ori_ori_n116_), .Y(ori_ori_n148_));
  NA2        o132(.A(ori_ori_n24_), .B(ori_ori_n18_), .Y(ori_ori_n149_));
  NA2        o133(.A(ori_ori_n24_), .B(ori_ori_n17_), .Y(ori_ori_n150_));
  NA3        o134(.A(ori_ori_n150_), .B(ori_ori_n149_), .C(ori_ori_n23_), .Y(ori_ori_n151_));
  AN2        o135(.A(ori_ori_n151_), .B(ori_ori_n120_), .Y(ori_ori_n152_));
  NA2        o136(.A(x8), .B(x0), .Y(ori_ori_n153_));
  NO2        o137(.A(ori_ori_n130_), .B(ori_ori_n24_), .Y(ori_ori_n154_));
  NA2        o138(.A(x2), .B(x0), .Y(ori_ori_n155_));
  NA2        o139(.A(x4), .B(x1), .Y(ori_ori_n156_));
  NAi21      o140(.An(ori_ori_n100_), .B(ori_ori_n156_), .Y(ori_ori_n157_));
  NOi31      o141(.An(ori_ori_n157_), .B(ori_ori_n133_), .C(ori_ori_n155_), .Y(ori_ori_n158_));
  NO3        o142(.A(ori_ori_n158_), .B(ori_ori_n152_), .C(ori_ori_n148_), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n159_), .B(ori_ori_n41_), .Y(ori_ori_n160_));
  NO2        o144(.A(ori_ori_n151_), .B(ori_ori_n69_), .Y(ori_ori_n161_));
  INV        o145(.A(ori_ori_n109_), .Y(ori_ori_n162_));
  NO2        o146(.A(ori_ori_n92_), .B(ori_ori_n17_), .Y(ori_ori_n163_));
  NA2        o147(.A(ori_ori_n157_), .B(ori_ori_n40_), .Y(ori_ori_n164_));
  OAI210     o148(.A0(ori_ori_n150_), .A1(ori_ori_n116_), .B0(ori_ori_n164_), .Y(ori_ori_n165_));
  NO2        o149(.A(ori_ori_n165_), .B(ori_ori_n161_), .Y(ori_ori_n166_));
  NO2        o150(.A(ori_ori_n166_), .B(x3), .Y(ori_ori_n167_));
  NO3        o151(.A(ori_ori_n167_), .B(ori_ori_n160_), .C(ori_ori_n147_), .Y(ori03));
  NO2        o152(.A(ori_ori_n46_), .B(x3), .Y(ori_ori_n169_));
  NO2        o153(.A(x6), .B(ori_ori_n24_), .Y(ori_ori_n170_));
  NO2        o154(.A(ori_ori_n52_), .B(x1), .Y(ori_ori_n171_));
  NA2        o155(.A(x6), .B(ori_ori_n24_), .Y(ori_ori_n172_));
  NO2        o156(.A(ori_ori_n172_), .B(x4), .Y(ori_ori_n173_));
  NO2        o157(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n174_));
  NA2        o158(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n175_));
  NO2        o159(.A(ori_ori_n175_), .B(ori_ori_n172_), .Y(ori_ori_n176_));
  NA2        o160(.A(x9), .B(ori_ori_n52_), .Y(ori_ori_n177_));
  NA2        o161(.A(ori_ori_n172_), .B(ori_ori_n74_), .Y(ori_ori_n178_));
  AOI210     o162(.A0(ori_ori_n24_), .A1(x3), .B0(ori_ori_n155_), .Y(ori_ori_n179_));
  AOI210     o163(.A0(ori_ori_n179_), .A1(ori_ori_n178_), .B0(ori_ori_n176_), .Y(ori_ori_n180_));
  NO3        o164(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n181_));
  NO2        o165(.A(x5), .B(x1), .Y(ori_ori_n182_));
  NO2        o166(.A(ori_ori_n175_), .B(ori_ori_n149_), .Y(ori_ori_n183_));
  NO3        o167(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n184_));
  AOI220     o168(.A0(ori_ori_n184_), .A1(ori_ori_n46_), .B0(ori_ori_n181_), .B1(ori_ori_n109_), .Y(ori_ori_n185_));
  NA2        o169(.A(ori_ori_n185_), .B(ori_ori_n180_), .Y(ori_ori_n186_));
  NO2        o170(.A(ori_ori_n46_), .B(ori_ori_n41_), .Y(ori_ori_n187_));
  NA2        o171(.A(ori_ori_n187_), .B(ori_ori_n19_), .Y(ori_ori_n188_));
  NO2        o172(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n189_));
  NO2        o173(.A(ori_ori_n189_), .B(x6), .Y(ori_ori_n190_));
  NOi21      o174(.An(ori_ori_n76_), .B(ori_ori_n190_), .Y(ori_ori_n191_));
  NA2        o175(.A(ori_ori_n60_), .B(ori_ori_n81_), .Y(ori_ori_n192_));
  NA3        o176(.A(ori_ori_n192_), .B(ori_ori_n189_), .C(x6), .Y(ori_ori_n193_));
  AOI210     o177(.A0(ori_ori_n193_), .A1(ori_ori_n191_), .B0(ori_ori_n130_), .Y(ori_ori_n194_));
  OR2        o178(.A(ori_ori_n194_), .B(ori_ori_n154_), .Y(ori_ori_n195_));
  NA2        o179(.A(ori_ori_n41_), .B(ori_ori_n52_), .Y(ori_ori_n196_));
  OAI210     o180(.A0(ori_ori_n196_), .A1(ori_ori_n24_), .B0(ori_ori_n150_), .Y(ori_ori_n197_));
  NO3        o181(.A(ori_ori_n156_), .B(ori_ori_n60_), .C(x6), .Y(ori_ori_n198_));
  AOI220     o182(.A0(ori_ori_n198_), .A1(ori_ori_n197_), .B0(ori_ori_n120_), .B1(ori_ori_n80_), .Y(ori_ori_n199_));
  NA2        o183(.A(x6), .B(ori_ori_n46_), .Y(ori_ori_n200_));
  OAI210     o184(.A0(ori_ori_n99_), .A1(ori_ori_n72_), .B0(x4), .Y(ori_ori_n201_));
  AOI210     o185(.A0(ori_ori_n201_), .A1(ori_ori_n200_), .B0(ori_ori_n71_), .Y(ori_ori_n202_));
  NO2        o186(.A(ori_ori_n60_), .B(x6), .Y(ori_ori_n203_));
  NO2        o187(.A(ori_ori_n138_), .B(ori_ori_n41_), .Y(ori_ori_n204_));
  OAI210     o188(.A0(ori_ori_n204_), .A1(ori_ori_n183_), .B0(ori_ori_n203_), .Y(ori_ori_n205_));
  NA2        o189(.A(ori_ori_n170_), .B(ori_ori_n114_), .Y(ori_ori_n206_));
  NA3        o190(.A(ori_ori_n175_), .B(ori_ori_n109_), .C(x6), .Y(ori_ori_n207_));
  INV        o191(.A(ori_ori_n62_), .Y(ori_ori_n208_));
  NA4        o192(.A(ori_ori_n208_), .B(ori_ori_n207_), .C(ori_ori_n206_), .D(ori_ori_n205_), .Y(ori_ori_n209_));
  OAI210     o193(.A0(ori_ori_n209_), .A1(ori_ori_n202_), .B0(x2), .Y(ori_ori_n210_));
  NA3        o194(.A(ori_ori_n210_), .B(ori_ori_n199_), .C(ori_ori_n195_), .Y(ori_ori_n211_));
  AOI210     o195(.A0(ori_ori_n186_), .A1(x8), .B0(ori_ori_n211_), .Y(ori_ori_n212_));
  NO2        o196(.A(ori_ori_n81_), .B(x3), .Y(ori_ori_n213_));
  NA2        o197(.A(ori_ori_n213_), .B(ori_ori_n173_), .Y(ori_ori_n214_));
  NO3        o198(.A(ori_ori_n79_), .B(ori_ori_n72_), .C(ori_ori_n24_), .Y(ori_ori_n215_));
  AOI210     o199(.A0(ori_ori_n190_), .A1(ori_ori_n133_), .B0(ori_ori_n215_), .Y(ori_ori_n216_));
  AOI210     o200(.A0(ori_ori_n216_), .A1(ori_ori_n214_), .B0(x2), .Y(ori_ori_n217_));
  NO2        o201(.A(x4), .B(ori_ori_n52_), .Y(ori_ori_n218_));
  AOI220     o202(.A0(ori_ori_n173_), .A1(ori_ori_n163_), .B0(ori_ori_n218_), .B1(ori_ori_n62_), .Y(ori_ori_n219_));
  NA2        o203(.A(ori_ori_n60_), .B(x6), .Y(ori_ori_n220_));
  NA3        o204(.A(ori_ori_n24_), .B(x3), .C(x2), .Y(ori_ori_n221_));
  AOI210     o205(.A0(ori_ori_n221_), .A1(ori_ori_n119_), .B0(ori_ori_n220_), .Y(ori_ori_n222_));
  NA2        o206(.A(ori_ori_n41_), .B(ori_ori_n17_), .Y(ori_ori_n223_));
  NO2        o207(.A(ori_ori_n223_), .B(ori_ori_n24_), .Y(ori_ori_n224_));
  OAI210     o208(.A0(ori_ori_n224_), .A1(ori_ori_n222_), .B0(ori_ori_n100_), .Y(ori_ori_n225_));
  NA2        o209(.A(ori_ori_n175_), .B(x6), .Y(ori_ori_n226_));
  NO2        o210(.A(ori_ori_n175_), .B(x6), .Y(ori_ori_n227_));
  INV        o211(.A(ori_ori_n227_), .Y(ori_ori_n228_));
  NA3        o212(.A(ori_ori_n228_), .B(ori_ori_n226_), .C(ori_ori_n124_), .Y(ori_ori_n229_));
  NA4        o213(.A(ori_ori_n229_), .B(ori_ori_n225_), .C(ori_ori_n219_), .D(ori_ori_n130_), .Y(ori_ori_n230_));
  NA2        o214(.A(ori_ori_n170_), .B(ori_ori_n189_), .Y(ori_ori_n231_));
  NO2        o215(.A(x9), .B(x6), .Y(ori_ori_n232_));
  NO2        o216(.A(ori_ori_n119_), .B(ori_ori_n18_), .Y(ori_ori_n233_));
  NAi21      o217(.An(ori_ori_n233_), .B(ori_ori_n221_), .Y(ori_ori_n234_));
  AOI220     o218(.A0(x2), .A1(x1), .B0(ori_ori_n234_), .B1(ori_ori_n232_), .Y(ori_ori_n235_));
  NA2        o219(.A(ori_ori_n235_), .B(ori_ori_n231_), .Y(ori_ori_n236_));
  NA2        o220(.A(ori_ori_n60_), .B(x2), .Y(ori_ori_n237_));
  NO2        o221(.A(ori_ori_n237_), .B(ori_ori_n231_), .Y(ori_ori_n238_));
  NA2        o222(.A(x6), .B(x2), .Y(ori_ori_n239_));
  OAI210     o223(.A0(x4), .A1(ori_ori_n238_), .B0(ori_ori_n236_), .Y(ori_ori_n240_));
  NA2        o224(.A(x4), .B(x0), .Y(ori_ori_n241_));
  NO2        o225(.A(ori_ori_n240_), .B(x8), .Y(ori_ori_n242_));
  INV        o226(.A(ori_ori_n220_), .Y(ori_ori_n243_));
  OAI210     o227(.A0(ori_ori_n233_), .A1(ori_ori_n182_), .B0(ori_ori_n243_), .Y(ori_ori_n244_));
  OAI210     o228(.A0(x0), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n245_));
  AOI210     o229(.A0(ori_ori_n245_), .A1(ori_ori_n244_), .B0(ori_ori_n196_), .Y(ori_ori_n246_));
  NO4        o230(.A(ori_ori_n246_), .B(ori_ori_n242_), .C(ori_ori_n230_), .D(ori_ori_n217_), .Y(ori_ori_n247_));
  INV        o231(.A(x1), .Y(ori_ori_n248_));
  OAI210     o232(.A0(x1), .A1(ori_ori_n227_), .B0(x2), .Y(ori_ori_n249_));
  OAI210     o233(.A0(x0), .A1(x6), .B0(ori_ori_n42_), .Y(ori_ori_n250_));
  AOI210     o234(.A0(ori_ori_n250_), .A1(ori_ori_n249_), .B0(ori_ori_n162_), .Y(ori_ori_n251_));
  NOi21      o235(.An(ori_ori_n239_), .B(ori_ori_n17_), .Y(ori_ori_n252_));
  NA3        o236(.A(ori_ori_n252_), .B(ori_ori_n182_), .C(ori_ori_n38_), .Y(ori_ori_n253_));
  AOI210     o237(.A0(ori_ori_n34_), .A1(ori_ori_n52_), .B0(x0), .Y(ori_ori_n254_));
  NA3        o238(.A(ori_ori_n254_), .B(ori_ori_n139_), .C(ori_ori_n31_), .Y(ori_ori_n255_));
  NA2        o239(.A(x3), .B(x2), .Y(ori_ori_n256_));
  AOI220     o240(.A0(ori_ori_n256_), .A1(ori_ori_n196_), .B0(ori_ori_n255_), .B1(ori_ori_n253_), .Y(ori_ori_n257_));
  NAi21      o241(.An(x4), .B(x0), .Y(ori_ori_n258_));
  NO3        o242(.A(ori_ori_n258_), .B(ori_ori_n42_), .C(x2), .Y(ori_ori_n259_));
  OAI210     o243(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n259_), .Y(ori_ori_n260_));
  OAI220     o244(.A0(ori_ori_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n261_));
  NO2        o245(.A(ori_ori_n254_), .B(ori_ori_n252_), .Y(ori_ori_n262_));
  AOI220     o246(.A0(ori_ori_n262_), .A1(ori_ori_n75_), .B0(ori_ori_n261_), .B1(ori_ori_n30_), .Y(ori_ori_n263_));
  AOI210     o247(.A0(ori_ori_n263_), .A1(ori_ori_n260_), .B0(ori_ori_n24_), .Y(ori_ori_n264_));
  NA3        o248(.A(ori_ori_n34_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n265_));
  NO2        o249(.A(ori_ori_n254_), .B(ori_ori_n252_), .Y(ori_ori_n266_));
  INV        o250(.A(ori_ori_n183_), .Y(ori_ori_n267_));
  NA2        o251(.A(ori_ori_n34_), .B(ori_ori_n41_), .Y(ori_ori_n268_));
  OR2        o252(.A(ori_ori_n268_), .B(ori_ori_n241_), .Y(ori_ori_n269_));
  OAI220     o253(.A0(ori_ori_n269_), .A1(ori_ori_n138_), .B0(ori_ori_n200_), .B1(ori_ori_n267_), .Y(ori_ori_n270_));
  AO210      o254(.A0(ori_ori_n266_), .A1(ori_ori_n126_), .B0(ori_ori_n270_), .Y(ori_ori_n271_));
  NO4        o255(.A(ori_ori_n271_), .B(ori_ori_n264_), .C(ori_ori_n257_), .D(ori_ori_n251_), .Y(ori_ori_n272_));
  OAI210     o256(.A0(ori_ori_n247_), .A1(ori_ori_n212_), .B0(ori_ori_n272_), .Y(ori04));
  NO2        o257(.A(x2), .B(x1), .Y(ori_ori_n274_));
  OAI210     o258(.A0(ori_ori_n223_), .A1(ori_ori_n274_), .B0(ori_ori_n34_), .Y(ori_ori_n275_));
  NO2        o259(.A(ori_ori_n274_), .B(ori_ori_n258_), .Y(ori_ori_n276_));
  OAI210     o260(.A0(ori_ori_n52_), .A1(ori_ori_n276_), .B0(ori_ori_n213_), .Y(ori_ori_n277_));
  NO2        o261(.A(ori_ori_n237_), .B(ori_ori_n79_), .Y(ori_ori_n278_));
  NO2        o262(.A(ori_ori_n278_), .B(ori_ori_n34_), .Y(ori_ori_n279_));
  NO2        o263(.A(ori_ori_n256_), .B(ori_ori_n174_), .Y(ori_ori_n280_));
  NA2        o264(.A(x9), .B(x0), .Y(ori_ori_n281_));
  AOI210     o265(.A0(ori_ori_n79_), .A1(ori_ori_n69_), .B0(ori_ori_n281_), .Y(ori_ori_n282_));
  OAI210     o266(.A0(ori_ori_n282_), .A1(ori_ori_n280_), .B0(ori_ori_n81_), .Y(ori_ori_n283_));
  NA3        o267(.A(ori_ori_n283_), .B(ori_ori_n279_), .C(ori_ori_n277_), .Y(ori_ori_n284_));
  NA2        o268(.A(ori_ori_n284_), .B(ori_ori_n275_), .Y(ori_ori_n285_));
  NO2        o269(.A(ori_ori_n177_), .B(ori_ori_n97_), .Y(ori_ori_n286_));
  NO3        o270(.A(ori_ori_n220_), .B(x2), .C(ori_ori_n18_), .Y(ori_ori_n287_));
  NO2        o271(.A(ori_ori_n287_), .B(ori_ori_n286_), .Y(ori_ori_n288_));
  OAI210     o272(.A0(ori_ori_n98_), .A1(ori_ori_n92_), .B0(ori_ori_n153_), .Y(ori_ori_n289_));
  NA3        o273(.A(ori_ori_n289_), .B(x6), .C(x3), .Y(ori_ori_n290_));
  NO2        o274(.A(ori_ori_n237_), .B(ori_ori_n265_), .Y(ori_ori_n291_));
  INV        o275(.A(ori_ori_n291_), .Y(ori_ori_n292_));
  NA2        o276(.A(ori_ori_n278_), .B(ori_ori_n81_), .Y(ori_ori_n293_));
  NA4        o277(.A(ori_ori_n293_), .B(ori_ori_n292_), .C(ori_ori_n290_), .D(ori_ori_n288_), .Y(ori_ori_n294_));
  NA2        o278(.A(ori_ori_n181_), .B(ori_ori_n76_), .Y(ori_ori_n295_));
  NA2        o279(.A(ori_ori_n295_), .B(ori_ori_n130_), .Y(ori_ori_n296_));
  AOI210     o280(.A0(ori_ori_n294_), .A1(x4), .B0(ori_ori_n296_), .Y(ori_ori_n297_));
  NA3        o281(.A(ori_ori_n276_), .B(ori_ori_n177_), .C(ori_ori_n81_), .Y(ori_ori_n298_));
  XO2        o282(.A(x4), .B(x0), .Y(ori_ori_n299_));
  NA2        o283(.A(x4), .B(ori_ori_n82_), .Y(ori_ori_n300_));
  AOI210     o284(.A0(ori_ori_n300_), .A1(ori_ori_n298_), .B0(x3), .Y(ori_ori_n301_));
  INV        o285(.A(ori_ori_n82_), .Y(ori_ori_n302_));
  NO2        o286(.A(ori_ori_n81_), .B(x4), .Y(ori_ori_n303_));
  AOI220     o287(.A0(ori_ori_n303_), .A1(ori_ori_n42_), .B0(ori_ori_n104_), .B1(ori_ori_n302_), .Y(ori_ori_n304_));
  NO2        o288(.A(ori_ori_n299_), .B(x2), .Y(ori_ori_n305_));
  NO3        o289(.A(ori_ori_n192_), .B(ori_ori_n27_), .C(ori_ori_n23_), .Y(ori_ori_n306_));
  NO2        o290(.A(ori_ori_n306_), .B(ori_ori_n305_), .Y(ori_ori_n307_));
  NA4        o291(.A(ori_ori_n307_), .B(ori_ori_n304_), .C(ori_ori_n188_), .D(x6), .Y(ori_ori_n308_));
  OAI220     o292(.A0(ori_ori_n258_), .A1(ori_ori_n79_), .B0(ori_ori_n155_), .B1(ori_ori_n81_), .Y(ori_ori_n309_));
  NO2        o293(.A(ori_ori_n41_), .B(x0), .Y(ori_ori_n310_));
  OR2        o294(.A(ori_ori_n303_), .B(ori_ori_n310_), .Y(ori_ori_n311_));
  NO2        o295(.A(ori_ori_n128_), .B(ori_ori_n92_), .Y(ori_ori_n312_));
  AOI220     o296(.A0(ori_ori_n312_), .A1(ori_ori_n311_), .B0(ori_ori_n309_), .B1(ori_ori_n59_), .Y(ori_ori_n313_));
  NO2        o297(.A(ori_ori_n33_), .B(x2), .Y(ori_ori_n314_));
  NO2        o298(.A(ori_ori_n313_), .B(ori_ori_n60_), .Y(ori_ori_n315_));
  OAI220     o299(.A0(ori_ori_n315_), .A1(x6), .B0(ori_ori_n308_), .B1(ori_ori_n301_), .Y(ori_ori_n316_));
  OAI210     o300(.A0(x6), .A1(ori_ori_n46_), .B0(ori_ori_n40_), .Y(ori_ori_n317_));
  OAI210     o301(.A0(ori_ori_n317_), .A1(ori_ori_n81_), .B0(ori_ori_n269_), .Y(ori_ori_n318_));
  AOI210     o302(.A0(ori_ori_n318_), .A1(ori_ori_n18_), .B0(ori_ori_n130_), .Y(ori_ori_n319_));
  AO220      o303(.A0(ori_ori_n319_), .A1(ori_ori_n316_), .B0(ori_ori_n297_), .B1(ori_ori_n285_), .Y(ori_ori_n320_));
  NA2        o304(.A(ori_ori_n314_), .B(x6), .Y(ori_ori_n321_));
  AOI210     o305(.A0(x6), .A1(x1), .B0(ori_ori_n129_), .Y(ori_ori_n322_));
  NA2        o306(.A(ori_ori_n303_), .B(x0), .Y(ori_ori_n323_));
  NA2        o307(.A(ori_ori_n76_), .B(x6), .Y(ori_ori_n324_));
  OAI210     o308(.A0(ori_ori_n323_), .A1(ori_ori_n322_), .B0(ori_ori_n324_), .Y(ori_ori_n325_));
  AOI220     o309(.A0(ori_ori_n325_), .A1(ori_ori_n321_), .B0(ori_ori_n184_), .B1(ori_ori_n47_), .Y(ori_ori_n326_));
  NA2        o310(.A(ori_ori_n326_), .B(ori_ori_n320_), .Y(ori_ori_n327_));
  OAI210     o311(.A0(ori_ori_n27_), .A1(x1), .B0(ori_ori_n196_), .Y(ori_ori_n328_));
  AO220      o312(.A0(ori_ori_n328_), .A1(ori_ori_n127_), .B0(ori_ori_n96_), .B1(x4), .Y(ori_ori_n329_));
  NA3        o313(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n330_));
  NA2        o314(.A(ori_ori_n187_), .B(x0), .Y(ori_ori_n331_));
  OAI220     o315(.A0(ori_ori_n331_), .A1(ori_ori_n177_), .B0(ori_ori_n330_), .B1(ori_ori_n302_), .Y(ori_ori_n332_));
  AOI210     o316(.A0(ori_ori_n329_), .A1(ori_ori_n99_), .B0(ori_ori_n332_), .Y(ori_ori_n333_));
  NO2        o317(.A(ori_ori_n333_), .B(ori_ori_n24_), .Y(ori_ori_n334_));
  OAI210     o318(.A0(ori_ori_n169_), .A1(ori_ori_n63_), .B0(ori_ori_n174_), .Y(ori_ori_n335_));
  NA3        o319(.A(ori_ori_n171_), .B(ori_ori_n189_), .C(x8), .Y(ori_ori_n336_));
  AOI210     o320(.A0(ori_ori_n336_), .A1(ori_ori_n335_), .B0(ori_ori_n24_), .Y(ori_ori_n337_));
  NO2        o321(.A(ori_ori_n310_), .B(ori_ori_n156_), .Y(ori_ori_n338_));
  OAI210     o322(.A0(ori_ori_n338_), .A1(ori_ori_n337_), .B0(ori_ori_n127_), .Y(ori_ori_n339_));
  NAi31      o323(.An(ori_ori_n48_), .B(ori_ori_n248_), .C(ori_ori_n154_), .Y(ori_ori_n340_));
  NA2        o324(.A(ori_ori_n340_), .B(ori_ori_n339_), .Y(ori_ori_n341_));
  OAI210     o325(.A0(ori_ori_n341_), .A1(ori_ori_n334_), .B0(x6), .Y(ori_ori_n342_));
  NA3        o326(.A(ori_ori_n53_), .B(ori_ori_n36_), .C(ori_ori_n30_), .Y(ori_ori_n343_));
  NO2        o327(.A(ori_ori_n343_), .B(ori_ori_n31_), .Y(ori_ori_n344_));
  NO2        o328(.A(ori_ori_n130_), .B(x0), .Y(ori_ori_n345_));
  AOI220     o329(.A0(ori_ori_n345_), .A1(ori_ori_n187_), .B0(ori_ori_n169_), .B1(ori_ori_n130_), .Y(ori_ori_n346_));
  AOI210     o330(.A0(ori_ori_n106_), .A1(ori_ori_n218_), .B0(x1), .Y(ori_ori_n347_));
  OAI210     o331(.A0(ori_ori_n346_), .A1(x8), .B0(ori_ori_n347_), .Y(ori_ori_n348_));
  NAi31      o332(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n349_));
  OAI210     o333(.A0(ori_ori_n349_), .A1(x4), .B0(ori_ori_n141_), .Y(ori_ori_n350_));
  NA3        o334(.A(ori_ori_n350_), .B(ori_ori_n125_), .C(x9), .Y(ori_ori_n351_));
  NO4        o335(.A(ori_ori_n105_), .B(ori_ori_n258_), .C(x9), .D(x2), .Y(ori_ori_n352_));
  NOi21      o336(.An(ori_ori_n103_), .B(ori_ori_n155_), .Y(ori_ori_n353_));
  NO3        o337(.A(ori_ori_n353_), .B(ori_ori_n352_), .C(ori_ori_n18_), .Y(ori_ori_n354_));
  NA3        o338(.A(ori_ori_n354_), .B(ori_ori_n351_), .C(ori_ori_n48_), .Y(ori_ori_n355_));
  OAI210     o339(.A0(ori_ori_n348_), .A1(ori_ori_n344_), .B0(ori_ori_n355_), .Y(ori_ori_n356_));
  AOI210     o340(.A0(ori_ori_n36_), .A1(x9), .B0(ori_ori_n113_), .Y(ori_ori_n357_));
  NO3        o341(.A(ori_ori_n357_), .B(ori_ori_n103_), .C(ori_ori_n41_), .Y(ori_ori_n358_));
  NOi31      o342(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n359_));
  AOI210     o343(.A0(x1), .A1(ori_ori_n58_), .B0(ori_ori_n102_), .Y(ori_ori_n360_));
  NO2        o344(.A(ori_ori_n360_), .B(x3), .Y(ori_ori_n361_));
  NO3        o345(.A(ori_ori_n361_), .B(ori_ori_n358_), .C(x2), .Y(ori_ori_n362_));
  OAI210     o346(.A0(ori_ori_n258_), .A1(ori_ori_n41_), .B0(ori_ori_n299_), .Y(ori_ori_n363_));
  AOI210     o347(.A0(x9), .A1(ori_ori_n46_), .B0(ori_ori_n330_), .Y(ori_ori_n364_));
  AOI220     o348(.A0(ori_ori_n364_), .A1(ori_ori_n81_), .B0(ori_ori_n363_), .B1(ori_ori_n130_), .Y(ori_ori_n365_));
  NO2        o349(.A(ori_ori_n365_), .B(ori_ori_n52_), .Y(ori_ori_n366_));
  NO2        o350(.A(ori_ori_n366_), .B(ori_ori_n362_), .Y(ori_ori_n367_));
  AOI210     o351(.A0(ori_ori_n367_), .A1(ori_ori_n356_), .B0(ori_ori_n24_), .Y(ori_ori_n368_));
  NA4        o352(.A(ori_ori_n30_), .B(ori_ori_n81_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n369_));
  NA2        o353(.A(ori_ori_n192_), .B(x7), .Y(ori_ori_n370_));
  NA3        o354(.A(ori_ori_n370_), .B(ori_ori_n129_), .C(ori_ori_n114_), .Y(ori_ori_n371_));
  NA2        o355(.A(ori_ori_n371_), .B(ori_ori_n369_), .Y(ori_ori_n372_));
  OAI210     o356(.A0(ori_ori_n372_), .A1(ori_ori_n368_), .B0(ori_ori_n34_), .Y(ori_ori_n373_));
  INV        o357(.A(ori_ori_n174_), .Y(ori_ori_n374_));
  NO4        o358(.A(ori_ori_n374_), .B(ori_ori_n71_), .C(x4), .D(ori_ori_n52_), .Y(ori_ori_n375_));
  NA2        o359(.A(ori_ori_n223_), .B(ori_ori_n21_), .Y(ori_ori_n376_));
  NO2        o360(.A(ori_ori_n138_), .B(ori_ori_n115_), .Y(ori_ori_n377_));
  NA2        o361(.A(ori_ori_n377_), .B(ori_ori_n376_), .Y(ori_ori_n378_));
  AOI210     o362(.A0(ori_ori_n378_), .A1(ori_ori_n144_), .B0(ori_ori_n27_), .Y(ori_ori_n379_));
  AOI220     o363(.A0(ori_ori_n310_), .A1(ori_ori_n81_), .B0(ori_ori_n128_), .B1(ori_ori_n171_), .Y(ori_ori_n380_));
  NA3        o364(.A(ori_ori_n380_), .B(ori_ori_n349_), .C(ori_ori_n79_), .Y(ori_ori_n381_));
  NA2        o365(.A(ori_ori_n381_), .B(ori_ori_n154_), .Y(ori_ori_n382_));
  NA2        o366(.A(x3), .B(ori_ori_n52_), .Y(ori_ori_n383_));
  OAI210     o367(.A0(ori_ori_n127_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n384_));
  NO3        o368(.A(ori_ori_n359_), .B(x3), .C(ori_ori_n52_), .Y(ori_ori_n385_));
  NA2        o369(.A(ori_ori_n385_), .B(ori_ori_n384_), .Y(ori_ori_n386_));
  OAI210     o370(.A0(ori_ori_n131_), .A1(ori_ori_n383_), .B0(ori_ori_n386_), .Y(ori_ori_n387_));
  NA2        o371(.A(ori_ori_n387_), .B(x0), .Y(ori_ori_n388_));
  AOI210     o372(.A0(ori_ori_n388_), .A1(ori_ori_n382_), .B0(ori_ori_n200_), .Y(ori_ori_n389_));
  NO3        o373(.A(ori_ori_n389_), .B(ori_ori_n379_), .C(ori_ori_n375_), .Y(ori_ori_n390_));
  NA3        o374(.A(ori_ori_n390_), .B(ori_ori_n373_), .C(ori_ori_n342_), .Y(ori_ori_n391_));
  AOI210     o375(.A0(ori_ori_n327_), .A1(ori_ori_n24_), .B0(ori_ori_n391_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO4        m012(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .D(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  NA2        m021(.A(x4), .B(x3), .Y(mai_mai_n38_));
  NO2        m022(.A(mai_mai_n23_), .B(mai_mai_n38_), .Y(mai_mai_n39_));
  NO2        m023(.A(x2), .B(x0), .Y(mai_mai_n40_));
  INV        m024(.A(x3), .Y(mai_mai_n41_));
  NO2        m025(.A(mai_mai_n41_), .B(mai_mai_n18_), .Y(mai_mai_n42_));
  INV        m026(.A(mai_mai_n42_), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n44_));
  OAI210     m028(.A0(mai_mai_n44_), .A1(mai_mai_n43_), .B0(mai_mai_n40_), .Y(mai_mai_n45_));
  INV        m029(.A(x4), .Y(mai_mai_n46_));
  NO2        m030(.A(mai_mai_n46_), .B(mai_mai_n17_), .Y(mai_mai_n47_));
  NA2        m031(.A(mai_mai_n47_), .B(x2), .Y(mai_mai_n48_));
  OAI210     m032(.A0(mai_mai_n48_), .A1(mai_mai_n20_), .B0(mai_mai_n45_), .Y(mai_mai_n49_));
  AOI210     m033(.A0(mai_mai_n22_), .A1(mai_mai_n19_), .B0(mai_mai_n35_), .Y(mai_mai_n50_));
  INV        m034(.A(x2), .Y(mai_mai_n51_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n17_), .Y(mai_mai_n52_));
  NA2        m036(.A(mai_mai_n41_), .B(mai_mai_n18_), .Y(mai_mai_n53_));
  NA2        m037(.A(mai_mai_n53_), .B(mai_mai_n52_), .Y(mai_mai_n54_));
  OAI210     m038(.A0(mai_mai_n50_), .A1(mai_mai_n32_), .B0(mai_mai_n54_), .Y(mai_mai_n55_));
  NO3        m039(.A(mai_mai_n55_), .B(mai_mai_n49_), .C(mai_mai_n39_), .Y(mai01));
  NA2        m040(.A(x8), .B(x7), .Y(mai_mai_n57_));
  NA2        m041(.A(mai_mai_n41_), .B(x1), .Y(mai_mai_n58_));
  INV        m042(.A(x9), .Y(mai_mai_n59_));
  NO2        m043(.A(mai_mai_n59_), .B(mai_mai_n36_), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n58_), .B(mai_mai_n57_), .Y(mai_mai_n61_));
  NO2        m045(.A(x7), .B(x6), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n58_), .B(x5), .Y(mai_mai_n63_));
  NO2        m047(.A(x8), .B(x2), .Y(mai_mai_n64_));
  INV        m048(.A(mai_mai_n64_), .Y(mai_mai_n65_));
  NO2        m049(.A(mai_mai_n65_), .B(x1), .Y(mai_mai_n66_));
  OA210      m050(.A0(mai_mai_n66_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .Y(mai_mai_n67_));
  OAI210     m051(.A0(mai_mai_n42_), .A1(mai_mai_n25_), .B0(mai_mai_n51_), .Y(mai_mai_n68_));
  OAI210     m052(.A0(mai_mai_n53_), .A1(mai_mai_n20_), .B0(mai_mai_n68_), .Y(mai_mai_n69_));
  NAi31      m053(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n70_));
  OAI220     m054(.A0(mai_mai_n70_), .A1(mai_mai_n41_), .B0(mai_mai_n69_), .B1(mai_mai_n67_), .Y(mai_mai_n71_));
  OAI210     m055(.A0(mai_mai_n71_), .A1(mai_mai_n61_), .B0(x4), .Y(mai_mai_n72_));
  NA2        m056(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n73_));
  OAI210     m057(.A0(mai_mai_n73_), .A1(mai_mai_n53_), .B0(x0), .Y(mai_mai_n74_));
  NA2        m058(.A(x5), .B(x3), .Y(mai_mai_n75_));
  NO2        m059(.A(x8), .B(x6), .Y(mai_mai_n76_));
  NO4        m060(.A(mai_mai_n76_), .B(mai_mai_n75_), .C(mai_mai_n62_), .D(mai_mai_n51_), .Y(mai_mai_n77_));
  NAi21      m061(.An(x4), .B(x3), .Y(mai_mai_n78_));
  INV        m062(.A(mai_mai_n78_), .Y(mai_mai_n79_));
  NO2        m063(.A(mai_mai_n79_), .B(mai_mai_n22_), .Y(mai_mai_n80_));
  NO2        m064(.A(x4), .B(x2), .Y(mai_mai_n81_));
  NO2        m065(.A(mai_mai_n81_), .B(x3), .Y(mai_mai_n82_));
  NO3        m066(.A(mai_mai_n82_), .B(mai_mai_n80_), .C(mai_mai_n18_), .Y(mai_mai_n83_));
  NO3        m067(.A(mai_mai_n83_), .B(mai_mai_n77_), .C(mai_mai_n74_), .Y(mai_mai_n84_));
  NO4        m068(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n41_), .D(x1), .Y(mai_mai_n85_));
  INV        m069(.A(x4), .Y(mai_mai_n86_));
  NA2        m070(.A(mai_mai_n85_), .B(mai_mai_n86_), .Y(mai_mai_n87_));
  NA2        m071(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n88_));
  NO2        m072(.A(mai_mai_n88_), .B(mai_mai_n25_), .Y(mai_mai_n89_));
  INV        m073(.A(x8), .Y(mai_mai_n90_));
  NA2        m074(.A(x2), .B(x1), .Y(mai_mai_n91_));
  NO2        m075(.A(mai_mai_n91_), .B(mai_mai_n90_), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n92_), .B(mai_mai_n89_), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n93_), .B(mai_mai_n26_), .Y(mai_mai_n94_));
  AOI210     m078(.A0(mai_mai_n53_), .A1(mai_mai_n25_), .B0(mai_mai_n51_), .Y(mai_mai_n95_));
  OAI210     m079(.A0(mai_mai_n43_), .A1(mai_mai_n37_), .B0(mai_mai_n46_), .Y(mai_mai_n96_));
  NO3        m080(.A(mai_mai_n96_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n97_));
  NA2        m081(.A(x4), .B(mai_mai_n41_), .Y(mai_mai_n98_));
  NO2        m082(.A(mai_mai_n46_), .B(mai_mai_n51_), .Y(mai_mai_n99_));
  NO2        m083(.A(mai_mai_n98_), .B(x1), .Y(mai_mai_n100_));
  NO2        m084(.A(x3), .B(x2), .Y(mai_mai_n101_));
  NA2        m085(.A(mai_mai_n101_), .B(mai_mai_n25_), .Y(mai_mai_n102_));
  AOI210     m086(.A0(x8), .A1(x6), .B0(mai_mai_n102_), .Y(mai_mai_n103_));
  NA2        m087(.A(mai_mai_n51_), .B(x1), .Y(mai_mai_n104_));
  OAI210     m088(.A0(mai_mai_n104_), .A1(mai_mai_n38_), .B0(mai_mai_n17_), .Y(mai_mai_n105_));
  NO4        m089(.A(mai_mai_n105_), .B(mai_mai_n103_), .C(mai_mai_n100_), .D(mai_mai_n97_), .Y(mai_mai_n106_));
  AO220      m090(.A0(mai_mai_n106_), .A1(mai_mai_n87_), .B0(mai_mai_n84_), .B1(mai_mai_n72_), .Y(mai02));
  NO2        m091(.A(x3), .B(mai_mai_n51_), .Y(mai_mai_n108_));
  NO2        m092(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n109_));
  NA2        m093(.A(mai_mai_n51_), .B(mai_mai_n17_), .Y(mai_mai_n110_));
  NA2        m094(.A(mai_mai_n41_), .B(x0), .Y(mai_mai_n111_));
  OAI210     m095(.A0(x4), .A1(mai_mai_n110_), .B0(mai_mai_n111_), .Y(mai_mai_n112_));
  AOI220     m096(.A0(mai_mai_n112_), .A1(mai_mai_n109_), .B0(mai_mai_n108_), .B1(x4), .Y(mai_mai_n113_));
  NO3        m097(.A(mai_mai_n113_), .B(x7), .C(x5), .Y(mai_mai_n114_));
  NA2        m098(.A(x9), .B(x2), .Y(mai_mai_n115_));
  OR2        m099(.A(x8), .B(x0), .Y(mai_mai_n116_));
  INV        m100(.A(mai_mai_n116_), .Y(mai_mai_n117_));
  NAi21      m101(.An(x2), .B(x8), .Y(mai_mai_n118_));
  INV        m102(.A(mai_mai_n118_), .Y(mai_mai_n119_));
  NO2        m103(.A(x4), .B(x1), .Y(mai_mai_n120_));
  NA3        m104(.A(mai_mai_n120_), .B(mai_mai_n414_), .C(mai_mai_n57_), .Y(mai_mai_n121_));
  NOi21      m105(.An(x0), .B(x1), .Y(mai_mai_n122_));
  NO3        m106(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n123_));
  NOi21      m107(.An(x0), .B(x4), .Y(mai_mai_n124_));
  NAi21      m108(.An(x8), .B(x7), .Y(mai_mai_n125_));
  NO2        m109(.A(mai_mai_n125_), .B(mai_mai_n59_), .Y(mai_mai_n126_));
  AOI220     m110(.A0(mai_mai_n126_), .A1(mai_mai_n124_), .B0(mai_mai_n123_), .B1(mai_mai_n122_), .Y(mai_mai_n127_));
  AOI210     m111(.A0(mai_mai_n127_), .A1(mai_mai_n121_), .B0(mai_mai_n75_), .Y(mai_mai_n128_));
  NO2        m112(.A(x5), .B(mai_mai_n46_), .Y(mai_mai_n129_));
  NA2        m113(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n130_));
  AOI210     m114(.A0(mai_mai_n130_), .A1(mai_mai_n104_), .B0(mai_mai_n111_), .Y(mai_mai_n131_));
  OAI210     m115(.A0(mai_mai_n131_), .A1(mai_mai_n35_), .B0(mai_mai_n129_), .Y(mai_mai_n132_));
  NAi21      m116(.An(x0), .B(x4), .Y(mai_mai_n133_));
  NO2        m117(.A(x7), .B(x0), .Y(mai_mai_n134_));
  NO2        m118(.A(mai_mai_n81_), .B(mai_mai_n99_), .Y(mai_mai_n135_));
  NO2        m119(.A(mai_mai_n135_), .B(x3), .Y(mai_mai_n136_));
  NA2        m120(.A(mai_mai_n134_), .B(mai_mai_n136_), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n21_), .B(mai_mai_n41_), .Y(mai_mai_n138_));
  NA2        m122(.A(x5), .B(x0), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n140_));
  NA3        m124(.A(mai_mai_n140_), .B(mai_mai_n139_), .C(mai_mai_n138_), .Y(mai_mai_n141_));
  NA4        m125(.A(mai_mai_n141_), .B(mai_mai_n137_), .C(mai_mai_n132_), .D(mai_mai_n36_), .Y(mai_mai_n142_));
  NO3        m126(.A(mai_mai_n142_), .B(mai_mai_n128_), .C(mai_mai_n114_), .Y(mai_mai_n143_));
  NO3        m127(.A(mai_mai_n75_), .B(mai_mai_n73_), .C(mai_mai_n24_), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n145_));
  AOI220     m129(.A0(mai_mai_n122_), .A1(mai_mai_n145_), .B0(mai_mai_n63_), .B1(mai_mai_n17_), .Y(mai_mai_n146_));
  NO3        m130(.A(mai_mai_n146_), .B(mai_mai_n57_), .C(mai_mai_n59_), .Y(mai_mai_n147_));
  NA2        m131(.A(x7), .B(x3), .Y(mai_mai_n148_));
  NO2        m132(.A(mai_mai_n98_), .B(x5), .Y(mai_mai_n149_));
  NO2        m133(.A(x9), .B(x7), .Y(mai_mai_n150_));
  NOi21      m134(.An(x8), .B(x0), .Y(mai_mai_n151_));
  AN2        m135(.A(x1), .B(mai_mai_n151_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n41_), .B(x2), .Y(mai_mai_n153_));
  INV        m137(.A(x7), .Y(mai_mai_n154_));
  NA2        m138(.A(mai_mai_n154_), .B(mai_mai_n18_), .Y(mai_mai_n155_));
  NA2        m139(.A(mai_mai_n155_), .B(mai_mai_n153_), .Y(mai_mai_n156_));
  NO2        m140(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n157_));
  NO2        m141(.A(mai_mai_n157_), .B(mai_mai_n124_), .Y(mai_mai_n158_));
  NO2        m142(.A(mai_mai_n158_), .B(mai_mai_n156_), .Y(mai_mai_n159_));
  AOI210     m143(.A0(mai_mai_n152_), .A1(mai_mai_n149_), .B0(mai_mai_n159_), .Y(mai_mai_n160_));
  OAI210     m144(.A0(mai_mai_n148_), .A1(mai_mai_n48_), .B0(mai_mai_n160_), .Y(mai_mai_n161_));
  NA2        m145(.A(x5), .B(x1), .Y(mai_mai_n162_));
  INV        m146(.A(mai_mai_n162_), .Y(mai_mai_n163_));
  AOI210     m147(.A0(mai_mai_n163_), .A1(mai_mai_n124_), .B0(mai_mai_n36_), .Y(mai_mai_n164_));
  NO2        m148(.A(mai_mai_n59_), .B(mai_mai_n90_), .Y(mai_mai_n165_));
  INV        m149(.A(mai_mai_n164_), .Y(mai_mai_n166_));
  NO4        m150(.A(mai_mai_n166_), .B(mai_mai_n161_), .C(mai_mai_n147_), .D(mai_mai_n144_), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n167_), .B(mai_mai_n143_), .Y(mai_mai_n168_));
  NO2        m152(.A(mai_mai_n139_), .B(mai_mai_n135_), .Y(mai_mai_n169_));
  NA2        m153(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n170_));
  NA2        m154(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n171_));
  NA3        m155(.A(mai_mai_n171_), .B(mai_mai_n170_), .C(mai_mai_n24_), .Y(mai_mai_n172_));
  AN2        m156(.A(mai_mai_n172_), .B(mai_mai_n140_), .Y(mai_mai_n173_));
  NA2        m157(.A(x8), .B(x0), .Y(mai_mai_n174_));
  NO2        m158(.A(mai_mai_n154_), .B(mai_mai_n25_), .Y(mai_mai_n175_));
  NO2        m159(.A(mai_mai_n122_), .B(x4), .Y(mai_mai_n176_));
  NA2        m160(.A(mai_mai_n176_), .B(mai_mai_n175_), .Y(mai_mai_n177_));
  AOI210     m161(.A0(mai_mai_n174_), .A1(mai_mai_n130_), .B0(mai_mai_n177_), .Y(mai_mai_n178_));
  NA2        m162(.A(x2), .B(x0), .Y(mai_mai_n179_));
  NA2        m163(.A(x4), .B(x1), .Y(mai_mai_n180_));
  NAi21      m164(.An(mai_mai_n120_), .B(mai_mai_n180_), .Y(mai_mai_n181_));
  NOi31      m165(.An(mai_mai_n181_), .B(mai_mai_n157_), .C(mai_mai_n179_), .Y(mai_mai_n182_));
  NO4        m166(.A(mai_mai_n182_), .B(mai_mai_n178_), .C(mai_mai_n173_), .D(mai_mai_n169_), .Y(mai_mai_n183_));
  NO2        m167(.A(mai_mai_n183_), .B(mai_mai_n41_), .Y(mai_mai_n184_));
  NO2        m168(.A(mai_mai_n172_), .B(mai_mai_n73_), .Y(mai_mai_n185_));
  INV        m169(.A(mai_mai_n129_), .Y(mai_mai_n186_));
  NO2        m170(.A(mai_mai_n104_), .B(mai_mai_n17_), .Y(mai_mai_n187_));
  AOI210     m171(.A0(mai_mai_n35_), .A1(mai_mai_n90_), .B0(mai_mai_n187_), .Y(mai_mai_n188_));
  NO3        m172(.A(mai_mai_n188_), .B(mai_mai_n186_), .C(x7), .Y(mai_mai_n189_));
  NA3        m173(.A(mai_mai_n181_), .B(mai_mai_n186_), .C(mai_mai_n40_), .Y(mai_mai_n190_));
  OAI210     m174(.A0(mai_mai_n171_), .A1(mai_mai_n135_), .B0(mai_mai_n190_), .Y(mai_mai_n191_));
  NO3        m175(.A(mai_mai_n191_), .B(mai_mai_n189_), .C(mai_mai_n185_), .Y(mai_mai_n192_));
  NO2        m176(.A(mai_mai_n192_), .B(x3), .Y(mai_mai_n193_));
  NO3        m177(.A(mai_mai_n193_), .B(mai_mai_n184_), .C(mai_mai_n168_), .Y(mai03));
  NO2        m178(.A(mai_mai_n46_), .B(x3), .Y(mai_mai_n195_));
  NO2        m179(.A(mai_mai_n51_), .B(x1), .Y(mai_mai_n196_));
  OAI210     m180(.A0(mai_mai_n196_), .A1(mai_mai_n25_), .B0(mai_mai_n60_), .Y(mai_mai_n197_));
  OAI220     m181(.A0(mai_mai_n197_), .A1(mai_mai_n17_), .B0(x6), .B1(mai_mai_n104_), .Y(mai_mai_n198_));
  NA2        m182(.A(mai_mai_n198_), .B(mai_mai_n195_), .Y(mai_mai_n199_));
  NO2        m183(.A(mai_mai_n75_), .B(x6), .Y(mai_mai_n200_));
  NA2        m184(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n201_), .B(x4), .Y(mai_mai_n202_));
  NO2        m186(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n203_));
  AN2        m187(.A(mai_mai_n200_), .B(mai_mai_n52_), .Y(mai_mai_n204_));
  INV        m188(.A(mai_mai_n204_), .Y(mai_mai_n205_));
  NA2        m189(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n206_));
  NO2        m190(.A(mai_mai_n206_), .B(mai_mai_n201_), .Y(mai_mai_n207_));
  NA2        m191(.A(x9), .B(mai_mai_n51_), .Y(mai_mai_n208_));
  NA2        m192(.A(mai_mai_n208_), .B(x4), .Y(mai_mai_n209_));
  NA2        m193(.A(mai_mai_n209_), .B(mai_mai_n207_), .Y(mai_mai_n210_));
  NO3        m194(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n211_));
  NO2        m195(.A(x5), .B(x1), .Y(mai_mai_n212_));
  AOI220     m196(.A0(mai_mai_n212_), .A1(mai_mai_n17_), .B0(mai_mai_n101_), .B1(x5), .Y(mai_mai_n213_));
  NO2        m197(.A(mai_mai_n206_), .B(mai_mai_n170_), .Y(mai_mai_n214_));
  AOI220     m198(.A0(mai_mai_n415_), .A1(mai_mai_n46_), .B0(mai_mai_n211_), .B1(mai_mai_n129_), .Y(mai_mai_n215_));
  NA4        m199(.A(mai_mai_n215_), .B(mai_mai_n210_), .C(mai_mai_n205_), .D(mai_mai_n199_), .Y(mai_mai_n216_));
  NO2        m200(.A(mai_mai_n46_), .B(mai_mai_n41_), .Y(mai_mai_n217_));
  NA2        m201(.A(mai_mai_n217_), .B(mai_mai_n19_), .Y(mai_mai_n218_));
  NO2        m202(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n219_));
  NO2        m203(.A(mai_mai_n219_), .B(x6), .Y(mai_mai_n220_));
  NOi21      m204(.An(mai_mai_n81_), .B(mai_mai_n220_), .Y(mai_mai_n221_));
  NA2        m205(.A(mai_mai_n59_), .B(mai_mai_n90_), .Y(mai_mai_n222_));
  NA2        m206(.A(mai_mai_n219_), .B(x6), .Y(mai_mai_n223_));
  AOI210     m207(.A0(mai_mai_n223_), .A1(mai_mai_n221_), .B0(mai_mai_n154_), .Y(mai_mai_n224_));
  AO210      m208(.A0(mai_mai_n224_), .A1(mai_mai_n218_), .B0(mai_mai_n175_), .Y(mai_mai_n225_));
  NA2        m209(.A(mai_mai_n41_), .B(mai_mai_n51_), .Y(mai_mai_n226_));
  NA2        m210(.A(mai_mai_n140_), .B(mai_mai_n89_), .Y(mai_mai_n227_));
  NA2        m211(.A(x6), .B(mai_mai_n46_), .Y(mai_mai_n228_));
  OAI210     m212(.A0(mai_mai_n117_), .A1(mai_mai_n76_), .B0(x4), .Y(mai_mai_n229_));
  AOI210     m213(.A0(mai_mai_n229_), .A1(mai_mai_n228_), .B0(mai_mai_n75_), .Y(mai_mai_n230_));
  NO2        m214(.A(mai_mai_n59_), .B(x6), .Y(mai_mai_n231_));
  NO2        m215(.A(mai_mai_n162_), .B(mai_mai_n41_), .Y(mai_mai_n232_));
  OAI210     m216(.A0(mai_mai_n232_), .A1(mai_mai_n214_), .B0(mai_mai_n231_), .Y(mai_mai_n233_));
  NA3        m217(.A(mai_mai_n206_), .B(mai_mai_n129_), .C(x6), .Y(mai_mai_n234_));
  OAI210     m218(.A0(mai_mai_n90_), .A1(mai_mai_n36_), .B0(mai_mai_n63_), .Y(mai_mai_n235_));
  NA3        m219(.A(mai_mai_n235_), .B(mai_mai_n234_), .C(mai_mai_n233_), .Y(mai_mai_n236_));
  OAI210     m220(.A0(mai_mai_n236_), .A1(mai_mai_n230_), .B0(x2), .Y(mai_mai_n237_));
  NA3        m221(.A(mai_mai_n237_), .B(mai_mai_n227_), .C(mai_mai_n225_), .Y(mai_mai_n238_));
  AOI210     m222(.A0(mai_mai_n216_), .A1(x8), .B0(mai_mai_n238_), .Y(mai_mai_n239_));
  NO2        m223(.A(mai_mai_n90_), .B(x3), .Y(mai_mai_n240_));
  NA2        m224(.A(mai_mai_n240_), .B(mai_mai_n202_), .Y(mai_mai_n241_));
  NO3        m225(.A(mai_mai_n88_), .B(mai_mai_n76_), .C(mai_mai_n25_), .Y(mai_mai_n242_));
  AOI210     m226(.A0(mai_mai_n220_), .A1(mai_mai_n157_), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  AOI210     m227(.A0(mai_mai_n243_), .A1(mai_mai_n241_), .B0(x2), .Y(mai_mai_n244_));
  NO2        m228(.A(x4), .B(mai_mai_n51_), .Y(mai_mai_n245_));
  AOI220     m229(.A0(mai_mai_n202_), .A1(mai_mai_n187_), .B0(mai_mai_n245_), .B1(mai_mai_n63_), .Y(mai_mai_n246_));
  NA2        m230(.A(mai_mai_n206_), .B(x6), .Y(mai_mai_n247_));
  NO2        m231(.A(mai_mai_n206_), .B(x6), .Y(mai_mai_n248_));
  NA2        m232(.A(mai_mai_n247_), .B(mai_mai_n145_), .Y(mai_mai_n249_));
  NA3        m233(.A(mai_mai_n249_), .B(mai_mai_n246_), .C(mai_mai_n154_), .Y(mai_mai_n250_));
  NAi21      m234(.An(x1), .B(x4), .Y(mai_mai_n251_));
  AOI210     m235(.A0(x3), .A1(x2), .B0(mai_mai_n46_), .Y(mai_mai_n252_));
  OAI210     m236(.A0(mai_mai_n139_), .A1(x3), .B0(mai_mai_n252_), .Y(mai_mai_n253_));
  NA2        m237(.A(mai_mai_n253_), .B(mai_mai_n251_), .Y(mai_mai_n254_));
  INV        m238(.A(mai_mai_n254_), .Y(mai_mai_n255_));
  NO2        m239(.A(x6), .B(x0), .Y(mai_mai_n256_));
  NA2        m240(.A(mai_mai_n104_), .B(mai_mai_n25_), .Y(mai_mai_n257_));
  NA2        m241(.A(x6), .B(x2), .Y(mai_mai_n258_));
  NO2        m242(.A(mai_mai_n258_), .B(mai_mai_n170_), .Y(mai_mai_n259_));
  AOI210     m243(.A0(mai_mai_n257_), .A1(mai_mai_n256_), .B0(mai_mai_n259_), .Y(mai_mai_n260_));
  OAI220     m244(.A0(mai_mai_n260_), .A1(mai_mai_n41_), .B0(mai_mai_n176_), .B1(mai_mai_n44_), .Y(mai_mai_n261_));
  NA2        m245(.A(mai_mai_n261_), .B(mai_mai_n255_), .Y(mai_mai_n262_));
  NA2        m246(.A(x9), .B(mai_mai_n41_), .Y(mai_mai_n263_));
  NO2        m247(.A(mai_mai_n263_), .B(mai_mai_n201_), .Y(mai_mai_n264_));
  OR3        m248(.A(mai_mai_n264_), .B(mai_mai_n200_), .C(mai_mai_n149_), .Y(mai_mai_n265_));
  NA2        m249(.A(x4), .B(x0), .Y(mai_mai_n266_));
  NO3        m250(.A(mai_mai_n70_), .B(mai_mai_n266_), .C(x6), .Y(mai_mai_n267_));
  AOI210     m251(.A0(mai_mai_n265_), .A1(mai_mai_n40_), .B0(mai_mai_n267_), .Y(mai_mai_n268_));
  AOI210     m252(.A0(mai_mai_n268_), .A1(mai_mai_n262_), .B0(x8), .Y(mai_mai_n269_));
  INV        m253(.A(mai_mai_n174_), .Y(mai_mai_n270_));
  NO3        m254(.A(mai_mai_n269_), .B(mai_mai_n250_), .C(mai_mai_n244_), .Y(mai_mai_n271_));
  NO2        m255(.A(mai_mai_n165_), .B(x1), .Y(mai_mai_n272_));
  NO3        m256(.A(mai_mai_n272_), .B(x3), .C(mai_mai_n36_), .Y(mai_mai_n273_));
  OAI210     m257(.A0(mai_mai_n273_), .A1(mai_mai_n248_), .B0(x2), .Y(mai_mai_n274_));
  OAI210     m258(.A0(mai_mai_n270_), .A1(x6), .B0(mai_mai_n42_), .Y(mai_mai_n275_));
  AOI210     m259(.A0(mai_mai_n275_), .A1(mai_mai_n274_), .B0(mai_mai_n186_), .Y(mai_mai_n276_));
  NOi21      m260(.An(mai_mai_n258_), .B(mai_mai_n17_), .Y(mai_mai_n277_));
  NA3        m261(.A(mai_mai_n277_), .B(mai_mai_n212_), .C(mai_mai_n38_), .Y(mai_mai_n278_));
  AOI210     m262(.A0(mai_mai_n36_), .A1(mai_mai_n51_), .B0(x0), .Y(mai_mai_n279_));
  NA3        m263(.A(mai_mai_n279_), .B(mai_mai_n163_), .C(mai_mai_n32_), .Y(mai_mai_n280_));
  NA2        m264(.A(x3), .B(x2), .Y(mai_mai_n281_));
  AOI220     m265(.A0(mai_mai_n281_), .A1(mai_mai_n226_), .B0(mai_mai_n280_), .B1(mai_mai_n278_), .Y(mai_mai_n282_));
  NAi21      m266(.An(x4), .B(x0), .Y(mai_mai_n283_));
  NO3        m267(.A(mai_mai_n283_), .B(mai_mai_n42_), .C(x2), .Y(mai_mai_n284_));
  OAI210     m268(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  NO2        m269(.A(x9), .B(x8), .Y(mai_mai_n286_));
  NA3        m270(.A(mai_mai_n286_), .B(mai_mai_n36_), .C(mai_mai_n51_), .Y(mai_mai_n287_));
  OAI210     m271(.A0(mai_mai_n279_), .A1(mai_mai_n277_), .B0(mai_mai_n287_), .Y(mai_mai_n288_));
  AOI220     m272(.A0(mai_mai_n288_), .A1(mai_mai_n79_), .B0(mai_mai_n18_), .B1(mai_mai_n31_), .Y(mai_mai_n289_));
  AOI210     m273(.A0(mai_mai_n289_), .A1(mai_mai_n285_), .B0(mai_mai_n25_), .Y(mai_mai_n290_));
  NO2        m274(.A(mai_mai_n279_), .B(mai_mai_n277_), .Y(mai_mai_n291_));
  NA2        m275(.A(mai_mai_n36_), .B(mai_mai_n41_), .Y(mai_mai_n292_));
  OR2        m276(.A(mai_mai_n292_), .B(mai_mai_n266_), .Y(mai_mai_n293_));
  NO2        m277(.A(mai_mai_n293_), .B(mai_mai_n162_), .Y(mai_mai_n294_));
  AO210      m278(.A0(mai_mai_n291_), .A1(mai_mai_n149_), .B0(mai_mai_n294_), .Y(mai_mai_n295_));
  NO4        m279(.A(mai_mai_n295_), .B(mai_mai_n290_), .C(mai_mai_n282_), .D(mai_mai_n276_), .Y(mai_mai_n296_));
  OAI210     m280(.A0(mai_mai_n271_), .A1(mai_mai_n239_), .B0(mai_mai_n296_), .Y(mai04));
  OAI210     m281(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n298_));
  NA3        m282(.A(mai_mai_n298_), .B(mai_mai_n256_), .C(mai_mai_n82_), .Y(mai_mai_n299_));
  AOI210     m283(.A0(mai_mai_n59_), .A1(x4), .B0(mai_mai_n110_), .Y(mai_mai_n300_));
  NA2        m284(.A(mai_mai_n300_), .B(mai_mai_n240_), .Y(mai_mai_n301_));
  NO2        m285(.A(mai_mai_n281_), .B(mai_mai_n203_), .Y(mai_mai_n302_));
  NA2        m286(.A(x9), .B(x0), .Y(mai_mai_n303_));
  AOI210     m287(.A0(mai_mai_n88_), .A1(mai_mai_n73_), .B0(mai_mai_n303_), .Y(mai_mai_n304_));
  OAI210     m288(.A0(mai_mai_n304_), .A1(mai_mai_n302_), .B0(mai_mai_n90_), .Y(mai_mai_n305_));
  NA3        m289(.A(mai_mai_n305_), .B(x6), .C(mai_mai_n301_), .Y(mai_mai_n306_));
  NA2        m290(.A(mai_mai_n306_), .B(x6), .Y(mai_mai_n307_));
  NO2        m291(.A(mai_mai_n208_), .B(mai_mai_n111_), .Y(mai_mai_n308_));
  NO3        m292(.A(x9), .B(mai_mai_n118_), .C(mai_mai_n18_), .Y(mai_mai_n309_));
  NO2        m293(.A(mai_mai_n309_), .B(mai_mai_n308_), .Y(mai_mai_n310_));
  OAI210     m294(.A0(mai_mai_n116_), .A1(mai_mai_n104_), .B0(mai_mai_n174_), .Y(mai_mai_n311_));
  NA3        m295(.A(mai_mai_n311_), .B(x6), .C(x3), .Y(mai_mai_n312_));
  NOi21      m296(.An(mai_mai_n151_), .B(mai_mai_n130_), .Y(mai_mai_n313_));
  INV        m297(.A(mai_mai_n292_), .Y(mai_mai_n314_));
  AOI210     m298(.A0(mai_mai_n313_), .A1(mai_mai_n60_), .B0(mai_mai_n314_), .Y(mai_mai_n315_));
  NA2        m299(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n316_));
  OAI210     m300(.A0(mai_mai_n104_), .A1(mai_mai_n17_), .B0(mai_mai_n316_), .Y(mai_mai_n317_));
  NA2        m301(.A(mai_mai_n317_), .B(mai_mai_n76_), .Y(mai_mai_n318_));
  NA4        m302(.A(mai_mai_n318_), .B(mai_mai_n315_), .C(mai_mai_n312_), .D(mai_mai_n310_), .Y(mai_mai_n319_));
  OAI210     m303(.A0(mai_mai_n109_), .A1(x3), .B0(mai_mai_n284_), .Y(mai_mai_n320_));
  NA3        m304(.A(mai_mai_n222_), .B(mai_mai_n211_), .C(mai_mai_n81_), .Y(mai_mai_n321_));
  NA3        m305(.A(mai_mai_n321_), .B(mai_mai_n320_), .C(mai_mai_n154_), .Y(mai_mai_n322_));
  AOI210     m306(.A0(mai_mai_n319_), .A1(x4), .B0(mai_mai_n322_), .Y(mai_mai_n323_));
  NOi21      m307(.An(x4), .B(x0), .Y(mai_mai_n324_));
  XO2        m308(.A(x4), .B(x0), .Y(mai_mai_n325_));
  OAI210     m309(.A0(mai_mai_n325_), .A1(mai_mai_n115_), .B0(mai_mai_n251_), .Y(mai_mai_n326_));
  AOI220     m310(.A0(mai_mai_n326_), .A1(x8), .B0(mai_mai_n324_), .B1(mai_mai_n91_), .Y(mai_mai_n327_));
  NO2        m311(.A(mai_mai_n327_), .B(x3), .Y(mai_mai_n328_));
  INV        m312(.A(mai_mai_n91_), .Y(mai_mai_n329_));
  NO2        m313(.A(mai_mai_n90_), .B(x4), .Y(mai_mai_n330_));
  AOI220     m314(.A0(mai_mai_n330_), .A1(mai_mai_n42_), .B0(mai_mai_n124_), .B1(mai_mai_n329_), .Y(mai_mai_n331_));
  NO3        m315(.A(mai_mai_n325_), .B(mai_mai_n165_), .C(x2), .Y(mai_mai_n332_));
  INV        m316(.A(mai_mai_n332_), .Y(mai_mai_n333_));
  NA4        m317(.A(mai_mai_n333_), .B(mai_mai_n331_), .C(mai_mai_n218_), .D(x6), .Y(mai_mai_n334_));
  NO2        m318(.A(mai_mai_n151_), .B(mai_mai_n78_), .Y(mai_mai_n335_));
  NO2        m319(.A(mai_mai_n35_), .B(x2), .Y(mai_mai_n336_));
  NOi21      m320(.An(mai_mai_n120_), .B(mai_mai_n27_), .Y(mai_mai_n337_));
  AOI210     m321(.A0(mai_mai_n336_), .A1(mai_mai_n335_), .B0(mai_mai_n337_), .Y(mai_mai_n338_));
  INV        m322(.A(mai_mai_n338_), .Y(mai_mai_n339_));
  OAI220     m323(.A0(mai_mai_n339_), .A1(x6), .B0(mai_mai_n334_), .B1(mai_mai_n328_), .Y(mai_mai_n340_));
  OAI210     m324(.A0(mai_mai_n60_), .A1(mai_mai_n46_), .B0(mai_mai_n40_), .Y(mai_mai_n341_));
  OAI210     m325(.A0(mai_mai_n341_), .A1(mai_mai_n90_), .B0(mai_mai_n293_), .Y(mai_mai_n342_));
  AOI210     m326(.A0(mai_mai_n342_), .A1(mai_mai_n18_), .B0(mai_mai_n154_), .Y(mai_mai_n343_));
  AO220      m327(.A0(mai_mai_n343_), .A1(mai_mai_n340_), .B0(mai_mai_n323_), .B1(mai_mai_n307_), .Y(mai_mai_n344_));
  NA2        m328(.A(mai_mai_n344_), .B(mai_mai_n299_), .Y(mai_mai_n345_));
  AOI210     m329(.A0(mai_mai_n196_), .A1(x8), .B0(mai_mai_n109_), .Y(mai_mai_n346_));
  NA2        m330(.A(mai_mai_n346_), .B(mai_mai_n316_), .Y(mai_mai_n347_));
  NA3        m331(.A(mai_mai_n347_), .B(mai_mai_n195_), .C(mai_mai_n154_), .Y(mai_mai_n348_));
  OAI210     m332(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n226_), .Y(mai_mai_n349_));
  AO220      m333(.A0(mai_mai_n349_), .A1(mai_mai_n150_), .B0(mai_mai_n108_), .B1(x4), .Y(mai_mai_n350_));
  NA3        m334(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n351_));
  NA2        m335(.A(mai_mai_n217_), .B(x0), .Y(mai_mai_n352_));
  OAI220     m336(.A0(mai_mai_n352_), .A1(mai_mai_n208_), .B0(mai_mai_n351_), .B1(mai_mai_n329_), .Y(mai_mai_n353_));
  AOI210     m337(.A0(mai_mai_n350_), .A1(mai_mai_n117_), .B0(mai_mai_n353_), .Y(mai_mai_n354_));
  AOI210     m338(.A0(mai_mai_n354_), .A1(mai_mai_n348_), .B0(mai_mai_n25_), .Y(mai_mai_n355_));
  NA3        m339(.A(mai_mai_n119_), .B(mai_mai_n217_), .C(x0), .Y(mai_mai_n356_));
  AOI210     m340(.A0(mai_mai_n118_), .A1(mai_mai_n116_), .B0(mai_mai_n40_), .Y(mai_mai_n357_));
  NAi31      m341(.An(mai_mai_n48_), .B(mai_mai_n272_), .C(mai_mai_n175_), .Y(mai_mai_n358_));
  NA2        m342(.A(mai_mai_n358_), .B(mai_mai_n356_), .Y(mai_mai_n359_));
  OAI210     m343(.A0(mai_mai_n359_), .A1(mai_mai_n355_), .B0(x6), .Y(mai_mai_n360_));
  INV        m344(.A(mai_mai_n134_), .Y(mai_mai_n361_));
  AOI210     m345(.A0(mai_mai_n38_), .A1(mai_mai_n32_), .B0(mai_mai_n361_), .Y(mai_mai_n362_));
  NO2        m346(.A(mai_mai_n154_), .B(x0), .Y(mai_mai_n363_));
  AOI220     m347(.A0(mai_mai_n363_), .A1(mai_mai_n217_), .B0(mai_mai_n195_), .B1(mai_mai_n154_), .Y(mai_mai_n364_));
  AOI210     m348(.A0(mai_mai_n126_), .A1(mai_mai_n245_), .B0(x1), .Y(mai_mai_n365_));
  OAI210     m349(.A0(mai_mai_n364_), .A1(x8), .B0(mai_mai_n365_), .Y(mai_mai_n366_));
  NO3        m350(.A(mai_mai_n125_), .B(mai_mai_n283_), .C(x2), .Y(mai_mai_n367_));
  NO2        m351(.A(mai_mai_n367_), .B(mai_mai_n18_), .Y(mai_mai_n368_));
  NO3        m352(.A(x9), .B(mai_mai_n154_), .C(x0), .Y(mai_mai_n369_));
  AOI220     m353(.A0(mai_mai_n369_), .A1(mai_mai_n240_), .B0(mai_mai_n335_), .B1(mai_mai_n154_), .Y(mai_mai_n370_));
  NA3        m354(.A(mai_mai_n370_), .B(mai_mai_n368_), .C(mai_mai_n48_), .Y(mai_mai_n371_));
  OAI210     m355(.A0(mai_mai_n366_), .A1(mai_mai_n362_), .B0(mai_mai_n371_), .Y(mai_mai_n372_));
  NOi31      m356(.An(mai_mai_n363_), .B(mai_mai_n32_), .C(x8), .Y(mai_mai_n373_));
  INV        m357(.A(mai_mai_n133_), .Y(mai_mai_n374_));
  NO3        m358(.A(mai_mai_n374_), .B(mai_mai_n123_), .C(mai_mai_n41_), .Y(mai_mai_n375_));
  NOi31      m359(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n376_));
  AOI220     m360(.A0(mai_mai_n376_), .A1(mai_mai_n324_), .B0(mai_mai_n124_), .B1(x3), .Y(mai_mai_n377_));
  AOI210     m361(.A0(mai_mai_n251_), .A1(mai_mai_n57_), .B0(mai_mai_n122_), .Y(mai_mai_n378_));
  OAI210     m362(.A0(mai_mai_n378_), .A1(x3), .B0(mai_mai_n377_), .Y(mai_mai_n379_));
  NO3        m363(.A(mai_mai_n379_), .B(mai_mai_n375_), .C(x2), .Y(mai_mai_n380_));
  OAI220     m364(.A0(mai_mai_n325_), .A1(mai_mai_n286_), .B0(mai_mai_n283_), .B1(mai_mai_n41_), .Y(mai_mai_n381_));
  NA2        m365(.A(mai_mai_n381_), .B(mai_mai_n154_), .Y(mai_mai_n382_));
  NO2        m366(.A(mai_mai_n382_), .B(mai_mai_n51_), .Y(mai_mai_n383_));
  NO3        m367(.A(mai_mai_n383_), .B(mai_mai_n380_), .C(mai_mai_n373_), .Y(mai_mai_n384_));
  AOI210     m368(.A0(mai_mai_n384_), .A1(mai_mai_n372_), .B0(mai_mai_n25_), .Y(mai_mai_n385_));
  NO3        m369(.A(mai_mai_n59_), .B(x4), .C(x1), .Y(mai_mai_n386_));
  NO3        m370(.A(mai_mai_n64_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n387_));
  AOI220     m371(.A0(mai_mai_n387_), .A1(mai_mai_n252_), .B0(mai_mai_n386_), .B1(mai_mai_n357_), .Y(mai_mai_n388_));
  NO2        m372(.A(mai_mai_n388_), .B(mai_mai_n101_), .Y(mai_mai_n389_));
  NO3        m373(.A(mai_mai_n413_), .B(mai_mai_n174_), .C(mai_mai_n38_), .Y(mai_mai_n390_));
  OAI210     m374(.A0(mai_mai_n390_), .A1(mai_mai_n389_), .B0(x7), .Y(mai_mai_n391_));
  INV        m375(.A(mai_mai_n391_), .Y(mai_mai_n392_));
  OAI210     m376(.A0(mai_mai_n392_), .A1(mai_mai_n385_), .B0(mai_mai_n36_), .Y(mai_mai_n393_));
  NO2        m377(.A(mai_mai_n369_), .B(mai_mai_n203_), .Y(mai_mai_n394_));
  NO4        m378(.A(mai_mai_n394_), .B(mai_mai_n75_), .C(x4), .D(mai_mai_n51_), .Y(mai_mai_n395_));
  INV        m379(.A(mai_mai_n88_), .Y(mai_mai_n396_));
  NA2        m380(.A(mai_mai_n396_), .B(mai_mai_n175_), .Y(mai_mai_n397_));
  OAI220     m381(.A0(mai_mai_n263_), .A1(mai_mai_n65_), .B0(mai_mai_n162_), .B1(mai_mai_n41_), .Y(mai_mai_n398_));
  NA2        m382(.A(x3), .B(mai_mai_n51_), .Y(mai_mai_n399_));
  INV        m383(.A(mai_mai_n70_), .Y(mai_mai_n400_));
  NO3        m384(.A(mai_mai_n376_), .B(x3), .C(mai_mai_n51_), .Y(mai_mai_n401_));
  NO2        m385(.A(mai_mai_n401_), .B(mai_mai_n400_), .Y(mai_mai_n402_));
  OAI210     m386(.A0(mai_mai_n155_), .A1(mai_mai_n399_), .B0(mai_mai_n402_), .Y(mai_mai_n403_));
  AOI220     m387(.A0(mai_mai_n403_), .A1(x0), .B0(mai_mai_n398_), .B1(mai_mai_n134_), .Y(mai_mai_n404_));
  AOI210     m388(.A0(mai_mai_n404_), .A1(mai_mai_n397_), .B0(mai_mai_n228_), .Y(mai_mai_n405_));
  INV        m389(.A(x5), .Y(mai_mai_n406_));
  NO4        m390(.A(mai_mai_n104_), .B(mai_mai_n406_), .C(mai_mai_n57_), .D(mai_mai_n32_), .Y(mai_mai_n407_));
  NO3        m391(.A(mai_mai_n407_), .B(mai_mai_n405_), .C(mai_mai_n395_), .Y(mai_mai_n408_));
  NA3        m392(.A(mai_mai_n408_), .B(mai_mai_n393_), .C(mai_mai_n360_), .Y(mai_mai_n409_));
  AOI210     m393(.A0(mai_mai_n345_), .A1(mai_mai_n25_), .B0(mai_mai_n409_), .Y(mai05));
  INV        m394(.A(x2), .Y(mai_mai_n413_));
  INV        m395(.A(mai_mai_n115_), .Y(mai_mai_n414_));
  INV        m396(.A(mai_mai_n213_), .Y(mai_mai_n415_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  INV        u012(.A(men_men_n24_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  AN2        u015(.A(men_men_n31_), .B(men_men_n19_), .Y(men_men_n32_));
  NOi31      u016(.An(men_men_n23_), .B(men_men_n32_), .C(men_men_n29_), .Y(men00));
  NO2        u017(.A(x1), .B(x0), .Y(men_men_n34_));
  INV        u018(.A(x6), .Y(men_men_n35_));
  NO2        u019(.A(men_men_n35_), .B(men_men_n25_), .Y(men_men_n36_));
  NA3        u020(.A(x7), .B(men_men_n36_), .C(men_men_n34_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  AOI210     u022(.A0(men_men_n37_), .A1(men_men_n23_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n36_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  NA2        u033(.A(x7), .B(men_men_n36_), .Y(men_men_n50_));
  AOI220     u034(.A0(men_men_n50_), .A1(men_men_n34_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n51_));
  INV        u035(.A(x2), .Y(men_men_n52_));
  NO2        u036(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  OAI210     u039(.A0(men_men_n51_), .A1(men_men_n31_), .B0(men_men_n55_), .Y(men_men_n56_));
  NO3        u040(.A(men_men_n56_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u041(.A(x8), .B(x7), .Y(men_men_n58_));
  NA2        u042(.A(men_men_n41_), .B(x1), .Y(men_men_n59_));
  INV        u043(.A(x9), .Y(men_men_n60_));
  NO2        u044(.A(men_men_n60_), .B(men_men_n35_), .Y(men_men_n61_));
  INV        u045(.A(men_men_n61_), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n62_), .B(men_men_n59_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n59_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  AN2        u051(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n68_));
  OAI210     u052(.A0(men_men_n42_), .A1(men_men_n25_), .B0(men_men_n52_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n54_), .A1(men_men_n20_), .B0(men_men_n69_), .Y(men_men_n70_));
  NAi31      u054(.An(x1), .B(x9), .C(x5), .Y(men_men_n71_));
  NO2        u055(.A(men_men_n70_), .B(men_men_n68_), .Y(men_men_n72_));
  OAI210     u056(.A0(men_men_n72_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n73_));
  NA2        u057(.A(men_men_n46_), .B(x2), .Y(men_men_n74_));
  OAI210     u058(.A0(men_men_n74_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n75_));
  NA2        u059(.A(x5), .B(x3), .Y(men_men_n76_));
  NO2        u060(.A(x8), .B(x6), .Y(men_men_n77_));
  NO4        u061(.A(men_men_n77_), .B(men_men_n76_), .C(men_men_n64_), .D(men_men_n52_), .Y(men_men_n78_));
  NAi21      u062(.An(x4), .B(x3), .Y(men_men_n79_));
  INV        u063(.A(men_men_n79_), .Y(men_men_n80_));
  NO2        u064(.A(men_men_n80_), .B(men_men_n22_), .Y(men_men_n81_));
  NO2        u065(.A(x4), .B(x2), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(x3), .Y(men_men_n83_));
  NO3        u067(.A(men_men_n83_), .B(men_men_n81_), .C(men_men_n18_), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n78_), .C(men_men_n75_), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n21_), .B(men_men_n41_), .C(x1), .Y(men_men_n86_));
  NA2        u070(.A(men_men_n60_), .B(men_men_n46_), .Y(men_men_n87_));
  INV        u071(.A(men_men_n87_), .Y(men_men_n88_));
  OAI210     u072(.A0(men_men_n86_), .A1(men_men_n65_), .B0(men_men_n88_), .Y(men_men_n89_));
  NA2        u073(.A(x3), .B(men_men_n18_), .Y(men_men_n90_));
  NO2        u074(.A(men_men_n90_), .B(men_men_n25_), .Y(men_men_n91_));
  INV        u075(.A(x8), .Y(men_men_n92_));
  NA2        u076(.A(x2), .B(x1), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n94_), .B(men_men_n91_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n26_), .Y(men_men_n96_));
  AOI210     u080(.A0(men_men_n54_), .A1(men_men_n25_), .B0(men_men_n52_), .Y(men_men_n97_));
  OAI210     u081(.A0(men_men_n43_), .A1(men_men_n36_), .B0(men_men_n46_), .Y(men_men_n98_));
  NO3        u082(.A(men_men_n98_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n99_));
  NA2        u083(.A(x4), .B(men_men_n41_), .Y(men_men_n100_));
  NO2        u084(.A(men_men_n46_), .B(men_men_n52_), .Y(men_men_n101_));
  OAI210     u085(.A0(men_men_n101_), .A1(men_men_n41_), .B0(men_men_n18_), .Y(men_men_n102_));
  AOI210     u086(.A0(men_men_n100_), .A1(men_men_n50_), .B0(men_men_n102_), .Y(men_men_n103_));
  NO2        u087(.A(x3), .B(x2), .Y(men_men_n104_));
  NA3        u088(.A(men_men_n104_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n105_));
  INV        u089(.A(men_men_n105_), .Y(men_men_n106_));
  NA2        u090(.A(men_men_n52_), .B(x1), .Y(men_men_n107_));
  OAI210     u091(.A0(men_men_n107_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n108_));
  NO4        u092(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n103_), .D(men_men_n99_), .Y(men_men_n109_));
  AO220      u093(.A0(men_men_n109_), .A1(men_men_n89_), .B0(men_men_n85_), .B1(men_men_n73_), .Y(men02));
  NO2        u094(.A(x3), .B(men_men_n52_), .Y(men_men_n111_));
  NO2        u095(.A(x8), .B(men_men_n18_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n41_), .B(x0), .Y(men_men_n113_));
  OAI210     u097(.A0(men_men_n87_), .A1(x2), .B0(men_men_n113_), .Y(men_men_n114_));
  AOI220     u098(.A0(men_men_n114_), .A1(men_men_n112_), .B0(men_men_n111_), .B1(x4), .Y(men_men_n115_));
  NO3        u099(.A(men_men_n115_), .B(x7), .C(x5), .Y(men_men_n116_));
  NA2        u100(.A(x9), .B(x2), .Y(men_men_n117_));
  OR2        u101(.A(x8), .B(x0), .Y(men_men_n118_));
  NAi21      u102(.An(x2), .B(x8), .Y(men_men_n119_));
  INV        u103(.A(men_men_n119_), .Y(men_men_n120_));
  NO2        u104(.A(x4), .B(x1), .Y(men_men_n121_));
  NA3        u105(.A(men_men_n121_), .B(men_men_n118_), .C(men_men_n58_), .Y(men_men_n122_));
  NOi21      u106(.An(x0), .B(x1), .Y(men_men_n123_));
  NO3        u107(.A(x9), .B(x8), .C(x7), .Y(men_men_n124_));
  NOi21      u108(.An(x0), .B(x4), .Y(men_men_n125_));
  NO2        u109(.A(men_men_n122_), .B(men_men_n76_), .Y(men_men_n126_));
  NO2        u110(.A(x5), .B(men_men_n46_), .Y(men_men_n127_));
  NA2        u111(.A(x2), .B(men_men_n18_), .Y(men_men_n128_));
  AOI210     u112(.A0(men_men_n128_), .A1(men_men_n107_), .B0(men_men_n113_), .Y(men_men_n129_));
  OAI210     u113(.A0(men_men_n129_), .A1(men_men_n34_), .B0(men_men_n127_), .Y(men_men_n130_));
  NAi21      u114(.An(x0), .B(x4), .Y(men_men_n131_));
  NO2        u115(.A(men_men_n131_), .B(x1), .Y(men_men_n132_));
  NO2        u116(.A(x7), .B(x0), .Y(men_men_n133_));
  NO2        u117(.A(men_men_n82_), .B(men_men_n101_), .Y(men_men_n134_));
  NO2        u118(.A(men_men_n134_), .B(x3), .Y(men_men_n135_));
  OAI210     u119(.A0(men_men_n133_), .A1(men_men_n132_), .B0(men_men_n135_), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n21_), .B(men_men_n41_), .Y(men_men_n137_));
  NA2        u121(.A(x5), .B(x0), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n46_), .B(x2), .Y(men_men_n139_));
  NA3        u123(.A(men_men_n139_), .B(men_men_n138_), .C(men_men_n137_), .Y(men_men_n140_));
  NA4        u124(.A(men_men_n140_), .B(men_men_n136_), .C(men_men_n130_), .D(men_men_n35_), .Y(men_men_n141_));
  NO3        u125(.A(men_men_n141_), .B(men_men_n126_), .C(men_men_n116_), .Y(men_men_n142_));
  NO2        u126(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n143_));
  AOI220     u127(.A0(men_men_n123_), .A1(men_men_n143_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n144_), .B(men_men_n58_), .Y(men_men_n145_));
  NA2        u129(.A(x7), .B(x3), .Y(men_men_n146_));
  NO2        u130(.A(men_men_n100_), .B(x5), .Y(men_men_n147_));
  NO2        u131(.A(x9), .B(x7), .Y(men_men_n148_));
  NOi21      u132(.An(x8), .B(x0), .Y(men_men_n149_));
  NO2        u133(.A(men_men_n41_), .B(x2), .Y(men_men_n150_));
  INV        u134(.A(x7), .Y(men_men_n151_));
  NA2        u135(.A(men_men_n151_), .B(men_men_n18_), .Y(men_men_n152_));
  AOI220     u136(.A0(men_men_n152_), .A1(men_men_n150_), .B0(men_men_n111_), .B1(x7), .Y(men_men_n153_));
  NO2        u137(.A(men_men_n25_), .B(x4), .Y(men_men_n154_));
  NO2        u138(.A(men_men_n154_), .B(men_men_n125_), .Y(men_men_n155_));
  NO2        u139(.A(men_men_n155_), .B(men_men_n153_), .Y(men_men_n156_));
  NA2        u140(.A(x5), .B(x1), .Y(men_men_n157_));
  INV        u141(.A(men_men_n157_), .Y(men_men_n158_));
  AOI210     u142(.A0(men_men_n158_), .A1(men_men_n125_), .B0(men_men_n35_), .Y(men_men_n159_));
  NO2        u143(.A(men_men_n60_), .B(men_men_n92_), .Y(men_men_n160_));
  NAi21      u144(.An(x2), .B(x7), .Y(men_men_n161_));
  NO3        u145(.A(men_men_n161_), .B(men_men_n160_), .C(men_men_n46_), .Y(men_men_n162_));
  NA2        u146(.A(men_men_n162_), .B(men_men_n65_), .Y(men_men_n163_));
  NAi31      u147(.An(men_men_n76_), .B(x7), .C(men_men_n34_), .Y(men_men_n164_));
  NA3        u148(.A(men_men_n164_), .B(men_men_n163_), .C(men_men_n159_), .Y(men_men_n165_));
  NO3        u149(.A(men_men_n165_), .B(men_men_n156_), .C(men_men_n145_), .Y(men_men_n166_));
  NO2        u150(.A(men_men_n166_), .B(men_men_n142_), .Y(men_men_n167_));
  NO2        u151(.A(men_men_n138_), .B(men_men_n134_), .Y(men_men_n168_));
  NA2        u152(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n169_));
  NA2        u153(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n170_));
  NA3        u154(.A(men_men_n170_), .B(men_men_n169_), .C(men_men_n24_), .Y(men_men_n171_));
  AN2        u155(.A(men_men_n171_), .B(men_men_n139_), .Y(men_men_n172_));
  NA2        u156(.A(x8), .B(x0), .Y(men_men_n173_));
  NO2        u157(.A(men_men_n151_), .B(men_men_n25_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n123_), .B(x4), .Y(men_men_n175_));
  NA2        u159(.A(men_men_n175_), .B(men_men_n174_), .Y(men_men_n176_));
  AOI210     u160(.A0(men_men_n173_), .A1(men_men_n128_), .B0(men_men_n176_), .Y(men_men_n177_));
  NA2        u161(.A(x2), .B(x0), .Y(men_men_n178_));
  NA2        u162(.A(x4), .B(x1), .Y(men_men_n179_));
  NAi21      u163(.An(men_men_n121_), .B(men_men_n179_), .Y(men_men_n180_));
  NOi31      u164(.An(men_men_n180_), .B(men_men_n154_), .C(men_men_n178_), .Y(men_men_n181_));
  NO4        u165(.A(men_men_n181_), .B(men_men_n177_), .C(men_men_n172_), .D(men_men_n168_), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n182_), .B(men_men_n41_), .Y(men_men_n183_));
  NO2        u167(.A(men_men_n171_), .B(men_men_n74_), .Y(men_men_n184_));
  INV        u168(.A(men_men_n127_), .Y(men_men_n185_));
  NO2        u169(.A(men_men_n107_), .B(men_men_n17_), .Y(men_men_n186_));
  NO2        u170(.A(men_men_n34_), .B(men_men_n186_), .Y(men_men_n187_));
  NO3        u171(.A(men_men_n187_), .B(men_men_n185_), .C(x7), .Y(men_men_n188_));
  NA3        u172(.A(men_men_n180_), .B(men_men_n185_), .C(men_men_n40_), .Y(men_men_n189_));
  OAI210     u173(.A0(men_men_n170_), .A1(men_men_n134_), .B0(men_men_n189_), .Y(men_men_n190_));
  NO3        u174(.A(men_men_n190_), .B(men_men_n188_), .C(men_men_n184_), .Y(men_men_n191_));
  NO2        u175(.A(men_men_n191_), .B(x3), .Y(men_men_n192_));
  NO3        u176(.A(men_men_n192_), .B(men_men_n183_), .C(men_men_n167_), .Y(men03));
  NO2        u177(.A(men_men_n46_), .B(x3), .Y(men_men_n194_));
  NO2        u178(.A(x6), .B(men_men_n25_), .Y(men_men_n195_));
  NO2        u179(.A(men_men_n52_), .B(x1), .Y(men_men_n196_));
  OAI210     u180(.A0(men_men_n196_), .A1(men_men_n25_), .B0(men_men_n61_), .Y(men_men_n197_));
  NO2        u181(.A(men_men_n197_), .B(men_men_n17_), .Y(men_men_n198_));
  NA2        u182(.A(men_men_n198_), .B(men_men_n194_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n76_), .B(x6), .Y(men_men_n200_));
  NA2        u184(.A(x6), .B(men_men_n25_), .Y(men_men_n201_));
  NO2        u185(.A(men_men_n201_), .B(x4), .Y(men_men_n202_));
  NO2        u186(.A(men_men_n18_), .B(x0), .Y(men_men_n203_));
  AO220      u187(.A0(men_men_n203_), .A1(men_men_n202_), .B0(men_men_n200_), .B1(men_men_n53_), .Y(men_men_n204_));
  NA2        u188(.A(men_men_n204_), .B(men_men_n60_), .Y(men_men_n205_));
  NA2        u189(.A(x3), .B(men_men_n17_), .Y(men_men_n206_));
  NA2        u190(.A(men_men_n201_), .B(men_men_n79_), .Y(men_men_n207_));
  AOI210     u191(.A0(men_men_n25_), .A1(x3), .B0(men_men_n178_), .Y(men_men_n208_));
  NA2        u192(.A(men_men_n208_), .B(men_men_n207_), .Y(men_men_n209_));
  NO2        u193(.A(x5), .B(x1), .Y(men_men_n210_));
  AOI220     u194(.A0(men_men_n210_), .A1(men_men_n17_), .B0(men_men_n104_), .B1(x5), .Y(men_men_n211_));
  NO2        u195(.A(men_men_n206_), .B(men_men_n169_), .Y(men_men_n212_));
  NO3        u196(.A(x3), .B(x2), .C(x1), .Y(men_men_n213_));
  NO2        u197(.A(men_men_n213_), .B(men_men_n212_), .Y(men_men_n214_));
  OAI210     u198(.A0(men_men_n211_), .A1(men_men_n62_), .B0(men_men_n214_), .Y(men_men_n215_));
  NA2        u199(.A(men_men_n215_), .B(men_men_n46_), .Y(men_men_n216_));
  NA4        u200(.A(men_men_n216_), .B(men_men_n209_), .C(men_men_n205_), .D(men_men_n199_), .Y(men_men_n217_));
  NO2        u201(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n218_));
  NA2        u202(.A(men_men_n218_), .B(men_men_n19_), .Y(men_men_n219_));
  NO2        u203(.A(x3), .B(men_men_n17_), .Y(men_men_n220_));
  NO2        u204(.A(men_men_n220_), .B(x6), .Y(men_men_n221_));
  NOi21      u205(.An(men_men_n82_), .B(men_men_n221_), .Y(men_men_n222_));
  NO2        u206(.A(men_men_n222_), .B(men_men_n151_), .Y(men_men_n223_));
  AO210      u207(.A0(men_men_n223_), .A1(men_men_n219_), .B0(men_men_n174_), .Y(men_men_n224_));
  NA2        u208(.A(men_men_n41_), .B(men_men_n52_), .Y(men_men_n225_));
  OAI210     u209(.A0(men_men_n225_), .A1(men_men_n25_), .B0(men_men_n170_), .Y(men_men_n226_));
  NO2        u210(.A(men_men_n179_), .B(x6), .Y(men_men_n227_));
  AOI220     u211(.A0(men_men_n227_), .A1(men_men_n226_), .B0(men_men_n139_), .B1(men_men_n91_), .Y(men_men_n228_));
  NA2        u212(.A(x6), .B(men_men_n46_), .Y(men_men_n229_));
  NA2        u213(.A(men_men_n77_), .B(x4), .Y(men_men_n230_));
  AOI210     u214(.A0(men_men_n230_), .A1(men_men_n229_), .B0(men_men_n76_), .Y(men_men_n231_));
  NA2        u215(.A(men_men_n195_), .B(men_men_n132_), .Y(men_men_n232_));
  OAI210     u216(.A0(men_men_n92_), .A1(men_men_n35_), .B0(men_men_n65_), .Y(men_men_n233_));
  NA2        u217(.A(men_men_n233_), .B(men_men_n232_), .Y(men_men_n234_));
  OAI210     u218(.A0(men_men_n234_), .A1(men_men_n231_), .B0(x2), .Y(men_men_n235_));
  NA3        u219(.A(men_men_n235_), .B(men_men_n228_), .C(men_men_n224_), .Y(men_men_n236_));
  AOI210     u220(.A0(men_men_n217_), .A1(x8), .B0(men_men_n236_), .Y(men_men_n237_));
  NO2        u221(.A(men_men_n90_), .B(men_men_n25_), .Y(men_men_n238_));
  AOI210     u222(.A0(men_men_n221_), .A1(men_men_n154_), .B0(men_men_n238_), .Y(men_men_n239_));
  NO2        u223(.A(men_men_n239_), .B(x2), .Y(men_men_n240_));
  NO2        u224(.A(x4), .B(men_men_n52_), .Y(men_men_n241_));
  AOI220     u225(.A0(men_men_n202_), .A1(men_men_n186_), .B0(men_men_n241_), .B1(men_men_n65_), .Y(men_men_n242_));
  NA2        u226(.A(men_men_n60_), .B(x6), .Y(men_men_n243_));
  NA3        u227(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n244_));
  AOI210     u228(.A0(men_men_n244_), .A1(men_men_n138_), .B0(men_men_n243_), .Y(men_men_n245_));
  NA2        u229(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n246_));
  NO2        u230(.A(men_men_n246_), .B(men_men_n25_), .Y(men_men_n247_));
  OAI210     u231(.A0(men_men_n247_), .A1(men_men_n245_), .B0(men_men_n121_), .Y(men_men_n248_));
  NA2        u232(.A(men_men_n206_), .B(x6), .Y(men_men_n249_));
  NO2        u233(.A(men_men_n206_), .B(x6), .Y(men_men_n250_));
  NAi21      u234(.An(men_men_n160_), .B(men_men_n250_), .Y(men_men_n251_));
  NA3        u235(.A(men_men_n251_), .B(men_men_n249_), .C(men_men_n143_), .Y(men_men_n252_));
  NA4        u236(.A(men_men_n252_), .B(men_men_n248_), .C(men_men_n242_), .D(men_men_n151_), .Y(men_men_n253_));
  NA2        u237(.A(men_men_n195_), .B(men_men_n220_), .Y(men_men_n254_));
  NO2        u238(.A(x9), .B(x6), .Y(men_men_n255_));
  NO2        u239(.A(men_men_n138_), .B(men_men_n18_), .Y(men_men_n256_));
  NAi21      u240(.An(men_men_n256_), .B(men_men_n244_), .Y(men_men_n257_));
  NAi21      u241(.An(x1), .B(x4), .Y(men_men_n258_));
  AOI210     u242(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n259_));
  OAI210     u243(.A0(men_men_n138_), .A1(x3), .B0(men_men_n259_), .Y(men_men_n260_));
  AOI220     u244(.A0(men_men_n260_), .A1(men_men_n258_), .B0(men_men_n257_), .B1(men_men_n255_), .Y(men_men_n261_));
  NA2        u245(.A(men_men_n261_), .B(men_men_n254_), .Y(men_men_n262_));
  NA2        u246(.A(men_men_n60_), .B(x2), .Y(men_men_n263_));
  NO2        u247(.A(men_men_n263_), .B(men_men_n254_), .Y(men_men_n264_));
  NO3        u248(.A(x9), .B(x6), .C(x0), .Y(men_men_n265_));
  NA2        u249(.A(x6), .B(x2), .Y(men_men_n266_));
  NO2        u250(.A(men_men_n266_), .B(men_men_n169_), .Y(men_men_n267_));
  NO2        u251(.A(men_men_n265_), .B(men_men_n267_), .Y(men_men_n268_));
  OAI220     u252(.A0(men_men_n268_), .A1(men_men_n41_), .B0(men_men_n175_), .B1(men_men_n44_), .Y(men_men_n269_));
  OAI210     u253(.A0(men_men_n269_), .A1(men_men_n264_), .B0(men_men_n262_), .Y(men_men_n270_));
  NO2        u254(.A(x3), .B(men_men_n201_), .Y(men_men_n271_));
  OR2        u255(.A(men_men_n271_), .B(men_men_n200_), .Y(men_men_n272_));
  NA2        u256(.A(men_men_n272_), .B(men_men_n40_), .Y(men_men_n273_));
  AOI210     u257(.A0(men_men_n273_), .A1(men_men_n270_), .B0(x8), .Y(men_men_n274_));
  OAI210     u258(.A0(men_men_n256_), .A1(men_men_n210_), .B0(x6), .Y(men_men_n275_));
  INV        u259(.A(men_men_n173_), .Y(men_men_n276_));
  OAI210     u260(.A0(men_men_n276_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n277_));
  AOI210     u261(.A0(men_men_n277_), .A1(men_men_n275_), .B0(men_men_n225_), .Y(men_men_n278_));
  NO4        u262(.A(men_men_n278_), .B(men_men_n274_), .C(men_men_n253_), .D(men_men_n240_), .Y(men_men_n279_));
  NO2        u263(.A(x3), .B(men_men_n35_), .Y(men_men_n280_));
  OAI210     u264(.A0(men_men_n280_), .A1(men_men_n250_), .B0(x2), .Y(men_men_n281_));
  OAI210     u265(.A0(men_men_n276_), .A1(x6), .B0(men_men_n42_), .Y(men_men_n282_));
  AOI210     u266(.A0(men_men_n282_), .A1(men_men_n281_), .B0(men_men_n185_), .Y(men_men_n283_));
  NOi21      u267(.An(men_men_n266_), .B(men_men_n17_), .Y(men_men_n284_));
  NA3        u268(.A(men_men_n284_), .B(men_men_n210_), .C(men_men_n38_), .Y(men_men_n285_));
  AOI210     u269(.A0(men_men_n35_), .A1(men_men_n52_), .B0(x0), .Y(men_men_n286_));
  NA3        u270(.A(men_men_n286_), .B(men_men_n158_), .C(men_men_n31_), .Y(men_men_n287_));
  NA2        u271(.A(x3), .B(x2), .Y(men_men_n288_));
  AOI220     u272(.A0(men_men_n288_), .A1(men_men_n225_), .B0(men_men_n287_), .B1(men_men_n285_), .Y(men_men_n289_));
  NAi21      u273(.An(x4), .B(x0), .Y(men_men_n290_));
  NO3        u274(.A(men_men_n290_), .B(men_men_n42_), .C(x2), .Y(men_men_n291_));
  OAI210     u275(.A0(x6), .A1(men_men_n18_), .B0(men_men_n291_), .Y(men_men_n292_));
  OAI220     u276(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n293_));
  NO2        u277(.A(x9), .B(x8), .Y(men_men_n294_));
  NA3        u278(.A(men_men_n294_), .B(men_men_n35_), .C(men_men_n52_), .Y(men_men_n295_));
  OAI210     u279(.A0(men_men_n286_), .A1(men_men_n284_), .B0(men_men_n295_), .Y(men_men_n296_));
  AOI220     u280(.A0(men_men_n296_), .A1(men_men_n80_), .B0(men_men_n293_), .B1(men_men_n30_), .Y(men_men_n297_));
  AOI210     u281(.A0(men_men_n297_), .A1(men_men_n292_), .B0(men_men_n25_), .Y(men_men_n298_));
  NA3        u282(.A(men_men_n35_), .B(x1), .C(men_men_n17_), .Y(men_men_n299_));
  OAI210     u283(.A0(men_men_n286_), .A1(men_men_n284_), .B0(men_men_n299_), .Y(men_men_n300_));
  INV        u284(.A(men_men_n212_), .Y(men_men_n301_));
  NA2        u285(.A(men_men_n35_), .B(men_men_n41_), .Y(men_men_n302_));
  NO2        u286(.A(men_men_n229_), .B(men_men_n301_), .Y(men_men_n303_));
  AO210      u287(.A0(men_men_n300_), .A1(men_men_n147_), .B0(men_men_n303_), .Y(men_men_n304_));
  NO4        u288(.A(men_men_n304_), .B(men_men_n298_), .C(men_men_n289_), .D(men_men_n283_), .Y(men_men_n305_));
  OAI210     u289(.A0(men_men_n279_), .A1(men_men_n237_), .B0(men_men_n305_), .Y(men04));
  OAI210     u290(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n307_));
  NA3        u291(.A(men_men_n307_), .B(men_men_n265_), .C(men_men_n83_), .Y(men_men_n308_));
  NO2        u292(.A(x2), .B(x1), .Y(men_men_n309_));
  OAI210     u293(.A0(men_men_n246_), .A1(men_men_n309_), .B0(men_men_n35_), .Y(men_men_n310_));
  NO2        u294(.A(men_men_n309_), .B(men_men_n290_), .Y(men_men_n311_));
  NA2        u295(.A(men_men_n311_), .B(men_men_n426_), .Y(men_men_n312_));
  NO2        u296(.A(men_men_n263_), .B(men_men_n90_), .Y(men_men_n313_));
  NO2        u297(.A(men_men_n313_), .B(men_men_n35_), .Y(men_men_n314_));
  NO2        u298(.A(men_men_n288_), .B(men_men_n203_), .Y(men_men_n315_));
  NA2        u299(.A(men_men_n315_), .B(men_men_n92_), .Y(men_men_n316_));
  NA3        u300(.A(men_men_n316_), .B(men_men_n314_), .C(men_men_n312_), .Y(men_men_n317_));
  NA2        u301(.A(men_men_n317_), .B(men_men_n310_), .Y(men_men_n318_));
  INV        u302(.A(men_men_n128_), .Y(men_men_n319_));
  AOI210     u303(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n320_));
  OAI220     u304(.A0(men_men_n320_), .A1(men_men_n302_), .B0(men_men_n263_), .B1(men_men_n299_), .Y(men_men_n321_));
  AOI210     u305(.A0(men_men_n319_), .A1(men_men_n61_), .B0(men_men_n321_), .Y(men_men_n322_));
  NA2        u306(.A(x2), .B(men_men_n17_), .Y(men_men_n323_));
  OAI210     u307(.A0(men_men_n107_), .A1(men_men_n17_), .B0(men_men_n323_), .Y(men_men_n324_));
  AOI220     u308(.A0(men_men_n324_), .A1(men_men_n77_), .B0(men_men_n313_), .B1(men_men_n92_), .Y(men_men_n325_));
  NA2        u309(.A(men_men_n325_), .B(men_men_n322_), .Y(men_men_n326_));
  OAI210     u310(.A0(men_men_n112_), .A1(x3), .B0(men_men_n291_), .Y(men_men_n327_));
  NA2        u311(.A(men_men_n327_), .B(men_men_n151_), .Y(men_men_n328_));
  AOI210     u312(.A0(men_men_n326_), .A1(x4), .B0(men_men_n328_), .Y(men_men_n329_));
  NA2        u313(.A(men_men_n311_), .B(men_men_n92_), .Y(men_men_n330_));
  NOi21      u314(.An(x4), .B(x0), .Y(men_men_n331_));
  XO2        u315(.A(x4), .B(x0), .Y(men_men_n332_));
  OAI210     u316(.A0(men_men_n332_), .A1(men_men_n117_), .B0(men_men_n258_), .Y(men_men_n333_));
  AOI220     u317(.A0(men_men_n333_), .A1(x8), .B0(men_men_n331_), .B1(men_men_n93_), .Y(men_men_n334_));
  AOI210     u318(.A0(men_men_n334_), .A1(men_men_n330_), .B0(x3), .Y(men_men_n335_));
  INV        u319(.A(men_men_n93_), .Y(men_men_n336_));
  NO2        u320(.A(men_men_n92_), .B(x4), .Y(men_men_n337_));
  NA2        u321(.A(men_men_n337_), .B(men_men_n42_), .Y(men_men_n338_));
  NO3        u322(.A(men_men_n332_), .B(men_men_n160_), .C(x2), .Y(men_men_n339_));
  NO3        u323(.A(x9), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n340_));
  NO2        u324(.A(men_men_n340_), .B(men_men_n339_), .Y(men_men_n341_));
  NA4        u325(.A(men_men_n341_), .B(men_men_n338_), .C(men_men_n219_), .D(x6), .Y(men_men_n342_));
  NO2        u326(.A(men_men_n41_), .B(x0), .Y(men_men_n343_));
  OR2        u327(.A(men_men_n337_), .B(men_men_n343_), .Y(men_men_n344_));
  NO2        u328(.A(men_men_n149_), .B(men_men_n107_), .Y(men_men_n345_));
  AOI220     u329(.A0(men_men_n345_), .A1(men_men_n344_), .B0(men_men_n427_), .B1(men_men_n59_), .Y(men_men_n346_));
  NO2        u330(.A(men_men_n149_), .B(men_men_n79_), .Y(men_men_n347_));
  NO2        u331(.A(men_men_n34_), .B(x2), .Y(men_men_n348_));
  NOi21      u332(.An(men_men_n121_), .B(men_men_n27_), .Y(men_men_n349_));
  AOI210     u333(.A0(men_men_n348_), .A1(men_men_n347_), .B0(men_men_n349_), .Y(men_men_n350_));
  OAI210     u334(.A0(men_men_n346_), .A1(men_men_n60_), .B0(men_men_n350_), .Y(men_men_n351_));
  OAI220     u335(.A0(men_men_n351_), .A1(x6), .B0(men_men_n342_), .B1(men_men_n335_), .Y(men_men_n352_));
  AO220      u336(.A0(x7), .A1(men_men_n352_), .B0(men_men_n329_), .B1(men_men_n318_), .Y(men_men_n353_));
  NA2        u337(.A(men_men_n348_), .B(x6), .Y(men_men_n354_));
  AOI210     u338(.A0(x6), .A1(x1), .B0(men_men_n150_), .Y(men_men_n355_));
  NA2        u339(.A(men_men_n337_), .B(x0), .Y(men_men_n356_));
  NA2        u340(.A(men_men_n82_), .B(x6), .Y(men_men_n357_));
  OAI210     u341(.A0(men_men_n356_), .A1(men_men_n355_), .B0(men_men_n357_), .Y(men_men_n358_));
  AOI220     u342(.A0(men_men_n358_), .A1(men_men_n354_), .B0(men_men_n213_), .B1(men_men_n47_), .Y(men_men_n359_));
  NA3        u343(.A(men_men_n359_), .B(men_men_n353_), .C(men_men_n308_), .Y(men_men_n360_));
  AOI210     u344(.A0(men_men_n196_), .A1(x8), .B0(men_men_n112_), .Y(men_men_n361_));
  NA2        u345(.A(men_men_n361_), .B(men_men_n323_), .Y(men_men_n362_));
  NA3        u346(.A(men_men_n362_), .B(men_men_n194_), .C(men_men_n151_), .Y(men_men_n363_));
  NA3        u347(.A(x7), .B(x3), .C(x0), .Y(men_men_n364_));
  NO2        u348(.A(men_men_n364_), .B(men_men_n336_), .Y(men_men_n365_));
  INV        u349(.A(men_men_n365_), .Y(men_men_n366_));
  AOI210     u350(.A0(men_men_n366_), .A1(men_men_n363_), .B0(men_men_n25_), .Y(men_men_n367_));
  NA3        u351(.A(men_men_n120_), .B(men_men_n218_), .C(x0), .Y(men_men_n368_));
  OAI210     u352(.A0(men_men_n194_), .A1(men_men_n66_), .B0(men_men_n203_), .Y(men_men_n369_));
  NA3        u353(.A(men_men_n196_), .B(men_men_n220_), .C(x8), .Y(men_men_n370_));
  AOI210     u354(.A0(men_men_n370_), .A1(men_men_n369_), .B0(men_men_n25_), .Y(men_men_n371_));
  AOI210     u355(.A0(men_men_n119_), .A1(men_men_n118_), .B0(men_men_n40_), .Y(men_men_n372_));
  NOi31      u356(.An(men_men_n372_), .B(men_men_n343_), .C(men_men_n179_), .Y(men_men_n373_));
  OAI210     u357(.A0(men_men_n373_), .A1(men_men_n371_), .B0(men_men_n148_), .Y(men_men_n374_));
  NA2        u358(.A(men_men_n374_), .B(men_men_n368_), .Y(men_men_n375_));
  OAI210     u359(.A0(men_men_n375_), .A1(men_men_n367_), .B0(x6), .Y(men_men_n376_));
  OAI210     u360(.A0(men_men_n160_), .A1(men_men_n46_), .B0(men_men_n133_), .Y(men_men_n377_));
  NA3        u361(.A(men_men_n53_), .B(x7), .C(men_men_n30_), .Y(men_men_n378_));
  AOI220     u362(.A0(men_men_n378_), .A1(men_men_n377_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n379_));
  NAi31      u363(.An(x2), .B(x8), .C(x0), .Y(men_men_n380_));
  OAI210     u364(.A0(men_men_n380_), .A1(x4), .B0(men_men_n161_), .Y(men_men_n381_));
  NA3        u365(.A(men_men_n381_), .B(men_men_n146_), .C(x9), .Y(men_men_n382_));
  NOi21      u366(.An(men_men_n124_), .B(men_men_n178_), .Y(men_men_n383_));
  NO2        u367(.A(men_men_n383_), .B(men_men_n18_), .Y(men_men_n384_));
  NO3        u368(.A(x9), .B(men_men_n151_), .C(x0), .Y(men_men_n385_));
  AOI220     u369(.A0(men_men_n385_), .A1(men_men_n426_), .B0(men_men_n347_), .B1(men_men_n151_), .Y(men_men_n386_));
  NA3        u370(.A(men_men_n386_), .B(men_men_n384_), .C(men_men_n382_), .Y(men_men_n387_));
  OAI210     u371(.A0(x1), .A1(men_men_n379_), .B0(men_men_n387_), .Y(men_men_n388_));
  OAI220     u372(.A0(men_men_n332_), .A1(men_men_n294_), .B0(men_men_n290_), .B1(men_men_n41_), .Y(men_men_n389_));
  INV        u373(.A(men_men_n364_), .Y(men_men_n390_));
  AOI220     u374(.A0(men_men_n390_), .A1(men_men_n92_), .B0(men_men_n389_), .B1(men_men_n151_), .Y(men_men_n391_));
  NO2        u375(.A(men_men_n391_), .B(men_men_n52_), .Y(men_men_n392_));
  INV        u376(.A(men_men_n392_), .Y(men_men_n393_));
  AOI210     u377(.A0(men_men_n393_), .A1(men_men_n388_), .B0(men_men_n25_), .Y(men_men_n394_));
  NA4        u378(.A(men_men_n30_), .B(men_men_n92_), .C(x2), .D(men_men_n17_), .Y(men_men_n395_));
  NO3        u379(.A(men_men_n60_), .B(x4), .C(x1), .Y(men_men_n396_));
  NO3        u380(.A(men_men_n66_), .B(men_men_n18_), .C(x0), .Y(men_men_n397_));
  AOI220     u381(.A0(men_men_n397_), .A1(men_men_n259_), .B0(men_men_n396_), .B1(men_men_n372_), .Y(men_men_n398_));
  NO2        u382(.A(men_men_n398_), .B(men_men_n104_), .Y(men_men_n399_));
  NO3        u383(.A(men_men_n263_), .B(men_men_n173_), .C(men_men_n38_), .Y(men_men_n400_));
  OAI210     u384(.A0(men_men_n400_), .A1(men_men_n399_), .B0(x7), .Y(men_men_n401_));
  NA2        u385(.A(x9), .B(x7), .Y(men_men_n402_));
  NA3        u386(.A(men_men_n402_), .B(men_men_n150_), .C(men_men_n132_), .Y(men_men_n403_));
  NA3        u387(.A(men_men_n403_), .B(men_men_n401_), .C(men_men_n395_), .Y(men_men_n404_));
  OAI210     u388(.A0(men_men_n404_), .A1(men_men_n394_), .B0(men_men_n35_), .Y(men_men_n405_));
  NO2        u389(.A(men_men_n385_), .B(men_men_n203_), .Y(men_men_n406_));
  NO4        u390(.A(men_men_n406_), .B(men_men_n76_), .C(x4), .D(men_men_n52_), .Y(men_men_n407_));
  NA2        u391(.A(men_men_n246_), .B(men_men_n21_), .Y(men_men_n408_));
  NO2        u392(.A(men_men_n157_), .B(men_men_n133_), .Y(men_men_n409_));
  NA2        u393(.A(men_men_n409_), .B(men_men_n408_), .Y(men_men_n410_));
  AOI210     u394(.A0(men_men_n410_), .A1(men_men_n164_), .B0(men_men_n28_), .Y(men_men_n411_));
  AOI220     u395(.A0(men_men_n343_), .A1(men_men_n92_), .B0(men_men_n149_), .B1(men_men_n196_), .Y(men_men_n412_));
  NA3        u396(.A(men_men_n412_), .B(men_men_n380_), .C(men_men_n90_), .Y(men_men_n413_));
  NA2        u397(.A(men_men_n413_), .B(men_men_n174_), .Y(men_men_n414_));
  OAI220     u398(.A0(x3), .A1(men_men_n67_), .B0(men_men_n157_), .B1(men_men_n41_), .Y(men_men_n415_));
  AOI210     u399(.A0(men_men_n161_), .A1(men_men_n27_), .B0(men_men_n71_), .Y(men_men_n416_));
  AOI220     u400(.A0(men_men_n416_), .A1(x0), .B0(men_men_n415_), .B1(men_men_n133_), .Y(men_men_n417_));
  AOI210     u401(.A0(men_men_n417_), .A1(men_men_n414_), .B0(men_men_n229_), .Y(men_men_n418_));
  NA2        u402(.A(x9), .B(x5), .Y(men_men_n419_));
  NO4        u403(.A(men_men_n107_), .B(men_men_n419_), .C(men_men_n58_), .D(men_men_n31_), .Y(men_men_n420_));
  NO4        u404(.A(men_men_n420_), .B(men_men_n418_), .C(men_men_n411_), .D(men_men_n407_), .Y(men_men_n421_));
  NA3        u405(.A(men_men_n421_), .B(men_men_n405_), .C(men_men_n376_), .Y(men_men_n422_));
  AOI210     u406(.A0(men_men_n360_), .A1(men_men_n25_), .B0(men_men_n422_), .Y(men05));
  INV        u407(.A(x3), .Y(men_men_n426_));
  INV        u408(.A(men_men_n178_), .Y(men_men_n427_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule