library verilog;
use verilog.vl_types.all;
entity primeiro_vlg_check_tst is
    port(
        s               : in     vl_logic;
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end primeiro_vlg_check_tst;
